module gen_p(
  input  [2:0]   io_src,
  input  [131:0] io_x,
  output [131:0] io_p,
  output         io_c
);
  wire [2:0] gen_sel_io_src; // @[wallace_mul.scala 71:17]
  wire [3:0] gen_sel_io_out; // @[wallace_mul.scala 71:17]
  wire  gen_p_i_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_1_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_1_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_1_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_1_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_2_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_2_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_2_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_2_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_3_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_3_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_3_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_3_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_4_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_4_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_4_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_4_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_5_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_5_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_5_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_5_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_6_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_6_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_6_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_6_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_7_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_7_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_7_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_7_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_8_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_8_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_8_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_8_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_9_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_9_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_9_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_9_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_10_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_10_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_10_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_10_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_11_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_11_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_11_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_11_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_12_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_12_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_12_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_12_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_13_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_13_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_13_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_13_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_14_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_14_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_14_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_14_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_15_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_15_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_15_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_15_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_16_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_16_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_16_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_16_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_17_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_17_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_17_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_17_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_18_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_18_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_18_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_18_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_19_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_19_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_19_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_19_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_20_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_20_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_20_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_20_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_21_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_21_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_21_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_21_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_22_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_22_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_22_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_22_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_23_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_23_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_23_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_23_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_24_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_24_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_24_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_24_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_25_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_25_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_25_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_25_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_26_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_26_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_26_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_26_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_27_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_27_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_27_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_27_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_28_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_28_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_28_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_28_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_29_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_29_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_29_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_29_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_30_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_30_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_30_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_30_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_31_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_31_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_31_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_31_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_32_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_32_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_32_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_32_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_33_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_33_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_33_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_33_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_34_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_34_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_34_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_34_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_35_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_35_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_35_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_35_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_36_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_36_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_36_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_36_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_37_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_37_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_37_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_37_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_38_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_38_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_38_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_38_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_39_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_39_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_39_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_39_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_40_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_40_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_40_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_40_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_41_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_41_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_41_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_41_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_42_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_42_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_42_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_42_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_43_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_43_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_43_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_43_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_44_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_44_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_44_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_44_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_45_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_45_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_45_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_45_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_46_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_46_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_46_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_46_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_47_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_47_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_47_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_47_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_48_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_48_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_48_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_48_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_49_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_49_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_49_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_49_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_50_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_50_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_50_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_50_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_51_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_51_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_51_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_51_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_52_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_52_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_52_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_52_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_53_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_53_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_53_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_53_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_54_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_54_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_54_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_54_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_55_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_55_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_55_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_55_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_56_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_56_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_56_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_56_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_57_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_57_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_57_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_57_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_58_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_58_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_58_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_58_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_59_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_59_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_59_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_59_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_60_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_60_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_60_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_60_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_61_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_61_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_61_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_61_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_62_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_62_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_62_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_62_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_63_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_63_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_63_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_63_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_64_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_64_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_64_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_64_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_65_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_65_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_65_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_65_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_66_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_66_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_66_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_66_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_67_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_67_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_67_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_67_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_68_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_68_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_68_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_68_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_69_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_69_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_69_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_69_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_70_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_70_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_70_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_70_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_71_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_71_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_71_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_71_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_72_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_72_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_72_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_72_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_73_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_73_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_73_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_73_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_74_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_74_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_74_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_74_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_75_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_75_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_75_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_75_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_76_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_76_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_76_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_76_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_77_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_77_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_77_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_77_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_78_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_78_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_78_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_78_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_79_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_79_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_79_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_79_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_80_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_80_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_80_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_80_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_81_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_81_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_81_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_81_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_82_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_82_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_82_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_82_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_83_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_83_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_83_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_83_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_84_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_84_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_84_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_84_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_85_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_85_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_85_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_85_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_86_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_86_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_86_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_86_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_87_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_87_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_87_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_87_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_88_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_88_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_88_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_88_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_89_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_89_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_89_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_89_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_90_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_90_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_90_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_90_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_91_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_91_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_91_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_91_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_92_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_92_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_92_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_92_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_93_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_93_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_93_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_93_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_94_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_94_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_94_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_94_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_95_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_95_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_95_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_95_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_96_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_96_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_96_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_96_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_97_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_97_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_97_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_97_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_98_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_98_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_98_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_98_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_99_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_99_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_99_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_99_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_100_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_100_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_100_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_100_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_101_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_101_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_101_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_101_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_102_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_102_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_102_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_102_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_103_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_103_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_103_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_103_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_104_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_104_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_104_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_104_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_105_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_105_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_105_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_105_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_106_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_106_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_106_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_106_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_107_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_107_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_107_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_107_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_108_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_108_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_108_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_108_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_109_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_109_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_109_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_109_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_110_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_110_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_110_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_110_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_111_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_111_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_111_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_111_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_112_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_112_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_112_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_112_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_113_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_113_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_113_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_113_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_114_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_114_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_114_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_114_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_115_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_115_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_115_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_115_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_116_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_116_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_116_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_116_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_117_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_117_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_117_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_117_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_118_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_118_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_118_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_118_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_119_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_119_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_119_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_119_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_120_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_120_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_120_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_120_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_121_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_121_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_121_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_121_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_122_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_122_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_122_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_122_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_123_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_123_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_123_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_123_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_124_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_124_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_124_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_124_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_125_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_125_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_125_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_125_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_126_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_126_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_126_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_126_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_127_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_127_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_127_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_127_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_128_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_128_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_128_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_128_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_129_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_129_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_129_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_129_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_130_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_130_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_130_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_130_io_p; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_131_io_x; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_131_io_x_sub; // @[wallace_mul.scala 72:29]
  wire [3:0] gen_p_i_131_io_sel; // @[wallace_mul.scala 72:29]
  wire  gen_p_i_131_io_p; // @[wallace_mul.scala 72:29]
  wire [7:0] io_p_lo_lo_lo_lo = {gen_p_i_7_io_p,gen_p_i_6_io_p,gen_p_i_5_io_p,gen_p_i_4_io_p,gen_p_i_3_io_p,
    gen_p_i_2_io_p,gen_p_i_1_io_p,gen_p_i_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_lo_hi_lo = {gen_p_i_23_io_p,gen_p_i_22_io_p,gen_p_i_21_io_p,gen_p_i_20_io_p,gen_p_i_19_io_p,
    gen_p_i_18_io_p,gen_p_i_17_io_p,gen_p_i_16_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_lo_lo_hi = {gen_p_i_32_io_p,gen_p_i_31_io_p,gen_p_i_30_io_p,gen_p_i_29_io_p,gen_p_i_28_io_p,
    gen_p_i_27_io_p,gen_p_i_26_io_p,gen_p_i_25_io_p,gen_p_i_24_io_p,io_p_lo_lo_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_lo_lo = {io_p_lo_lo_hi,gen_p_i_15_io_p,gen_p_i_14_io_p,gen_p_i_13_io_p,gen_p_i_12_io_p,
    gen_p_i_11_io_p,gen_p_i_10_io_p,gen_p_i_9_io_p,gen_p_i_8_io_p,io_p_lo_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_hi_lo_lo = {gen_p_i_40_io_p,gen_p_i_39_io_p,gen_p_i_38_io_p,gen_p_i_37_io_p,gen_p_i_36_io_p,
    gen_p_i_35_io_p,gen_p_i_34_io_p,gen_p_i_33_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_hi_hi_lo = {gen_p_i_56_io_p,gen_p_i_55_io_p,gen_p_i_54_io_p,gen_p_i_53_io_p,gen_p_i_52_io_p,
    gen_p_i_51_io_p,gen_p_i_50_io_p,gen_p_i_49_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_lo_hi_hi = {gen_p_i_65_io_p,gen_p_i_64_io_p,gen_p_i_63_io_p,gen_p_i_62_io_p,gen_p_i_61_io_p,
    gen_p_i_60_io_p,gen_p_i_59_io_p,gen_p_i_58_io_p,gen_p_i_57_io_p,io_p_lo_hi_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_lo_hi = {io_p_lo_hi_hi,gen_p_i_48_io_p,gen_p_i_47_io_p,gen_p_i_46_io_p,gen_p_i_45_io_p,
    gen_p_i_44_io_p,gen_p_i_43_io_p,gen_p_i_42_io_p,gen_p_i_41_io_p,io_p_lo_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [65:0] io_p_lo = {io_p_lo_hi,io_p_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_lo_lo_lo = {gen_p_i_73_io_p,gen_p_i_72_io_p,gen_p_i_71_io_p,gen_p_i_70_io_p,gen_p_i_69_io_p,
    gen_p_i_68_io_p,gen_p_i_67_io_p,gen_p_i_66_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_lo_hi_lo = {gen_p_i_89_io_p,gen_p_i_88_io_p,gen_p_i_87_io_p,gen_p_i_86_io_p,gen_p_i_85_io_p,
    gen_p_i_84_io_p,gen_p_i_83_io_p,gen_p_i_82_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_hi_lo_hi = {gen_p_i_98_io_p,gen_p_i_97_io_p,gen_p_i_96_io_p,gen_p_i_95_io_p,gen_p_i_94_io_p,
    gen_p_i_93_io_p,gen_p_i_92_io_p,gen_p_i_91_io_p,gen_p_i_90_io_p,io_p_hi_lo_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_hi_lo = {io_p_hi_lo_hi,gen_p_i_81_io_p,gen_p_i_80_io_p,gen_p_i_79_io_p,gen_p_i_78_io_p,
    gen_p_i_77_io_p,gen_p_i_76_io_p,gen_p_i_75_io_p,gen_p_i_74_io_p,io_p_hi_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_hi_lo_lo = {gen_p_i_106_io_p,gen_p_i_105_io_p,gen_p_i_104_io_p,gen_p_i_103_io_p,gen_p_i_102_io_p,
    gen_p_i_101_io_p,gen_p_i_100_io_p,gen_p_i_99_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_hi_hi_lo = {gen_p_i_122_io_p,gen_p_i_121_io_p,gen_p_i_120_io_p,gen_p_i_119_io_p,gen_p_i_118_io_p,
    gen_p_i_117_io_p,gen_p_i_116_io_p,gen_p_i_115_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_hi_hi_hi = {gen_p_i_131_io_p,gen_p_i_130_io_p,gen_p_i_129_io_p,gen_p_i_128_io_p,gen_p_i_127_io_p,
    gen_p_i_126_io_p,gen_p_i_125_io_p,gen_p_i_124_io_p,gen_p_i_123_io_p,io_p_hi_hi_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_hi_hi = {io_p_hi_hi_hi,gen_p_i_114_io_p,gen_p_i_113_io_p,gen_p_i_112_io_p,gen_p_i_111_io_p,
    gen_p_i_110_io_p,gen_p_i_109_io_p,gen_p_i_108_io_p,gen_p_i_107_io_p,io_p_hi_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [65:0] io_p_hi = {io_p_hi_hi,io_p_hi_lo}; // @[Cat.scala 33:92]
  gen_sel gen_sel ( // @[wallace_mul.scala 71:17]
    .io_src(gen_sel_io_src),
    .io_out(gen_sel_io_out)
  );
  gen_p_i gen_p_i ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_io_x),
    .io_x_sub(gen_p_i_io_x_sub),
    .io_sel(gen_p_i_io_sel),
    .io_p(gen_p_i_io_p)
  );
  gen_p_i gen_p_i_1 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_1_io_x),
    .io_x_sub(gen_p_i_1_io_x_sub),
    .io_sel(gen_p_i_1_io_sel),
    .io_p(gen_p_i_1_io_p)
  );
  gen_p_i gen_p_i_2 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_2_io_x),
    .io_x_sub(gen_p_i_2_io_x_sub),
    .io_sel(gen_p_i_2_io_sel),
    .io_p(gen_p_i_2_io_p)
  );
  gen_p_i gen_p_i_3 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_3_io_x),
    .io_x_sub(gen_p_i_3_io_x_sub),
    .io_sel(gen_p_i_3_io_sel),
    .io_p(gen_p_i_3_io_p)
  );
  gen_p_i gen_p_i_4 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_4_io_x),
    .io_x_sub(gen_p_i_4_io_x_sub),
    .io_sel(gen_p_i_4_io_sel),
    .io_p(gen_p_i_4_io_p)
  );
  gen_p_i gen_p_i_5 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_5_io_x),
    .io_x_sub(gen_p_i_5_io_x_sub),
    .io_sel(gen_p_i_5_io_sel),
    .io_p(gen_p_i_5_io_p)
  );
  gen_p_i gen_p_i_6 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_6_io_x),
    .io_x_sub(gen_p_i_6_io_x_sub),
    .io_sel(gen_p_i_6_io_sel),
    .io_p(gen_p_i_6_io_p)
  );
  gen_p_i gen_p_i_7 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_7_io_x),
    .io_x_sub(gen_p_i_7_io_x_sub),
    .io_sel(gen_p_i_7_io_sel),
    .io_p(gen_p_i_7_io_p)
  );
  gen_p_i gen_p_i_8 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_8_io_x),
    .io_x_sub(gen_p_i_8_io_x_sub),
    .io_sel(gen_p_i_8_io_sel),
    .io_p(gen_p_i_8_io_p)
  );
  gen_p_i gen_p_i_9 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_9_io_x),
    .io_x_sub(gen_p_i_9_io_x_sub),
    .io_sel(gen_p_i_9_io_sel),
    .io_p(gen_p_i_9_io_p)
  );
  gen_p_i gen_p_i_10 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_10_io_x),
    .io_x_sub(gen_p_i_10_io_x_sub),
    .io_sel(gen_p_i_10_io_sel),
    .io_p(gen_p_i_10_io_p)
  );
  gen_p_i gen_p_i_11 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_11_io_x),
    .io_x_sub(gen_p_i_11_io_x_sub),
    .io_sel(gen_p_i_11_io_sel),
    .io_p(gen_p_i_11_io_p)
  );
  gen_p_i gen_p_i_12 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_12_io_x),
    .io_x_sub(gen_p_i_12_io_x_sub),
    .io_sel(gen_p_i_12_io_sel),
    .io_p(gen_p_i_12_io_p)
  );
  gen_p_i gen_p_i_13 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_13_io_x),
    .io_x_sub(gen_p_i_13_io_x_sub),
    .io_sel(gen_p_i_13_io_sel),
    .io_p(gen_p_i_13_io_p)
  );
  gen_p_i gen_p_i_14 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_14_io_x),
    .io_x_sub(gen_p_i_14_io_x_sub),
    .io_sel(gen_p_i_14_io_sel),
    .io_p(gen_p_i_14_io_p)
  );
  gen_p_i gen_p_i_15 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_15_io_x),
    .io_x_sub(gen_p_i_15_io_x_sub),
    .io_sel(gen_p_i_15_io_sel),
    .io_p(gen_p_i_15_io_p)
  );
  gen_p_i gen_p_i_16 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_16_io_x),
    .io_x_sub(gen_p_i_16_io_x_sub),
    .io_sel(gen_p_i_16_io_sel),
    .io_p(gen_p_i_16_io_p)
  );
  gen_p_i gen_p_i_17 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_17_io_x),
    .io_x_sub(gen_p_i_17_io_x_sub),
    .io_sel(gen_p_i_17_io_sel),
    .io_p(gen_p_i_17_io_p)
  );
  gen_p_i gen_p_i_18 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_18_io_x),
    .io_x_sub(gen_p_i_18_io_x_sub),
    .io_sel(gen_p_i_18_io_sel),
    .io_p(gen_p_i_18_io_p)
  );
  gen_p_i gen_p_i_19 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_19_io_x),
    .io_x_sub(gen_p_i_19_io_x_sub),
    .io_sel(gen_p_i_19_io_sel),
    .io_p(gen_p_i_19_io_p)
  );
  gen_p_i gen_p_i_20 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_20_io_x),
    .io_x_sub(gen_p_i_20_io_x_sub),
    .io_sel(gen_p_i_20_io_sel),
    .io_p(gen_p_i_20_io_p)
  );
  gen_p_i gen_p_i_21 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_21_io_x),
    .io_x_sub(gen_p_i_21_io_x_sub),
    .io_sel(gen_p_i_21_io_sel),
    .io_p(gen_p_i_21_io_p)
  );
  gen_p_i gen_p_i_22 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_22_io_x),
    .io_x_sub(gen_p_i_22_io_x_sub),
    .io_sel(gen_p_i_22_io_sel),
    .io_p(gen_p_i_22_io_p)
  );
  gen_p_i gen_p_i_23 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_23_io_x),
    .io_x_sub(gen_p_i_23_io_x_sub),
    .io_sel(gen_p_i_23_io_sel),
    .io_p(gen_p_i_23_io_p)
  );
  gen_p_i gen_p_i_24 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_24_io_x),
    .io_x_sub(gen_p_i_24_io_x_sub),
    .io_sel(gen_p_i_24_io_sel),
    .io_p(gen_p_i_24_io_p)
  );
  gen_p_i gen_p_i_25 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_25_io_x),
    .io_x_sub(gen_p_i_25_io_x_sub),
    .io_sel(gen_p_i_25_io_sel),
    .io_p(gen_p_i_25_io_p)
  );
  gen_p_i gen_p_i_26 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_26_io_x),
    .io_x_sub(gen_p_i_26_io_x_sub),
    .io_sel(gen_p_i_26_io_sel),
    .io_p(gen_p_i_26_io_p)
  );
  gen_p_i gen_p_i_27 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_27_io_x),
    .io_x_sub(gen_p_i_27_io_x_sub),
    .io_sel(gen_p_i_27_io_sel),
    .io_p(gen_p_i_27_io_p)
  );
  gen_p_i gen_p_i_28 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_28_io_x),
    .io_x_sub(gen_p_i_28_io_x_sub),
    .io_sel(gen_p_i_28_io_sel),
    .io_p(gen_p_i_28_io_p)
  );
  gen_p_i gen_p_i_29 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_29_io_x),
    .io_x_sub(gen_p_i_29_io_x_sub),
    .io_sel(gen_p_i_29_io_sel),
    .io_p(gen_p_i_29_io_p)
  );
  gen_p_i gen_p_i_30 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_30_io_x),
    .io_x_sub(gen_p_i_30_io_x_sub),
    .io_sel(gen_p_i_30_io_sel),
    .io_p(gen_p_i_30_io_p)
  );
  gen_p_i gen_p_i_31 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_31_io_x),
    .io_x_sub(gen_p_i_31_io_x_sub),
    .io_sel(gen_p_i_31_io_sel),
    .io_p(gen_p_i_31_io_p)
  );
  gen_p_i gen_p_i_32 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_32_io_x),
    .io_x_sub(gen_p_i_32_io_x_sub),
    .io_sel(gen_p_i_32_io_sel),
    .io_p(gen_p_i_32_io_p)
  );
  gen_p_i gen_p_i_33 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_33_io_x),
    .io_x_sub(gen_p_i_33_io_x_sub),
    .io_sel(gen_p_i_33_io_sel),
    .io_p(gen_p_i_33_io_p)
  );
  gen_p_i gen_p_i_34 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_34_io_x),
    .io_x_sub(gen_p_i_34_io_x_sub),
    .io_sel(gen_p_i_34_io_sel),
    .io_p(gen_p_i_34_io_p)
  );
  gen_p_i gen_p_i_35 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_35_io_x),
    .io_x_sub(gen_p_i_35_io_x_sub),
    .io_sel(gen_p_i_35_io_sel),
    .io_p(gen_p_i_35_io_p)
  );
  gen_p_i gen_p_i_36 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_36_io_x),
    .io_x_sub(gen_p_i_36_io_x_sub),
    .io_sel(gen_p_i_36_io_sel),
    .io_p(gen_p_i_36_io_p)
  );
  gen_p_i gen_p_i_37 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_37_io_x),
    .io_x_sub(gen_p_i_37_io_x_sub),
    .io_sel(gen_p_i_37_io_sel),
    .io_p(gen_p_i_37_io_p)
  );
  gen_p_i gen_p_i_38 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_38_io_x),
    .io_x_sub(gen_p_i_38_io_x_sub),
    .io_sel(gen_p_i_38_io_sel),
    .io_p(gen_p_i_38_io_p)
  );
  gen_p_i gen_p_i_39 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_39_io_x),
    .io_x_sub(gen_p_i_39_io_x_sub),
    .io_sel(gen_p_i_39_io_sel),
    .io_p(gen_p_i_39_io_p)
  );
  gen_p_i gen_p_i_40 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_40_io_x),
    .io_x_sub(gen_p_i_40_io_x_sub),
    .io_sel(gen_p_i_40_io_sel),
    .io_p(gen_p_i_40_io_p)
  );
  gen_p_i gen_p_i_41 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_41_io_x),
    .io_x_sub(gen_p_i_41_io_x_sub),
    .io_sel(gen_p_i_41_io_sel),
    .io_p(gen_p_i_41_io_p)
  );
  gen_p_i gen_p_i_42 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_42_io_x),
    .io_x_sub(gen_p_i_42_io_x_sub),
    .io_sel(gen_p_i_42_io_sel),
    .io_p(gen_p_i_42_io_p)
  );
  gen_p_i gen_p_i_43 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_43_io_x),
    .io_x_sub(gen_p_i_43_io_x_sub),
    .io_sel(gen_p_i_43_io_sel),
    .io_p(gen_p_i_43_io_p)
  );
  gen_p_i gen_p_i_44 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_44_io_x),
    .io_x_sub(gen_p_i_44_io_x_sub),
    .io_sel(gen_p_i_44_io_sel),
    .io_p(gen_p_i_44_io_p)
  );
  gen_p_i gen_p_i_45 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_45_io_x),
    .io_x_sub(gen_p_i_45_io_x_sub),
    .io_sel(gen_p_i_45_io_sel),
    .io_p(gen_p_i_45_io_p)
  );
  gen_p_i gen_p_i_46 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_46_io_x),
    .io_x_sub(gen_p_i_46_io_x_sub),
    .io_sel(gen_p_i_46_io_sel),
    .io_p(gen_p_i_46_io_p)
  );
  gen_p_i gen_p_i_47 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_47_io_x),
    .io_x_sub(gen_p_i_47_io_x_sub),
    .io_sel(gen_p_i_47_io_sel),
    .io_p(gen_p_i_47_io_p)
  );
  gen_p_i gen_p_i_48 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_48_io_x),
    .io_x_sub(gen_p_i_48_io_x_sub),
    .io_sel(gen_p_i_48_io_sel),
    .io_p(gen_p_i_48_io_p)
  );
  gen_p_i gen_p_i_49 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_49_io_x),
    .io_x_sub(gen_p_i_49_io_x_sub),
    .io_sel(gen_p_i_49_io_sel),
    .io_p(gen_p_i_49_io_p)
  );
  gen_p_i gen_p_i_50 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_50_io_x),
    .io_x_sub(gen_p_i_50_io_x_sub),
    .io_sel(gen_p_i_50_io_sel),
    .io_p(gen_p_i_50_io_p)
  );
  gen_p_i gen_p_i_51 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_51_io_x),
    .io_x_sub(gen_p_i_51_io_x_sub),
    .io_sel(gen_p_i_51_io_sel),
    .io_p(gen_p_i_51_io_p)
  );
  gen_p_i gen_p_i_52 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_52_io_x),
    .io_x_sub(gen_p_i_52_io_x_sub),
    .io_sel(gen_p_i_52_io_sel),
    .io_p(gen_p_i_52_io_p)
  );
  gen_p_i gen_p_i_53 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_53_io_x),
    .io_x_sub(gen_p_i_53_io_x_sub),
    .io_sel(gen_p_i_53_io_sel),
    .io_p(gen_p_i_53_io_p)
  );
  gen_p_i gen_p_i_54 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_54_io_x),
    .io_x_sub(gen_p_i_54_io_x_sub),
    .io_sel(gen_p_i_54_io_sel),
    .io_p(gen_p_i_54_io_p)
  );
  gen_p_i gen_p_i_55 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_55_io_x),
    .io_x_sub(gen_p_i_55_io_x_sub),
    .io_sel(gen_p_i_55_io_sel),
    .io_p(gen_p_i_55_io_p)
  );
  gen_p_i gen_p_i_56 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_56_io_x),
    .io_x_sub(gen_p_i_56_io_x_sub),
    .io_sel(gen_p_i_56_io_sel),
    .io_p(gen_p_i_56_io_p)
  );
  gen_p_i gen_p_i_57 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_57_io_x),
    .io_x_sub(gen_p_i_57_io_x_sub),
    .io_sel(gen_p_i_57_io_sel),
    .io_p(gen_p_i_57_io_p)
  );
  gen_p_i gen_p_i_58 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_58_io_x),
    .io_x_sub(gen_p_i_58_io_x_sub),
    .io_sel(gen_p_i_58_io_sel),
    .io_p(gen_p_i_58_io_p)
  );
  gen_p_i gen_p_i_59 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_59_io_x),
    .io_x_sub(gen_p_i_59_io_x_sub),
    .io_sel(gen_p_i_59_io_sel),
    .io_p(gen_p_i_59_io_p)
  );
  gen_p_i gen_p_i_60 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_60_io_x),
    .io_x_sub(gen_p_i_60_io_x_sub),
    .io_sel(gen_p_i_60_io_sel),
    .io_p(gen_p_i_60_io_p)
  );
  gen_p_i gen_p_i_61 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_61_io_x),
    .io_x_sub(gen_p_i_61_io_x_sub),
    .io_sel(gen_p_i_61_io_sel),
    .io_p(gen_p_i_61_io_p)
  );
  gen_p_i gen_p_i_62 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_62_io_x),
    .io_x_sub(gen_p_i_62_io_x_sub),
    .io_sel(gen_p_i_62_io_sel),
    .io_p(gen_p_i_62_io_p)
  );
  gen_p_i gen_p_i_63 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_63_io_x),
    .io_x_sub(gen_p_i_63_io_x_sub),
    .io_sel(gen_p_i_63_io_sel),
    .io_p(gen_p_i_63_io_p)
  );
  gen_p_i gen_p_i_64 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_64_io_x),
    .io_x_sub(gen_p_i_64_io_x_sub),
    .io_sel(gen_p_i_64_io_sel),
    .io_p(gen_p_i_64_io_p)
  );
  gen_p_i gen_p_i_65 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_65_io_x),
    .io_x_sub(gen_p_i_65_io_x_sub),
    .io_sel(gen_p_i_65_io_sel),
    .io_p(gen_p_i_65_io_p)
  );
  gen_p_i gen_p_i_66 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_66_io_x),
    .io_x_sub(gen_p_i_66_io_x_sub),
    .io_sel(gen_p_i_66_io_sel),
    .io_p(gen_p_i_66_io_p)
  );
  gen_p_i gen_p_i_67 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_67_io_x),
    .io_x_sub(gen_p_i_67_io_x_sub),
    .io_sel(gen_p_i_67_io_sel),
    .io_p(gen_p_i_67_io_p)
  );
  gen_p_i gen_p_i_68 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_68_io_x),
    .io_x_sub(gen_p_i_68_io_x_sub),
    .io_sel(gen_p_i_68_io_sel),
    .io_p(gen_p_i_68_io_p)
  );
  gen_p_i gen_p_i_69 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_69_io_x),
    .io_x_sub(gen_p_i_69_io_x_sub),
    .io_sel(gen_p_i_69_io_sel),
    .io_p(gen_p_i_69_io_p)
  );
  gen_p_i gen_p_i_70 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_70_io_x),
    .io_x_sub(gen_p_i_70_io_x_sub),
    .io_sel(gen_p_i_70_io_sel),
    .io_p(gen_p_i_70_io_p)
  );
  gen_p_i gen_p_i_71 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_71_io_x),
    .io_x_sub(gen_p_i_71_io_x_sub),
    .io_sel(gen_p_i_71_io_sel),
    .io_p(gen_p_i_71_io_p)
  );
  gen_p_i gen_p_i_72 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_72_io_x),
    .io_x_sub(gen_p_i_72_io_x_sub),
    .io_sel(gen_p_i_72_io_sel),
    .io_p(gen_p_i_72_io_p)
  );
  gen_p_i gen_p_i_73 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_73_io_x),
    .io_x_sub(gen_p_i_73_io_x_sub),
    .io_sel(gen_p_i_73_io_sel),
    .io_p(gen_p_i_73_io_p)
  );
  gen_p_i gen_p_i_74 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_74_io_x),
    .io_x_sub(gen_p_i_74_io_x_sub),
    .io_sel(gen_p_i_74_io_sel),
    .io_p(gen_p_i_74_io_p)
  );
  gen_p_i gen_p_i_75 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_75_io_x),
    .io_x_sub(gen_p_i_75_io_x_sub),
    .io_sel(gen_p_i_75_io_sel),
    .io_p(gen_p_i_75_io_p)
  );
  gen_p_i gen_p_i_76 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_76_io_x),
    .io_x_sub(gen_p_i_76_io_x_sub),
    .io_sel(gen_p_i_76_io_sel),
    .io_p(gen_p_i_76_io_p)
  );
  gen_p_i gen_p_i_77 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_77_io_x),
    .io_x_sub(gen_p_i_77_io_x_sub),
    .io_sel(gen_p_i_77_io_sel),
    .io_p(gen_p_i_77_io_p)
  );
  gen_p_i gen_p_i_78 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_78_io_x),
    .io_x_sub(gen_p_i_78_io_x_sub),
    .io_sel(gen_p_i_78_io_sel),
    .io_p(gen_p_i_78_io_p)
  );
  gen_p_i gen_p_i_79 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_79_io_x),
    .io_x_sub(gen_p_i_79_io_x_sub),
    .io_sel(gen_p_i_79_io_sel),
    .io_p(gen_p_i_79_io_p)
  );
  gen_p_i gen_p_i_80 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_80_io_x),
    .io_x_sub(gen_p_i_80_io_x_sub),
    .io_sel(gen_p_i_80_io_sel),
    .io_p(gen_p_i_80_io_p)
  );
  gen_p_i gen_p_i_81 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_81_io_x),
    .io_x_sub(gen_p_i_81_io_x_sub),
    .io_sel(gen_p_i_81_io_sel),
    .io_p(gen_p_i_81_io_p)
  );
  gen_p_i gen_p_i_82 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_82_io_x),
    .io_x_sub(gen_p_i_82_io_x_sub),
    .io_sel(gen_p_i_82_io_sel),
    .io_p(gen_p_i_82_io_p)
  );
  gen_p_i gen_p_i_83 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_83_io_x),
    .io_x_sub(gen_p_i_83_io_x_sub),
    .io_sel(gen_p_i_83_io_sel),
    .io_p(gen_p_i_83_io_p)
  );
  gen_p_i gen_p_i_84 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_84_io_x),
    .io_x_sub(gen_p_i_84_io_x_sub),
    .io_sel(gen_p_i_84_io_sel),
    .io_p(gen_p_i_84_io_p)
  );
  gen_p_i gen_p_i_85 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_85_io_x),
    .io_x_sub(gen_p_i_85_io_x_sub),
    .io_sel(gen_p_i_85_io_sel),
    .io_p(gen_p_i_85_io_p)
  );
  gen_p_i gen_p_i_86 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_86_io_x),
    .io_x_sub(gen_p_i_86_io_x_sub),
    .io_sel(gen_p_i_86_io_sel),
    .io_p(gen_p_i_86_io_p)
  );
  gen_p_i gen_p_i_87 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_87_io_x),
    .io_x_sub(gen_p_i_87_io_x_sub),
    .io_sel(gen_p_i_87_io_sel),
    .io_p(gen_p_i_87_io_p)
  );
  gen_p_i gen_p_i_88 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_88_io_x),
    .io_x_sub(gen_p_i_88_io_x_sub),
    .io_sel(gen_p_i_88_io_sel),
    .io_p(gen_p_i_88_io_p)
  );
  gen_p_i gen_p_i_89 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_89_io_x),
    .io_x_sub(gen_p_i_89_io_x_sub),
    .io_sel(gen_p_i_89_io_sel),
    .io_p(gen_p_i_89_io_p)
  );
  gen_p_i gen_p_i_90 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_90_io_x),
    .io_x_sub(gen_p_i_90_io_x_sub),
    .io_sel(gen_p_i_90_io_sel),
    .io_p(gen_p_i_90_io_p)
  );
  gen_p_i gen_p_i_91 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_91_io_x),
    .io_x_sub(gen_p_i_91_io_x_sub),
    .io_sel(gen_p_i_91_io_sel),
    .io_p(gen_p_i_91_io_p)
  );
  gen_p_i gen_p_i_92 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_92_io_x),
    .io_x_sub(gen_p_i_92_io_x_sub),
    .io_sel(gen_p_i_92_io_sel),
    .io_p(gen_p_i_92_io_p)
  );
  gen_p_i gen_p_i_93 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_93_io_x),
    .io_x_sub(gen_p_i_93_io_x_sub),
    .io_sel(gen_p_i_93_io_sel),
    .io_p(gen_p_i_93_io_p)
  );
  gen_p_i gen_p_i_94 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_94_io_x),
    .io_x_sub(gen_p_i_94_io_x_sub),
    .io_sel(gen_p_i_94_io_sel),
    .io_p(gen_p_i_94_io_p)
  );
  gen_p_i gen_p_i_95 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_95_io_x),
    .io_x_sub(gen_p_i_95_io_x_sub),
    .io_sel(gen_p_i_95_io_sel),
    .io_p(gen_p_i_95_io_p)
  );
  gen_p_i gen_p_i_96 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_96_io_x),
    .io_x_sub(gen_p_i_96_io_x_sub),
    .io_sel(gen_p_i_96_io_sel),
    .io_p(gen_p_i_96_io_p)
  );
  gen_p_i gen_p_i_97 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_97_io_x),
    .io_x_sub(gen_p_i_97_io_x_sub),
    .io_sel(gen_p_i_97_io_sel),
    .io_p(gen_p_i_97_io_p)
  );
  gen_p_i gen_p_i_98 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_98_io_x),
    .io_x_sub(gen_p_i_98_io_x_sub),
    .io_sel(gen_p_i_98_io_sel),
    .io_p(gen_p_i_98_io_p)
  );
  gen_p_i gen_p_i_99 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_99_io_x),
    .io_x_sub(gen_p_i_99_io_x_sub),
    .io_sel(gen_p_i_99_io_sel),
    .io_p(gen_p_i_99_io_p)
  );
  gen_p_i gen_p_i_100 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_100_io_x),
    .io_x_sub(gen_p_i_100_io_x_sub),
    .io_sel(gen_p_i_100_io_sel),
    .io_p(gen_p_i_100_io_p)
  );
  gen_p_i gen_p_i_101 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_101_io_x),
    .io_x_sub(gen_p_i_101_io_x_sub),
    .io_sel(gen_p_i_101_io_sel),
    .io_p(gen_p_i_101_io_p)
  );
  gen_p_i gen_p_i_102 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_102_io_x),
    .io_x_sub(gen_p_i_102_io_x_sub),
    .io_sel(gen_p_i_102_io_sel),
    .io_p(gen_p_i_102_io_p)
  );
  gen_p_i gen_p_i_103 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_103_io_x),
    .io_x_sub(gen_p_i_103_io_x_sub),
    .io_sel(gen_p_i_103_io_sel),
    .io_p(gen_p_i_103_io_p)
  );
  gen_p_i gen_p_i_104 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_104_io_x),
    .io_x_sub(gen_p_i_104_io_x_sub),
    .io_sel(gen_p_i_104_io_sel),
    .io_p(gen_p_i_104_io_p)
  );
  gen_p_i gen_p_i_105 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_105_io_x),
    .io_x_sub(gen_p_i_105_io_x_sub),
    .io_sel(gen_p_i_105_io_sel),
    .io_p(gen_p_i_105_io_p)
  );
  gen_p_i gen_p_i_106 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_106_io_x),
    .io_x_sub(gen_p_i_106_io_x_sub),
    .io_sel(gen_p_i_106_io_sel),
    .io_p(gen_p_i_106_io_p)
  );
  gen_p_i gen_p_i_107 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_107_io_x),
    .io_x_sub(gen_p_i_107_io_x_sub),
    .io_sel(gen_p_i_107_io_sel),
    .io_p(gen_p_i_107_io_p)
  );
  gen_p_i gen_p_i_108 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_108_io_x),
    .io_x_sub(gen_p_i_108_io_x_sub),
    .io_sel(gen_p_i_108_io_sel),
    .io_p(gen_p_i_108_io_p)
  );
  gen_p_i gen_p_i_109 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_109_io_x),
    .io_x_sub(gen_p_i_109_io_x_sub),
    .io_sel(gen_p_i_109_io_sel),
    .io_p(gen_p_i_109_io_p)
  );
  gen_p_i gen_p_i_110 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_110_io_x),
    .io_x_sub(gen_p_i_110_io_x_sub),
    .io_sel(gen_p_i_110_io_sel),
    .io_p(gen_p_i_110_io_p)
  );
  gen_p_i gen_p_i_111 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_111_io_x),
    .io_x_sub(gen_p_i_111_io_x_sub),
    .io_sel(gen_p_i_111_io_sel),
    .io_p(gen_p_i_111_io_p)
  );
  gen_p_i gen_p_i_112 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_112_io_x),
    .io_x_sub(gen_p_i_112_io_x_sub),
    .io_sel(gen_p_i_112_io_sel),
    .io_p(gen_p_i_112_io_p)
  );
  gen_p_i gen_p_i_113 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_113_io_x),
    .io_x_sub(gen_p_i_113_io_x_sub),
    .io_sel(gen_p_i_113_io_sel),
    .io_p(gen_p_i_113_io_p)
  );
  gen_p_i gen_p_i_114 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_114_io_x),
    .io_x_sub(gen_p_i_114_io_x_sub),
    .io_sel(gen_p_i_114_io_sel),
    .io_p(gen_p_i_114_io_p)
  );
  gen_p_i gen_p_i_115 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_115_io_x),
    .io_x_sub(gen_p_i_115_io_x_sub),
    .io_sel(gen_p_i_115_io_sel),
    .io_p(gen_p_i_115_io_p)
  );
  gen_p_i gen_p_i_116 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_116_io_x),
    .io_x_sub(gen_p_i_116_io_x_sub),
    .io_sel(gen_p_i_116_io_sel),
    .io_p(gen_p_i_116_io_p)
  );
  gen_p_i gen_p_i_117 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_117_io_x),
    .io_x_sub(gen_p_i_117_io_x_sub),
    .io_sel(gen_p_i_117_io_sel),
    .io_p(gen_p_i_117_io_p)
  );
  gen_p_i gen_p_i_118 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_118_io_x),
    .io_x_sub(gen_p_i_118_io_x_sub),
    .io_sel(gen_p_i_118_io_sel),
    .io_p(gen_p_i_118_io_p)
  );
  gen_p_i gen_p_i_119 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_119_io_x),
    .io_x_sub(gen_p_i_119_io_x_sub),
    .io_sel(gen_p_i_119_io_sel),
    .io_p(gen_p_i_119_io_p)
  );
  gen_p_i gen_p_i_120 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_120_io_x),
    .io_x_sub(gen_p_i_120_io_x_sub),
    .io_sel(gen_p_i_120_io_sel),
    .io_p(gen_p_i_120_io_p)
  );
  gen_p_i gen_p_i_121 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_121_io_x),
    .io_x_sub(gen_p_i_121_io_x_sub),
    .io_sel(gen_p_i_121_io_sel),
    .io_p(gen_p_i_121_io_p)
  );
  gen_p_i gen_p_i_122 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_122_io_x),
    .io_x_sub(gen_p_i_122_io_x_sub),
    .io_sel(gen_p_i_122_io_sel),
    .io_p(gen_p_i_122_io_p)
  );
  gen_p_i gen_p_i_123 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_123_io_x),
    .io_x_sub(gen_p_i_123_io_x_sub),
    .io_sel(gen_p_i_123_io_sel),
    .io_p(gen_p_i_123_io_p)
  );
  gen_p_i gen_p_i_124 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_124_io_x),
    .io_x_sub(gen_p_i_124_io_x_sub),
    .io_sel(gen_p_i_124_io_sel),
    .io_p(gen_p_i_124_io_p)
  );
  gen_p_i gen_p_i_125 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_125_io_x),
    .io_x_sub(gen_p_i_125_io_x_sub),
    .io_sel(gen_p_i_125_io_sel),
    .io_p(gen_p_i_125_io_p)
  );
  gen_p_i gen_p_i_126 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_126_io_x),
    .io_x_sub(gen_p_i_126_io_x_sub),
    .io_sel(gen_p_i_126_io_sel),
    .io_p(gen_p_i_126_io_p)
  );
  gen_p_i gen_p_i_127 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_127_io_x),
    .io_x_sub(gen_p_i_127_io_x_sub),
    .io_sel(gen_p_i_127_io_sel),
    .io_p(gen_p_i_127_io_p)
  );
  gen_p_i gen_p_i_128 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_128_io_x),
    .io_x_sub(gen_p_i_128_io_x_sub),
    .io_sel(gen_p_i_128_io_sel),
    .io_p(gen_p_i_128_io_p)
  );
  gen_p_i gen_p_i_129 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_129_io_x),
    .io_x_sub(gen_p_i_129_io_x_sub),
    .io_sel(gen_p_i_129_io_sel),
    .io_p(gen_p_i_129_io_p)
  );
  gen_p_i gen_p_i_130 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_130_io_x),
    .io_x_sub(gen_p_i_130_io_x_sub),
    .io_sel(gen_p_i_130_io_sel),
    .io_p(gen_p_i_130_io_p)
  );
  gen_p_i gen_p_i_131 ( // @[wallace_mul.scala 72:29]
    .io_x(gen_p_i_131_io_x),
    .io_x_sub(gen_p_i_131_io_x_sub),
    .io_sel(gen_p_i_131_io_sel),
    .io_p(gen_p_i_131_io_p)
  );
  assign io_p = {io_p_hi,io_p_lo}; // @[Cat.scala 33:92]
  assign io_c = gen_sel_io_out[0] | gen_sel_io_out[2]; // @[wallace_mul.scala 88:21]
  assign gen_sel_io_src = io_src; // @[wallace_mul.scala 74:10]
  assign gen_p_i_io_x = io_x[0]; // @[wallace_mul.scala 76:16]
  assign gen_p_i_io_x_sub = 1'h0; // @[wallace_mul.scala 77:14]
  assign gen_p_i_io_sel = gen_sel_io_out; // @[wallace_mul.scala 78:11]
  assign gen_p_i_1_io_x = io_x[1]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_1_io_x_sub = io_x[0]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_1_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_2_io_x = io_x[2]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_2_io_x_sub = io_x[1]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_2_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_3_io_x = io_x[3]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_3_io_x_sub = io_x[2]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_3_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_4_io_x = io_x[4]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_4_io_x_sub = io_x[3]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_4_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_5_io_x = io_x[5]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_5_io_x_sub = io_x[4]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_5_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_6_io_x = io_x[6]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_6_io_x_sub = io_x[5]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_6_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_7_io_x = io_x[7]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_7_io_x_sub = io_x[6]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_7_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_8_io_x = io_x[8]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_8_io_x_sub = io_x[7]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_8_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_9_io_x = io_x[9]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_9_io_x_sub = io_x[8]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_9_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_10_io_x = io_x[10]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_10_io_x_sub = io_x[9]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_10_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_11_io_x = io_x[11]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_11_io_x_sub = io_x[10]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_11_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_12_io_x = io_x[12]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_12_io_x_sub = io_x[11]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_12_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_13_io_x = io_x[13]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_13_io_x_sub = io_x[12]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_13_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_14_io_x = io_x[14]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_14_io_x_sub = io_x[13]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_14_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_15_io_x = io_x[15]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_15_io_x_sub = io_x[14]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_15_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_16_io_x = io_x[16]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_16_io_x_sub = io_x[15]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_16_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_17_io_x = io_x[17]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_17_io_x_sub = io_x[16]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_17_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_18_io_x = io_x[18]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_18_io_x_sub = io_x[17]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_18_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_19_io_x = io_x[19]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_19_io_x_sub = io_x[18]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_19_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_20_io_x = io_x[20]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_20_io_x_sub = io_x[19]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_20_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_21_io_x = io_x[21]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_21_io_x_sub = io_x[20]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_21_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_22_io_x = io_x[22]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_22_io_x_sub = io_x[21]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_22_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_23_io_x = io_x[23]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_23_io_x_sub = io_x[22]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_23_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_24_io_x = io_x[24]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_24_io_x_sub = io_x[23]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_24_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_25_io_x = io_x[25]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_25_io_x_sub = io_x[24]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_25_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_26_io_x = io_x[26]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_26_io_x_sub = io_x[25]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_26_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_27_io_x = io_x[27]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_27_io_x_sub = io_x[26]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_27_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_28_io_x = io_x[28]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_28_io_x_sub = io_x[27]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_28_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_29_io_x = io_x[29]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_29_io_x_sub = io_x[28]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_29_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_30_io_x = io_x[30]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_30_io_x_sub = io_x[29]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_30_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_31_io_x = io_x[31]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_31_io_x_sub = io_x[30]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_31_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_32_io_x = io_x[32]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_32_io_x_sub = io_x[31]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_32_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_33_io_x = io_x[33]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_33_io_x_sub = io_x[32]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_33_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_34_io_x = io_x[34]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_34_io_x_sub = io_x[33]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_34_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_35_io_x = io_x[35]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_35_io_x_sub = io_x[34]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_35_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_36_io_x = io_x[36]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_36_io_x_sub = io_x[35]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_36_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_37_io_x = io_x[37]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_37_io_x_sub = io_x[36]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_37_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_38_io_x = io_x[38]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_38_io_x_sub = io_x[37]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_38_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_39_io_x = io_x[39]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_39_io_x_sub = io_x[38]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_39_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_40_io_x = io_x[40]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_40_io_x_sub = io_x[39]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_40_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_41_io_x = io_x[41]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_41_io_x_sub = io_x[40]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_41_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_42_io_x = io_x[42]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_42_io_x_sub = io_x[41]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_42_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_43_io_x = io_x[43]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_43_io_x_sub = io_x[42]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_43_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_44_io_x = io_x[44]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_44_io_x_sub = io_x[43]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_44_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_45_io_x = io_x[45]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_45_io_x_sub = io_x[44]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_45_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_46_io_x = io_x[46]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_46_io_x_sub = io_x[45]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_46_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_47_io_x = io_x[47]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_47_io_x_sub = io_x[46]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_47_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_48_io_x = io_x[48]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_48_io_x_sub = io_x[47]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_48_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_49_io_x = io_x[49]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_49_io_x_sub = io_x[48]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_49_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_50_io_x = io_x[50]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_50_io_x_sub = io_x[49]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_50_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_51_io_x = io_x[51]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_51_io_x_sub = io_x[50]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_51_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_52_io_x = io_x[52]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_52_io_x_sub = io_x[51]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_52_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_53_io_x = io_x[53]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_53_io_x_sub = io_x[52]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_53_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_54_io_x = io_x[54]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_54_io_x_sub = io_x[53]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_54_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_55_io_x = io_x[55]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_55_io_x_sub = io_x[54]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_55_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_56_io_x = io_x[56]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_56_io_x_sub = io_x[55]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_56_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_57_io_x = io_x[57]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_57_io_x_sub = io_x[56]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_57_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_58_io_x = io_x[58]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_58_io_x_sub = io_x[57]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_58_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_59_io_x = io_x[59]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_59_io_x_sub = io_x[58]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_59_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_60_io_x = io_x[60]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_60_io_x_sub = io_x[59]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_60_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_61_io_x = io_x[61]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_61_io_x_sub = io_x[60]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_61_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_62_io_x = io_x[62]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_62_io_x_sub = io_x[61]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_62_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_63_io_x = io_x[63]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_63_io_x_sub = io_x[62]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_63_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_64_io_x = io_x[64]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_64_io_x_sub = io_x[63]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_64_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_65_io_x = io_x[65]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_65_io_x_sub = io_x[64]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_65_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_66_io_x = io_x[66]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_66_io_x_sub = io_x[65]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_66_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_67_io_x = io_x[67]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_67_io_x_sub = io_x[66]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_67_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_68_io_x = io_x[68]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_68_io_x_sub = io_x[67]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_68_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_69_io_x = io_x[69]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_69_io_x_sub = io_x[68]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_69_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_70_io_x = io_x[70]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_70_io_x_sub = io_x[69]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_70_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_71_io_x = io_x[71]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_71_io_x_sub = io_x[70]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_71_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_72_io_x = io_x[72]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_72_io_x_sub = io_x[71]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_72_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_73_io_x = io_x[73]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_73_io_x_sub = io_x[72]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_73_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_74_io_x = io_x[74]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_74_io_x_sub = io_x[73]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_74_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_75_io_x = io_x[75]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_75_io_x_sub = io_x[74]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_75_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_76_io_x = io_x[76]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_76_io_x_sub = io_x[75]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_76_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_77_io_x = io_x[77]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_77_io_x_sub = io_x[76]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_77_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_78_io_x = io_x[78]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_78_io_x_sub = io_x[77]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_78_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_79_io_x = io_x[79]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_79_io_x_sub = io_x[78]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_79_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_80_io_x = io_x[80]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_80_io_x_sub = io_x[79]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_80_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_81_io_x = io_x[81]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_81_io_x_sub = io_x[80]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_81_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_82_io_x = io_x[82]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_82_io_x_sub = io_x[81]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_82_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_83_io_x = io_x[83]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_83_io_x_sub = io_x[82]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_83_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_84_io_x = io_x[84]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_84_io_x_sub = io_x[83]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_84_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_85_io_x = io_x[85]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_85_io_x_sub = io_x[84]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_85_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_86_io_x = io_x[86]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_86_io_x_sub = io_x[85]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_86_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_87_io_x = io_x[87]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_87_io_x_sub = io_x[86]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_87_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_88_io_x = io_x[88]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_88_io_x_sub = io_x[87]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_88_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_89_io_x = io_x[89]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_89_io_x_sub = io_x[88]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_89_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_90_io_x = io_x[90]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_90_io_x_sub = io_x[89]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_90_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_91_io_x = io_x[91]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_91_io_x_sub = io_x[90]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_91_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_92_io_x = io_x[92]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_92_io_x_sub = io_x[91]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_92_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_93_io_x = io_x[93]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_93_io_x_sub = io_x[92]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_93_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_94_io_x = io_x[94]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_94_io_x_sub = io_x[93]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_94_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_95_io_x = io_x[95]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_95_io_x_sub = io_x[94]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_95_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_96_io_x = io_x[96]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_96_io_x_sub = io_x[95]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_96_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_97_io_x = io_x[97]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_97_io_x_sub = io_x[96]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_97_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_98_io_x = io_x[98]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_98_io_x_sub = io_x[97]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_98_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_99_io_x = io_x[99]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_99_io_x_sub = io_x[98]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_99_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_100_io_x = io_x[100]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_100_io_x_sub = io_x[99]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_100_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_101_io_x = io_x[101]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_101_io_x_sub = io_x[100]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_101_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_102_io_x = io_x[102]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_102_io_x_sub = io_x[101]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_102_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_103_io_x = io_x[103]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_103_io_x_sub = io_x[102]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_103_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_104_io_x = io_x[104]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_104_io_x_sub = io_x[103]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_104_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_105_io_x = io_x[105]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_105_io_x_sub = io_x[104]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_105_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_106_io_x = io_x[106]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_106_io_x_sub = io_x[105]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_106_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_107_io_x = io_x[107]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_107_io_x_sub = io_x[106]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_107_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_108_io_x = io_x[108]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_108_io_x_sub = io_x[107]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_108_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_109_io_x = io_x[109]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_109_io_x_sub = io_x[108]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_109_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_110_io_x = io_x[110]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_110_io_x_sub = io_x[109]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_110_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_111_io_x = io_x[111]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_111_io_x_sub = io_x[110]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_111_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_112_io_x = io_x[112]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_112_io_x_sub = io_x[111]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_112_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_113_io_x = io_x[113]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_113_io_x_sub = io_x[112]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_113_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_114_io_x = io_x[114]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_114_io_x_sub = io_x[113]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_114_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_115_io_x = io_x[115]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_115_io_x_sub = io_x[114]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_115_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_116_io_x = io_x[116]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_116_io_x_sub = io_x[115]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_116_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_117_io_x = io_x[117]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_117_io_x_sub = io_x[116]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_117_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_118_io_x = io_x[118]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_118_io_x_sub = io_x[117]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_118_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_119_io_x = io_x[119]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_119_io_x_sub = io_x[118]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_119_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_120_io_x = io_x[120]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_120_io_x_sub = io_x[119]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_120_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_121_io_x = io_x[121]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_121_io_x_sub = io_x[120]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_121_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_122_io_x = io_x[122]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_122_io_x_sub = io_x[121]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_122_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_123_io_x = io_x[123]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_123_io_x_sub = io_x[122]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_123_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_124_io_x = io_x[124]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_124_io_x_sub = io_x[123]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_124_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_125_io_x = io_x[125]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_125_io_x_sub = io_x[124]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_125_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_126_io_x = io_x[126]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_126_io_x_sub = io_x[125]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_126_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_127_io_x = io_x[127]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_127_io_x_sub = io_x[126]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_127_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_128_io_x = io_x[128]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_128_io_x_sub = io_x[127]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_128_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_129_io_x = io_x[129]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_129_io_x_sub = io_x[128]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_129_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_130_io_x = io_x[130]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_130_io_x_sub = io_x[129]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_130_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
  assign gen_p_i_131_io_x = io_x[131]; // @[wallace_mul.scala 81:18]
  assign gen_p_i_131_io_x_sub = io_x[130]; // @[wallace_mul.scala 82:23]
  assign gen_p_i_131_io_sel = gen_sel_io_out; // @[wallace_mul.scala 83:13]
endmodule
