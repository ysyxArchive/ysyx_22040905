module ps2_keyboard(
  input        clock,
  input        io_ps2_clk,
  input        io_ps2_data,
  input        io_nextdata_n,
  output [7:0] io_data,
  output       io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg  rea; // @[ps2.scala 144:16]
  reg  buffer_0; // @[ps2.scala 152:19]
  reg  buffer_1; // @[ps2.scala 152:19]
  reg  buffer_2; // @[ps2.scala 152:19]
  reg  buffer_3; // @[ps2.scala 152:19]
  reg  buffer_4; // @[ps2.scala 152:19]
  reg  buffer_5; // @[ps2.scala 152:19]
  reg  buffer_6; // @[ps2.scala 152:19]
  reg  buffer_7; // @[ps2.scala 152:19]
  reg  buffer_8; // @[ps2.scala 152:19]
  reg  buffer_9; // @[ps2.scala 152:19]
  reg [7:0] fifo_0; // @[ps2.scala 153:17]
  reg [7:0] fifo_1; // @[ps2.scala 153:17]
  reg [7:0] fifo_2; // @[ps2.scala 153:17]
  reg [7:0] fifo_3; // @[ps2.scala 153:17]
  reg [7:0] fifo_4; // @[ps2.scala 153:17]
  reg [7:0] fifo_5; // @[ps2.scala 153:17]
  reg [7:0] fifo_6; // @[ps2.scala 153:17]
  reg [7:0] fifo_7; // @[ps2.scala 153:17]
  reg [2:0] w_ptr; // @[ps2.scala 154:18]
  reg [2:0] r_ptr; // @[ps2.scala 155:18]
  reg [3:0] count; // @[ps2.scala 156:18]
  reg [2:0] ps2_clk_sync; // @[ps2.scala 157:25]
  wire [1:0] ps2_clk_sync_hi = ps2_clk_sync[1:0]; // @[ps2.scala 159:35]
  wire  sampling = ps2_clk_sync[2] & ~ps2_clk_sync[1]; // @[ps2.scala 161:30]
  wire [2:0] _r_ptr_T_1 = r_ptr + 3'h1; // @[ps2.scala 171:29]
  wire  _GEN_0 = w_ptr == _r_ptr_T_1 ? 1'h0 : rea; // @[ps2.scala 172:42 ps2.scala 173:24 ps2.scala 144:16]
  wire  _GEN_3 = ~io_nextdata_n ? _GEN_0 : rea; // @[ps2.scala 170:38 ps2.scala 144:16]
  wire  _GEN_6 = rea ? _GEN_3 : rea; // @[ps2.scala 169:24 ps2.scala 144:16]
  wire [7:0] _fifo_T = {buffer_8,buffer_7,buffer_6,buffer_5,buffer_4,buffer_3,buffer_2,buffer_1}; // @[Cat.scala 30:58]
  wire [2:0] _w_ptr_T_1 = w_ptr + 3'h1; // @[ps2.scala 182:33]
  wire  _GEN_25 = ~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3
     ^ buffer_2 ^ buffer_1) | _GEN_6; // @[ps2.scala 180:162 ps2.scala 183:24]
  wire [3:0] _count_T_1 = count + 4'h1; // @[ps2.scala 189:29]
  wire [7:0] _GEN_106 = 3'h1 == r_ptr ? fifo_1 : fifo_0; // @[ps2.scala 193:12 ps2.scala 193:12]
  wire [7:0] _GEN_107 = 3'h2 == r_ptr ? fifo_2 : _GEN_106; // @[ps2.scala 193:12 ps2.scala 193:12]
  wire [7:0] _GEN_108 = 3'h3 == r_ptr ? fifo_3 : _GEN_107; // @[ps2.scala 193:12 ps2.scala 193:12]
  wire [7:0] _GEN_109 = 3'h4 == r_ptr ? fifo_4 : _GEN_108; // @[ps2.scala 193:12 ps2.scala 193:12]
  wire [7:0] _GEN_110 = 3'h5 == r_ptr ? fifo_5 : _GEN_109; // @[ps2.scala 193:12 ps2.scala 193:12]
  wire [7:0] _GEN_111 = 3'h6 == r_ptr ? fifo_6 : _GEN_110; // @[ps2.scala 193:12 ps2.scala 193:12]
  assign io_data = 3'h7 == r_ptr ? fifo_7 : _GEN_111; // @[ps2.scala 193:12 ps2.scala 193:12]
  assign io_ready = rea; // @[ps2.scala 162:24 ps2.scala 150:13]
  always @(posedge clock) begin
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        rea <= _GEN_25;
      end else begin
        rea <= _GEN_6;
      end
    end else begin
      rea <= _GEN_6;
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h0 == count) begin // @[ps2.scala 188:30]
          buffer_0 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h1 == count) begin // @[ps2.scala 188:30]
          buffer_1 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h2 == count) begin // @[ps2.scala 188:30]
          buffer_2 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h3 == count) begin // @[ps2.scala 188:30]
          buffer_3 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h4 == count) begin // @[ps2.scala 188:30]
          buffer_4 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h5 == count) begin // @[ps2.scala 188:30]
          buffer_5 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h6 == count) begin // @[ps2.scala 188:30]
          buffer_6 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h7 == count) begin // @[ps2.scala 188:30]
          buffer_7 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h8 == count) begin // @[ps2.scala 188:30]
          buffer_8 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 179:31]
        if (4'h9 == count) begin // @[ps2.scala 188:30]
          buffer_9 <= io_ps2_data; // @[ps2.scala 188:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h0 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_0 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h1 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_1 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h2 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_2 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h3 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_3 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h4 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_4 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h5 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_5 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h6 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_6 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          if (3'h7 == w_ptr) begin // @[ps2.scala 181:32]
            fifo_7 <= _fifo_T; // @[ps2.scala 181:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 180:162]
          w_ptr <= _w_ptr_T_1; // @[ps2.scala 182:26]
        end
      end
    end
    if (rea) begin // @[ps2.scala 169:24]
      if (~io_nextdata_n) begin // @[ps2.scala 170:38]
        r_ptr <= _r_ptr_T_1; // @[ps2.scala 171:22]
      end
    end
    if (sampling) begin // @[ps2.scala 178:29]
      if (count == 4'ha) begin // @[ps2.scala 179:31]
        count <= 4'h0; // @[ps2.scala 186:22]
      end else begin
        count <= _count_T_1; // @[ps2.scala 189:22]
      end
    end
    ps2_clk_sync <= {ps2_clk_sync_hi,io_ps2_clk}; // @[Cat.scala 30:58]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rea = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  fifo_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  fifo_1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  fifo_2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  fifo_3 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  fifo_4 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  fifo_5 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  fifo_6 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  fifo_7 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  w_ptr = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  r_ptr = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  count = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  ps2_clk_sync = _RAND_22[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ps2ascii(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [255:0] _RAND_0;
  reg [255:0] _RAND_1;
  reg [255:0] _RAND_2;
  reg [255:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [255:0] _RAND_5;
  reg [255:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [255:0] _RAND_9;
  reg [255:0] _RAND_10;
  reg [255:0] _RAND_11;
  reg [255:0] _RAND_12;
  reg [255:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [255:0] _RAND_15;
  reg [255:0] _RAND_16;
  reg [255:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [255:0] _RAND_19;
  reg [255:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [255:0] _RAND_22;
  reg [255:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [255:0] _RAND_25;
  reg [255:0] _RAND_26;
  reg [255:0] _RAND_27;
  reg [255:0] _RAND_28;
  reg [255:0] _RAND_29;
  reg [255:0] _RAND_30;
  reg [255:0] _RAND_31;
  reg [255:0] _RAND_32;
  reg [255:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [255:0] _RAND_35;
  reg [255:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  reg [255:0] table_21; // @[ps2.scala 201:22]
  reg [255:0] table_22; // @[ps2.scala 201:22]
  reg [255:0] table_26; // @[ps2.scala 201:22]
  reg [255:0] table_27; // @[ps2.scala 201:22]
  reg [255:0] table_28; // @[ps2.scala 201:22]
  reg [255:0] table_29; // @[ps2.scala 201:22]
  reg [255:0] table_30; // @[ps2.scala 201:22]
  reg [255:0] table_33; // @[ps2.scala 201:22]
  reg [255:0] table_34; // @[ps2.scala 201:22]
  reg [255:0] table_35; // @[ps2.scala 201:22]
  reg [255:0] table_36; // @[ps2.scala 201:22]
  reg [255:0] table_37; // @[ps2.scala 201:22]
  reg [255:0] table_38; // @[ps2.scala 201:22]
  reg [255:0] table_42; // @[ps2.scala 201:22]
  reg [255:0] table_43; // @[ps2.scala 201:22]
  reg [255:0] table_44; // @[ps2.scala 201:22]
  reg [255:0] table_45; // @[ps2.scala 201:22]
  reg [255:0] table_46; // @[ps2.scala 201:22]
  reg [255:0] table_49; // @[ps2.scala 201:22]
  reg [255:0] table_50; // @[ps2.scala 201:22]
  reg [255:0] table_51; // @[ps2.scala 201:22]
  reg [255:0] table_52; // @[ps2.scala 201:22]
  reg [255:0] table_53; // @[ps2.scala 201:22]
  reg [255:0] table_54; // @[ps2.scala 201:22]
  reg [255:0] table_58; // @[ps2.scala 201:22]
  reg [255:0] table_59; // @[ps2.scala 201:22]
  reg [255:0] table_60; // @[ps2.scala 201:22]
  reg [255:0] table_61; // @[ps2.scala 201:22]
  reg [255:0] table_62; // @[ps2.scala 201:22]
  reg [255:0] table_66; // @[ps2.scala 201:22]
  reg [255:0] table_67; // @[ps2.scala 201:22]
  reg [255:0] table_68; // @[ps2.scala 201:22]
  reg [255:0] table_69; // @[ps2.scala 201:22]
  reg [255:0] table_70; // @[ps2.scala 201:22]
  reg [255:0] table_75; // @[ps2.scala 201:22]
  reg [255:0] table_77; // @[ps2.scala 201:22]
  reg [255:0] table_90; // @[ps2.scala 201:22]
  wire [255:0] _GEN_21 = 8'h15 == io_in ? table_21 : 256'h0; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_22 = 8'h16 == io_in ? table_22 : _GEN_21; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_23 = 8'h17 == io_in ? 256'h0 : _GEN_22; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_24 = 8'h18 == io_in ? 256'h0 : _GEN_23; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_25 = 8'h19 == io_in ? 256'h0 : _GEN_24; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_26 = 8'h1a == io_in ? table_26 : _GEN_25; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_27 = 8'h1b == io_in ? table_27 : _GEN_26; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_28 = 8'h1c == io_in ? table_28 : _GEN_27; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_29 = 8'h1d == io_in ? table_29 : _GEN_28; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_30 = 8'h1e == io_in ? table_30 : _GEN_29; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_31 = 8'h1f == io_in ? 256'h0 : _GEN_30; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_32 = 8'h20 == io_in ? 256'h0 : _GEN_31; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_33 = 8'h21 == io_in ? table_33 : _GEN_32; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_34 = 8'h22 == io_in ? table_34 : _GEN_33; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_35 = 8'h23 == io_in ? table_35 : _GEN_34; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_36 = 8'h24 == io_in ? table_36 : _GEN_35; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_37 = 8'h25 == io_in ? table_37 : _GEN_36; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_38 = 8'h26 == io_in ? table_38 : _GEN_37; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_39 = 8'h27 == io_in ? 256'h0 : _GEN_38; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_40 = 8'h28 == io_in ? 256'h0 : _GEN_39; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_41 = 8'h29 == io_in ? 256'h0 : _GEN_40; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_42 = 8'h2a == io_in ? table_42 : _GEN_41; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_43 = 8'h2b == io_in ? table_43 : _GEN_42; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_44 = 8'h2c == io_in ? table_44 : _GEN_43; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_45 = 8'h2d == io_in ? table_45 : _GEN_44; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_46 = 8'h2e == io_in ? table_46 : _GEN_45; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_47 = 8'h2f == io_in ? 256'h0 : _GEN_46; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_48 = 8'h30 == io_in ? 256'h0 : _GEN_47; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_49 = 8'h31 == io_in ? table_49 : _GEN_48; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_50 = 8'h32 == io_in ? table_50 : _GEN_49; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_51 = 8'h33 == io_in ? table_51 : _GEN_50; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_52 = 8'h34 == io_in ? table_52 : _GEN_51; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_53 = 8'h35 == io_in ? table_53 : _GEN_52; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_54 = 8'h36 == io_in ? table_54 : _GEN_53; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_55 = 8'h37 == io_in ? 256'h0 : _GEN_54; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_56 = 8'h38 == io_in ? 256'h0 : _GEN_55; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_57 = 8'h39 == io_in ? 256'h0 : _GEN_56; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_58 = 8'h3a == io_in ? table_58 : _GEN_57; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_59 = 8'h3b == io_in ? table_59 : _GEN_58; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_60 = 8'h3c == io_in ? table_60 : _GEN_59; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_61 = 8'h3d == io_in ? table_61 : _GEN_60; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_62 = 8'h3e == io_in ? table_62 : _GEN_61; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_63 = 8'h3f == io_in ? 256'h0 : _GEN_62; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_64 = 8'h40 == io_in ? 256'h0 : _GEN_63; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_65 = 8'h41 == io_in ? 256'h0 : _GEN_64; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_66 = 8'h42 == io_in ? table_66 : _GEN_65; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_67 = 8'h43 == io_in ? table_67 : _GEN_66; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_68 = 8'h44 == io_in ? table_68 : _GEN_67; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_69 = 8'h45 == io_in ? table_69 : _GEN_68; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_70 = 8'h46 == io_in ? table_70 : _GEN_69; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_71 = 8'h47 == io_in ? 256'h0 : _GEN_70; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_72 = 8'h48 == io_in ? 256'h0 : _GEN_71; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_73 = 8'h49 == io_in ? 256'h0 : _GEN_72; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_74 = 8'h4a == io_in ? 256'h0 : _GEN_73; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_75 = 8'h4b == io_in ? table_75 : _GEN_74; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_76 = 8'h4c == io_in ? 256'h0 : _GEN_75; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_77 = 8'h4d == io_in ? table_77 : _GEN_76; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_78 = 8'h4e == io_in ? 256'h0 : _GEN_77; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_79 = 8'h4f == io_in ? 256'h0 : _GEN_78; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_80 = 8'h50 == io_in ? 256'h0 : _GEN_79; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_81 = 8'h51 == io_in ? 256'h0 : _GEN_80; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_82 = 8'h52 == io_in ? 256'h0 : _GEN_81; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_83 = 8'h53 == io_in ? 256'h0 : _GEN_82; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_84 = 8'h54 == io_in ? 256'h0 : _GEN_83; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_85 = 8'h55 == io_in ? 256'h0 : _GEN_84; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_86 = 8'h56 == io_in ? 256'h0 : _GEN_85; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_87 = 8'h57 == io_in ? 256'h0 : _GEN_86; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_88 = 8'h58 == io_in ? 256'h0 : _GEN_87; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_89 = 8'h59 == io_in ? 256'h0 : _GEN_88; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_90 = 8'h5a == io_in ? table_90 : _GEN_89; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_91 = 8'h5b == io_in ? 256'h0 : _GEN_90; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_92 = 8'h5c == io_in ? 256'h0 : _GEN_91; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_93 = 8'h5d == io_in ? 256'h0 : _GEN_92; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_94 = 8'h5e == io_in ? 256'h0 : _GEN_93; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_95 = 8'h5f == io_in ? 256'h0 : _GEN_94; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_96 = 8'h60 == io_in ? 256'h0 : _GEN_95; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_97 = 8'h61 == io_in ? 256'h0 : _GEN_96; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_98 = 8'h62 == io_in ? 256'h0 : _GEN_97; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_99 = 8'h63 == io_in ? 256'h0 : _GEN_98; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_100 = 8'h64 == io_in ? 256'h0 : _GEN_99; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_101 = 8'h65 == io_in ? 256'h0 : _GEN_100; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_102 = 8'h66 == io_in ? 256'h0 : _GEN_101; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_103 = 8'h67 == io_in ? 256'h0 : _GEN_102; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_104 = 8'h68 == io_in ? 256'h0 : _GEN_103; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_105 = 8'h69 == io_in ? 256'h0 : _GEN_104; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_106 = 8'h6a == io_in ? 256'h0 : _GEN_105; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_107 = 8'h6b == io_in ? 256'h0 : _GEN_106; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_108 = 8'h6c == io_in ? 256'h0 : _GEN_107; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_109 = 8'h6d == io_in ? 256'h0 : _GEN_108; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_110 = 8'h6e == io_in ? 256'h0 : _GEN_109; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_111 = 8'h6f == io_in ? 256'h0 : _GEN_110; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_112 = 8'h70 == io_in ? 256'h0 : _GEN_111; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_113 = 8'h71 == io_in ? 256'h0 : _GEN_112; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_114 = 8'h72 == io_in ? 256'h0 : _GEN_113; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_115 = 8'h73 == io_in ? 256'h0 : _GEN_114; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_116 = 8'h74 == io_in ? 256'h0 : _GEN_115; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_117 = 8'h75 == io_in ? 256'h0 : _GEN_116; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_118 = 8'h76 == io_in ? 256'h0 : _GEN_117; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_119 = 8'h77 == io_in ? 256'h0 : _GEN_118; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_120 = 8'h78 == io_in ? 256'h0 : _GEN_119; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_121 = 8'h79 == io_in ? 256'h0 : _GEN_120; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_122 = 8'h7a == io_in ? 256'h0 : _GEN_121; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_123 = 8'h7b == io_in ? 256'h0 : _GEN_122; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_124 = 8'h7c == io_in ? 256'h0 : _GEN_123; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_125 = 8'h7d == io_in ? 256'h0 : _GEN_124; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_126 = 8'h7e == io_in ? 256'h0 : _GEN_125; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_127 = 8'h7f == io_in ? 256'h0 : _GEN_126; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_128 = 8'h80 == io_in ? 256'h0 : _GEN_127; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_129 = 8'h81 == io_in ? 256'h0 : _GEN_128; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_130 = 8'h82 == io_in ? 256'h0 : _GEN_129; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_131 = 8'h83 == io_in ? 256'h0 : _GEN_130; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_132 = 8'h84 == io_in ? 256'h0 : _GEN_131; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_133 = 8'h85 == io_in ? 256'h0 : _GEN_132; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_134 = 8'h86 == io_in ? 256'h0 : _GEN_133; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_135 = 8'h87 == io_in ? 256'h0 : _GEN_134; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_136 = 8'h88 == io_in ? 256'h0 : _GEN_135; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_137 = 8'h89 == io_in ? 256'h0 : _GEN_136; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_138 = 8'h8a == io_in ? 256'h0 : _GEN_137; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_139 = 8'h8b == io_in ? 256'h0 : _GEN_138; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_140 = 8'h8c == io_in ? 256'h0 : _GEN_139; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_141 = 8'h8d == io_in ? 256'h0 : _GEN_140; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_142 = 8'h8e == io_in ? 256'h0 : _GEN_141; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_143 = 8'h8f == io_in ? 256'h0 : _GEN_142; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_144 = 8'h90 == io_in ? 256'h0 : _GEN_143; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_145 = 8'h91 == io_in ? 256'h0 : _GEN_144; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_146 = 8'h92 == io_in ? 256'h0 : _GEN_145; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_147 = 8'h93 == io_in ? 256'h0 : _GEN_146; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_148 = 8'h94 == io_in ? 256'h0 : _GEN_147; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_149 = 8'h95 == io_in ? 256'h0 : _GEN_148; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_150 = 8'h96 == io_in ? 256'h0 : _GEN_149; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_151 = 8'h97 == io_in ? 256'h0 : _GEN_150; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_152 = 8'h98 == io_in ? 256'h0 : _GEN_151; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_153 = 8'h99 == io_in ? 256'h0 : _GEN_152; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_154 = 8'h9a == io_in ? 256'h0 : _GEN_153; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_155 = 8'h9b == io_in ? 256'h0 : _GEN_154; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_156 = 8'h9c == io_in ? 256'h0 : _GEN_155; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_157 = 8'h9d == io_in ? 256'h0 : _GEN_156; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_158 = 8'h9e == io_in ? 256'h0 : _GEN_157; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_159 = 8'h9f == io_in ? 256'h0 : _GEN_158; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_160 = 8'ha0 == io_in ? 256'h0 : _GEN_159; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_161 = 8'ha1 == io_in ? 256'h0 : _GEN_160; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_162 = 8'ha2 == io_in ? 256'h0 : _GEN_161; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_163 = 8'ha3 == io_in ? 256'h0 : _GEN_162; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_164 = 8'ha4 == io_in ? 256'h0 : _GEN_163; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_165 = 8'ha5 == io_in ? 256'h0 : _GEN_164; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_166 = 8'ha6 == io_in ? 256'h0 : _GEN_165; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_167 = 8'ha7 == io_in ? 256'h0 : _GEN_166; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_168 = 8'ha8 == io_in ? 256'h0 : _GEN_167; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_169 = 8'ha9 == io_in ? 256'h0 : _GEN_168; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_170 = 8'haa == io_in ? 256'h0 : _GEN_169; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_171 = 8'hab == io_in ? 256'h0 : _GEN_170; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_172 = 8'hac == io_in ? 256'h0 : _GEN_171; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_173 = 8'had == io_in ? 256'h0 : _GEN_172; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_174 = 8'hae == io_in ? 256'h0 : _GEN_173; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_175 = 8'haf == io_in ? 256'h0 : _GEN_174; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_176 = 8'hb0 == io_in ? 256'h0 : _GEN_175; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_177 = 8'hb1 == io_in ? 256'h0 : _GEN_176; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_178 = 8'hb2 == io_in ? 256'h0 : _GEN_177; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_179 = 8'hb3 == io_in ? 256'h0 : _GEN_178; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_180 = 8'hb4 == io_in ? 256'h0 : _GEN_179; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_181 = 8'hb5 == io_in ? 256'h0 : _GEN_180; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_182 = 8'hb6 == io_in ? 256'h0 : _GEN_181; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_183 = 8'hb7 == io_in ? 256'h0 : _GEN_182; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_184 = 8'hb8 == io_in ? 256'h0 : _GEN_183; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_185 = 8'hb9 == io_in ? 256'h0 : _GEN_184; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_186 = 8'hba == io_in ? 256'h0 : _GEN_185; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_187 = 8'hbb == io_in ? 256'h0 : _GEN_186; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_188 = 8'hbc == io_in ? 256'h0 : _GEN_187; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_189 = 8'hbd == io_in ? 256'h0 : _GEN_188; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_190 = 8'hbe == io_in ? 256'h0 : _GEN_189; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_191 = 8'hbf == io_in ? 256'h0 : _GEN_190; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_192 = 8'hc0 == io_in ? 256'h0 : _GEN_191; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_193 = 8'hc1 == io_in ? 256'h0 : _GEN_192; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_194 = 8'hc2 == io_in ? 256'h0 : _GEN_193; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_195 = 8'hc3 == io_in ? 256'h0 : _GEN_194; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_196 = 8'hc4 == io_in ? 256'h0 : _GEN_195; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_197 = 8'hc5 == io_in ? 256'h0 : _GEN_196; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_198 = 8'hc6 == io_in ? 256'h0 : _GEN_197; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_199 = 8'hc7 == io_in ? 256'h0 : _GEN_198; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_200 = 8'hc8 == io_in ? 256'h0 : _GEN_199; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_201 = 8'hc9 == io_in ? 256'h0 : _GEN_200; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_202 = 8'hca == io_in ? 256'h0 : _GEN_201; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_203 = 8'hcb == io_in ? 256'h0 : _GEN_202; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_204 = 8'hcc == io_in ? 256'h0 : _GEN_203; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_205 = 8'hcd == io_in ? 256'h0 : _GEN_204; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_206 = 8'hce == io_in ? 256'h0 : _GEN_205; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_207 = 8'hcf == io_in ? 256'h0 : _GEN_206; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_208 = 8'hd0 == io_in ? 256'h0 : _GEN_207; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_209 = 8'hd1 == io_in ? 256'h0 : _GEN_208; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_210 = 8'hd2 == io_in ? 256'h0 : _GEN_209; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_211 = 8'hd3 == io_in ? 256'h0 : _GEN_210; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_212 = 8'hd4 == io_in ? 256'h0 : _GEN_211; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_213 = 8'hd5 == io_in ? 256'h0 : _GEN_212; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_214 = 8'hd6 == io_in ? 256'h0 : _GEN_213; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_215 = 8'hd7 == io_in ? 256'h0 : _GEN_214; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_216 = 8'hd8 == io_in ? 256'h0 : _GEN_215; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_217 = 8'hd9 == io_in ? 256'h0 : _GEN_216; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_218 = 8'hda == io_in ? 256'h0 : _GEN_217; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_219 = 8'hdb == io_in ? 256'h0 : _GEN_218; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_220 = 8'hdc == io_in ? 256'h0 : _GEN_219; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_221 = 8'hdd == io_in ? 256'h0 : _GEN_220; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_222 = 8'hde == io_in ? 256'h0 : _GEN_221; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_223 = 8'hdf == io_in ? 256'h0 : _GEN_222; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_224 = 8'he0 == io_in ? 256'h0 : _GEN_223; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_225 = 8'he1 == io_in ? 256'h0 : _GEN_224; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_226 = 8'he2 == io_in ? 256'h0 : _GEN_225; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_227 = 8'he3 == io_in ? 256'h0 : _GEN_226; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_228 = 8'he4 == io_in ? 256'h0 : _GEN_227; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_229 = 8'he5 == io_in ? 256'h0 : _GEN_228; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_230 = 8'he6 == io_in ? 256'h0 : _GEN_229; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_231 = 8'he7 == io_in ? 256'h0 : _GEN_230; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_232 = 8'he8 == io_in ? 256'h0 : _GEN_231; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_233 = 8'he9 == io_in ? 256'h0 : _GEN_232; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_234 = 8'hea == io_in ? 256'h0 : _GEN_233; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_235 = 8'heb == io_in ? 256'h0 : _GEN_234; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_236 = 8'hec == io_in ? 256'h0 : _GEN_235; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_237 = 8'hed == io_in ? 256'h0 : _GEN_236; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_238 = 8'hee == io_in ? 256'h0 : _GEN_237; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_239 = 8'hef == io_in ? 256'h0 : _GEN_238; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_240 = 8'hf0 == io_in ? 256'h0 : _GEN_239; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_241 = 8'hf1 == io_in ? 256'h0 : _GEN_240; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_242 = 8'hf2 == io_in ? 256'h0 : _GEN_241; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_243 = 8'hf3 == io_in ? 256'h0 : _GEN_242; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_244 = 8'hf4 == io_in ? 256'h0 : _GEN_243; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_245 = 8'hf5 == io_in ? 256'h0 : _GEN_244; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_246 = 8'hf6 == io_in ? 256'h0 : _GEN_245; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_247 = 8'hf7 == io_in ? 256'h0 : _GEN_246; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_248 = 8'hf8 == io_in ? 256'h0 : _GEN_247; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_249 = 8'hf9 == io_in ? 256'h0 : _GEN_248; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_250 = 8'hfa == io_in ? 256'h0 : _GEN_249; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_251 = 8'hfb == io_in ? 256'h0 : _GEN_250; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_252 = 8'hfc == io_in ? 256'h0 : _GEN_251; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_253 = 8'hfd == io_in ? 256'h0 : _GEN_252; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_254 = 8'hfe == io_in ? 256'h0 : _GEN_253; // @[ps2.scala 242:11 ps2.scala 242:11]
  wire [255:0] _GEN_255 = 8'hff == io_in ? 256'h0 : _GEN_254; // @[ps2.scala 242:11 ps2.scala 242:11]
  assign io_out = _GEN_255[7:0]; // @[ps2.scala 242:11]
  always @(posedge clock) begin
    if (reset) begin // @[ps2.scala 201:22]
      table_21 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_21 <= 256'h71; // @[ps2.scala 220:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_22 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_22 <= 256'h31; // @[ps2.scala 232:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_26 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_26 <= 256'h7a; // @[ps2.scala 229:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_27 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_27 <= 256'h73; // @[ps2.scala 222:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_28 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_28 <= 256'h61; // @[ps2.scala 204:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_29 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_29 <= 256'h77; // @[ps2.scala 226:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_30 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_30 <= 256'h32; // @[ps2.scala 233:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_33 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_33 <= 256'h63; // @[ps2.scala 206:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_34 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_34 <= 256'h78; // @[ps2.scala 227:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_35 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_35 <= 256'h64; // @[ps2.scala 207:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_36 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_36 <= 256'h65; // @[ps2.scala 208:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_37 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_37 <= 256'h34; // @[ps2.scala 235:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_38 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_38 <= 256'h33; // @[ps2.scala 234:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_42 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_42 <= 256'h76; // @[ps2.scala 225:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_43 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_43 <= 256'h66; // @[ps2.scala 209:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_44 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_44 <= 256'h74; // @[ps2.scala 223:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_45 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_45 <= 256'h72; // @[ps2.scala 221:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_46 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_46 <= 256'h35; // @[ps2.scala 236:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_49 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_49 <= 256'h6e; // @[ps2.scala 217:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_50 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_50 <= 256'h62; // @[ps2.scala 205:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_51 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_51 <= 256'h68; // @[ps2.scala 211:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_52 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_52 <= 256'h67; // @[ps2.scala 210:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_53 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_53 <= 256'h79; // @[ps2.scala 228:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_54 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_54 <= 256'h36; // @[ps2.scala 237:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_58 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_58 <= 256'h6d; // @[ps2.scala 216:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_59 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_59 <= 256'h6a; // @[ps2.scala 213:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_60 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_60 <= 256'h75; // @[ps2.scala 224:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_61 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_61 <= 256'h37; // @[ps2.scala 238:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_62 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_62 <= 256'h38; // @[ps2.scala 239:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_66 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_66 <= 256'h6b; // @[ps2.scala 214:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_67 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_67 <= 256'h69; // @[ps2.scala 212:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_68 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_68 <= 256'h6f; // @[ps2.scala 218:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_69 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_69 <= 256'h30; // @[ps2.scala 231:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_70 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_70 <= 256'h39; // @[ps2.scala 240:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_75 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_75 <= 256'h6c; // @[ps2.scala 215:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_77 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_77 <= 256'h70; // @[ps2.scala 219:19]
    end
    if (reset) begin // @[ps2.scala 201:22]
      table_90 <= 256'h0; // @[ps2.scala 201:22]
    end else begin
      table_90 <= 256'ha; // @[ps2.scala 202:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  table_21 = _RAND_0[255:0];
  _RAND_1 = {8{`RANDOM}};
  table_22 = _RAND_1[255:0];
  _RAND_2 = {8{`RANDOM}};
  table_26 = _RAND_2[255:0];
  _RAND_3 = {8{`RANDOM}};
  table_27 = _RAND_3[255:0];
  _RAND_4 = {8{`RANDOM}};
  table_28 = _RAND_4[255:0];
  _RAND_5 = {8{`RANDOM}};
  table_29 = _RAND_5[255:0];
  _RAND_6 = {8{`RANDOM}};
  table_30 = _RAND_6[255:0];
  _RAND_7 = {8{`RANDOM}};
  table_33 = _RAND_7[255:0];
  _RAND_8 = {8{`RANDOM}};
  table_34 = _RAND_8[255:0];
  _RAND_9 = {8{`RANDOM}};
  table_35 = _RAND_9[255:0];
  _RAND_10 = {8{`RANDOM}};
  table_36 = _RAND_10[255:0];
  _RAND_11 = {8{`RANDOM}};
  table_37 = _RAND_11[255:0];
  _RAND_12 = {8{`RANDOM}};
  table_38 = _RAND_12[255:0];
  _RAND_13 = {8{`RANDOM}};
  table_42 = _RAND_13[255:0];
  _RAND_14 = {8{`RANDOM}};
  table_43 = _RAND_14[255:0];
  _RAND_15 = {8{`RANDOM}};
  table_44 = _RAND_15[255:0];
  _RAND_16 = {8{`RANDOM}};
  table_45 = _RAND_16[255:0];
  _RAND_17 = {8{`RANDOM}};
  table_46 = _RAND_17[255:0];
  _RAND_18 = {8{`RANDOM}};
  table_49 = _RAND_18[255:0];
  _RAND_19 = {8{`RANDOM}};
  table_50 = _RAND_19[255:0];
  _RAND_20 = {8{`RANDOM}};
  table_51 = _RAND_20[255:0];
  _RAND_21 = {8{`RANDOM}};
  table_52 = _RAND_21[255:0];
  _RAND_22 = {8{`RANDOM}};
  table_53 = _RAND_22[255:0];
  _RAND_23 = {8{`RANDOM}};
  table_54 = _RAND_23[255:0];
  _RAND_24 = {8{`RANDOM}};
  table_58 = _RAND_24[255:0];
  _RAND_25 = {8{`RANDOM}};
  table_59 = _RAND_25[255:0];
  _RAND_26 = {8{`RANDOM}};
  table_60 = _RAND_26[255:0];
  _RAND_27 = {8{`RANDOM}};
  table_61 = _RAND_27[255:0];
  _RAND_28 = {8{`RANDOM}};
  table_62 = _RAND_28[255:0];
  _RAND_29 = {8{`RANDOM}};
  table_66 = _RAND_29[255:0];
  _RAND_30 = {8{`RANDOM}};
  table_67 = _RAND_30[255:0];
  _RAND_31 = {8{`RANDOM}};
  table_68 = _RAND_31[255:0];
  _RAND_32 = {8{`RANDOM}};
  table_69 = _RAND_32[255:0];
  _RAND_33 = {8{`RANDOM}};
  table_70 = _RAND_33[255:0];
  _RAND_34 = {8{`RANDOM}};
  table_75 = _RAND_34[255:0];
  _RAND_35 = {8{`RANDOM}};
  table_77 = _RAND_35[255:0];
  _RAND_36 = {8{`RANDOM}};
  table_90 = _RAND_36[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module seg(
  input  [3:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_0 = io_in == 4'hf ? 8'h8e : 8'hff; // @[ps2.scala 286:33 ps2.scala 287:19 ps2.scala 254:11]
  wire [7:0] _GEN_1 = io_in == 4'he ? 8'h86 : _GEN_0; // @[ps2.scala 284:33 ps2.scala 285:19]
  wire [7:0] _GEN_2 = io_in == 4'hd ? 8'ha1 : _GEN_1; // @[ps2.scala 282:33 ps2.scala 283:19]
  wire [7:0] _GEN_3 = io_in == 4'hc ? 8'hc6 : _GEN_2; // @[ps2.scala 280:33 ps2.scala 281:19]
  wire [7:0] _GEN_4 = io_in == 4'hb ? 8'h83 : _GEN_3; // @[ps2.scala 278:33 ps2.scala 279:19]
  wire [7:0] _GEN_5 = io_in == 4'ha ? 8'h88 : _GEN_4; // @[ps2.scala 276:33 ps2.scala 277:19]
  wire [7:0] _GEN_6 = io_in == 4'h9 ? 8'h90 : _GEN_5; // @[ps2.scala 274:32 ps2.scala 275:19]
  wire [7:0] _GEN_7 = io_in == 4'h8 ? 8'h80 : _GEN_6; // @[ps2.scala 272:32 ps2.scala 273:19]
  wire [7:0] _GEN_8 = io_in == 4'h7 ? 8'hf8 : _GEN_7; // @[ps2.scala 270:32 ps2.scala 271:19]
  wire [7:0] _GEN_9 = io_in == 4'h6 ? 8'h82 : _GEN_8; // @[ps2.scala 268:32 ps2.scala 269:19]
  wire [7:0] _GEN_10 = io_in == 4'h5 ? 8'h92 : _GEN_9; // @[ps2.scala 266:32 ps2.scala 267:19]
  wire [7:0] _GEN_11 = io_in == 4'h4 ? 8'h99 : _GEN_10; // @[ps2.scala 264:32 ps2.scala 265:19]
  wire [7:0] _GEN_12 = io_in == 4'h3 ? 8'hb0 : _GEN_11; // @[ps2.scala 262:32 ps2.scala 263:19]
  wire [7:0] _GEN_13 = io_in == 4'h2 ? 8'ha4 : _GEN_12; // @[ps2.scala 260:32 ps2.scala 261:19]
  wire [7:0] _GEN_14 = io_in == 4'h1 ? 8'hf9 : _GEN_13; // @[ps2.scala 258:32 ps2.scala 259:19]
  assign io_out = io_in == 4'h0 ? 8'hc0 : _GEN_14; // @[ps2.scala 256:26 ps2.scala 257:19]
endmodule
module ps2(
  input        clock,
  input        reset,
  input        io_ps2_clk,
  input        io_ps2_data,
  output [7:0] io_ascii,
  output       io_ready,
  output [7:0] io_bcd8seg_0,
  output [7:0] io_bcd8seg_1,
  output [7:0] io_bcd8seg_2,
  output [7:0] io_bcd8seg_3,
  output [7:0] io_bcd8seg_4,
  output [7:0] io_bcd8seg_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ps2_clock; // @[ps2.scala 16:19]
  wire  ps2_io_ps2_clk; // @[ps2.scala 16:19]
  wire  ps2_io_ps2_data; // @[ps2.scala 16:19]
  wire  ps2_io_nextdata_n; // @[ps2.scala 16:19]
  wire [7:0] ps2_io_data; // @[ps2.scala 16:19]
  wire  ps2_io_ready; // @[ps2.scala 16:19]
  wire  mm_clock; // @[ps2.scala 93:18]
  wire  mm_reset; // @[ps2.scala 93:18]
  wire [7:0] mm_io_in; // @[ps2.scala 93:18]
  wire [7:0] mm_io_out; // @[ps2.scala 93:18]
  wire [3:0] m0_io_in; // @[ps2.scala 98:18]
  wire [7:0] m0_io_out; // @[ps2.scala 98:18]
  wire [3:0] m1_io_in; // @[ps2.scala 102:18]
  wire [7:0] m1_io_out; // @[ps2.scala 102:18]
  wire [3:0] m2_io_in; // @[ps2.scala 106:18]
  wire [7:0] m2_io_out; // @[ps2.scala 106:18]
  wire [3:0] m3_io_in; // @[ps2.scala 110:18]
  wire [7:0] m3_io_out; // @[ps2.scala 110:18]
  wire [3:0] m4_io_in; // @[ps2.scala 114:18]
  wire [7:0] m4_io_out; // @[ps2.scala 114:18]
  wire [3:0] m5_io_in; // @[ps2.scala 118:18]
  wire [7:0] m5_io_out; // @[ps2.scala 118:18]
  reg [7:0] data; // @[ps2.scala 12:21]
  reg  ready; // @[ps2.scala 13:18]
  reg  nextdata; // @[ps2.scala 15:21]
  reg [3:0] now; // @[ps2.scala 30:20]
  reg [3:0] next; // @[ps2.scala 31:21]
  wire  _T = now == 4'h1; // @[ps2.scala 33:13]
  wire [1:0] _GEN_0 = ready ? 2'h2 : 2'h1; // @[ps2.scala 34:26 ps2.scala 35:17 ps2.scala 37:17]
  wire  _T_2 = now == 4'h2; // @[ps2.scala 39:19]
  wire  _T_3 = now == 4'h4; // @[ps2.scala 41:19]
  wire  _T_4 = now == 4'h8; // @[ps2.scala 43:19]
  reg [23:0] ps2segdata; // @[ps2.scala 48:27]
  wire [15:0] ps2segdata_hi = ps2segdata[15:0]; // @[ps2.scala 54:35]
  wire [23:0] _ps2segdata_T = {ps2segdata_hi,data}; // @[Cat.scala 30:58]
  wire  _GEN_6 = _T_2 ? nextdata : 1'h1; // @[ps2.scala 53:25 ps2.scala 15:21 ps2.scala 56:17]
  wire  _GEN_7 = _T_3 | _T_4 ? 1'h0 : _GEN_6; // @[ps2.scala 51:35 ps2.scala 52:17]
  reg [99:0] num; // @[ps2.scala 61:16]
  reg  segen; // @[ps2.scala 64:22]
  reg [1:0] ss; // @[ps2.scala 65:19]
  wire [99:0] _num_T_1 = num + 100'h1; // @[ps2.scala 67:17]
  wire  _T_13 = ps2segdata[23:16] == 8'hf0; // @[ps2.scala 69:36]
  wire  _T_18 = ss == 2'h2; // @[ps2.scala 74:20]
  wire [99:0] _GEN_1 = num % 100'hc350; // @[ps2.scala 78:21]
  wire [15:0] _T_19 = _GEN_1[15:0]; // @[ps2.scala 78:21]
  wire  _T_20 = _T_19 == 16'h0; // @[ps2.scala 78:29]
  wire  _GEN_15 = _T_13 ? 1'h0 : _T_20; // @[ps2.scala 81:46 ps2.scala 83:25]
  wire  _GEN_17 = num < 100'h2710 ? _T_18 : _GEN_15; // @[ps2.scala 68:26]
  wire  ss_hi = ss[0]; // @[ps2.scala 88:15]
  wire [1:0] _ss_T = {ss_hi,segen}; // @[Cat.scala 30:58]
  reg [7:0] ascii; // @[ps2.scala 92:22]
  ps2_keyboard ps2 ( // @[ps2.scala 16:19]
    .clock(ps2_clock),
    .io_ps2_clk(ps2_io_ps2_clk),
    .io_ps2_data(ps2_io_ps2_data),
    .io_nextdata_n(ps2_io_nextdata_n),
    .io_data(ps2_io_data),
    .io_ready(ps2_io_ready)
  );
  ps2ascii mm ( // @[ps2.scala 93:18]
    .clock(mm_clock),
    .reset(mm_reset),
    .io_in(mm_io_in),
    .io_out(mm_io_out)
  );
  seg m0 ( // @[ps2.scala 98:18]
    .io_in(m0_io_in),
    .io_out(m0_io_out)
  );
  seg m1 ( // @[ps2.scala 102:18]
    .io_in(m1_io_in),
    .io_out(m1_io_out)
  );
  seg m2 ( // @[ps2.scala 106:18]
    .io_in(m2_io_in),
    .io_out(m2_io_out)
  );
  seg m3 ( // @[ps2.scala 110:18]
    .io_in(m3_io_in),
    .io_out(m3_io_out)
  );
  seg m4 ( // @[ps2.scala 114:18]
    .io_in(m4_io_in),
    .io_out(m4_io_out)
  );
  seg m5 ( // @[ps2.scala 118:18]
    .io_in(m5_io_in),
    .io_out(m5_io_out)
  );
  assign io_ascii = ascii; // @[ps2.scala 96:13]
  assign io_ready = data != 8'h0 & _GEN_17; // @[ps2.scala 66:21 ps2.scala 59:13]
  assign io_bcd8seg_0 = m0_io_out; // @[ps2.scala 101:18]
  assign io_bcd8seg_1 = m1_io_out; // @[ps2.scala 105:18]
  assign io_bcd8seg_2 = m2_io_out; // @[ps2.scala 109:18]
  assign io_bcd8seg_3 = m3_io_out; // @[ps2.scala 113:18]
  assign io_bcd8seg_4 = m4_io_out; // @[ps2.scala 117:18]
  assign io_bcd8seg_5 = m5_io_out; // @[ps2.scala 121:18]
  assign ps2_clock = clock;
  assign ps2_io_ps2_clk = io_ps2_clk; // @[ps2.scala 18:19]
  assign ps2_io_ps2_data = io_ps2_data; // @[ps2.scala 19:20]
  assign ps2_io_nextdata_n = nextdata; // @[ps2.scala 20:22]
  assign mm_clock = clock;
  assign mm_reset = reset;
  assign mm_io_in = ps2segdata[7:0]; // @[ps2.scala 94:25]
  assign m0_io_in = ps2segdata[3:0]; // @[ps2.scala 100:25]
  assign m1_io_in = ps2segdata[7:4]; // @[ps2.scala 104:25]
  assign m2_io_in = ps2segdata[11:8]; // @[ps2.scala 108:25]
  assign m3_io_in = ps2segdata[15:12]; // @[ps2.scala 112:25]
  assign m4_io_in = ps2segdata[19:16]; // @[ps2.scala 116:25]
  assign m5_io_in = ps2segdata[23:20]; // @[ps2.scala 120:25]
  always @(posedge clock) begin
    if (reset) begin // @[ps2.scala 12:21]
      data <= 8'h0; // @[ps2.scala 12:21]
    end else begin
      data <= ps2_io_data; // @[ps2.scala 21:9]
    end
    ready <= ps2_io_ready; // @[ps2.scala 22:10]
    nextdata <= _T | _GEN_7; // @[ps2.scala 49:19 ps2.scala 50:17]
    if (reset) begin // @[ps2.scala 30:20]
      now <= 4'h1; // @[ps2.scala 30:20]
    end else begin
      now <= next; // @[ps2.scala 32:8]
    end
    if (reset) begin // @[ps2.scala 31:21]
      next <= 4'h1; // @[ps2.scala 31:21]
    end else if (now == 4'h1) begin // @[ps2.scala 33:19]
      next <= {{2'd0}, _GEN_0};
    end else if (now == 4'h2) begin // @[ps2.scala 39:25]
      next <= 4'h4; // @[ps2.scala 40:13]
    end else if (now == 4'h4) begin // @[ps2.scala 41:25]
      next <= 4'h8; // @[ps2.scala 42:13]
    end else begin
      next <= 4'h1;
    end
    if (reset) begin // @[ps2.scala 48:27]
      ps2segdata <= 24'h0; // @[ps2.scala 48:27]
    end else if (!(_T)) begin // @[ps2.scala 49:19]
      if (!(_T_3 | _T_4)) begin // @[ps2.scala 51:35]
        if (_T_2) begin // @[ps2.scala 53:25]
          ps2segdata <= _ps2segdata_T; // @[ps2.scala 54:19]
        end
      end
    end
    if (data != 8'h0) begin // @[ps2.scala 66:21]
      if (num < 100'h2710) begin // @[ps2.scala 68:26]
        num <= _num_T_1; // @[ps2.scala 67:12]
      end else if (_T_13) begin // @[ps2.scala 81:46]
        num <= 100'h0; // @[ps2.scala 82:20]
      end else begin
        num <= _num_T_1; // @[ps2.scala 67:12]
      end
    end else begin
      num <= 100'h0; // @[ps2.scala 63:8]
    end
    if (reset) begin // @[ps2.scala 64:22]
      segen <= 1'h0; // @[ps2.scala 64:22]
    end else if (data != 8'h0) begin // @[ps2.scala 66:21]
      if (num < 100'h2710) begin // @[ps2.scala 68:26]
        if (ps2segdata[23:16] == 8'hf0 & ps2segdata[15:8] == ps2segdata[7:0]) begin // @[ps2.scala 69:86]
          segen <= 1'h0; // @[ps2.scala 70:22]
        end else begin
          segen <= 1'h1; // @[ps2.scala 72:22]
        end
      end
    end
    if (reset) begin // @[ps2.scala 65:19]
      ss <= 2'h0; // @[ps2.scala 65:19]
    end else begin
      ss <= _ss_T; // @[ps2.scala 88:7]
    end
    if (reset) begin // @[ps2.scala 92:22]
      ascii <= 8'h0; // @[ps2.scala 92:22]
    end else begin
      ascii <= mm_io_out; // @[ps2.scala 95:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  ready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  nextdata = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  now = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  next = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  ps2segdata = _RAND_5[23:0];
  _RAND_6 = {4{`RANDOM}};
  num = _RAND_6[99:0];
  _RAND_7 = {1{`RANDOM}};
  segen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ss = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ascii = _RAND_9[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vmem(
  input         clock,
  input         reset,
  input  [9:0]  io_h_addr,
  input  [8:0]  io_v_addr,
  input  [7:0]  io_ascii,
  input         io_w_en,
  output [23:0] io_vga_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
`endif // RANDOMIZE_REG_INIT
  reg [11:0] vga_mem [0:4095]; // @[vga.scala 16:30]
  wire [11:0] vga_mem_MPORT_data; // @[vga.scala 16:30]
  wire [11:0] vga_mem_MPORT_addr; // @[vga.scala 16:30]
  reg [11:0] vga_mem_MPORT_addr_pipe_0;
  reg [23:0] rdwrPort; // @[vga.scala 13:27]
  reg [7:0] ram_0; // @[vga.scala 14:20]
  reg [7:0] ram_1; // @[vga.scala 14:20]
  reg [7:0] ram_2; // @[vga.scala 14:20]
  reg [7:0] ram_3; // @[vga.scala 14:20]
  reg [7:0] ram_4; // @[vga.scala 14:20]
  reg [7:0] ram_5; // @[vga.scala 14:20]
  reg [7:0] ram_6; // @[vga.scala 14:20]
  reg [7:0] ram_7; // @[vga.scala 14:20]
  reg [7:0] ram_8; // @[vga.scala 14:20]
  reg [7:0] ram_9; // @[vga.scala 14:20]
  reg [7:0] ram_10; // @[vga.scala 14:20]
  reg [7:0] ram_11; // @[vga.scala 14:20]
  reg [7:0] ram_12; // @[vga.scala 14:20]
  reg [7:0] ram_13; // @[vga.scala 14:20]
  reg [7:0] ram_14; // @[vga.scala 14:20]
  reg [7:0] ram_15; // @[vga.scala 14:20]
  reg [7:0] ram_16; // @[vga.scala 14:20]
  reg [7:0] ram_17; // @[vga.scala 14:20]
  reg [7:0] ram_18; // @[vga.scala 14:20]
  reg [7:0] ram_19; // @[vga.scala 14:20]
  reg [7:0] ram_20; // @[vga.scala 14:20]
  reg [7:0] ram_21; // @[vga.scala 14:20]
  reg [7:0] ram_22; // @[vga.scala 14:20]
  reg [7:0] ram_23; // @[vga.scala 14:20]
  reg [7:0] ram_24; // @[vga.scala 14:20]
  reg [7:0] ram_25; // @[vga.scala 14:20]
  reg [7:0] ram_26; // @[vga.scala 14:20]
  reg [7:0] ram_27; // @[vga.scala 14:20]
  reg [7:0] ram_28; // @[vga.scala 14:20]
  reg [7:0] ram_29; // @[vga.scala 14:20]
  reg [7:0] ram_30; // @[vga.scala 14:20]
  reg [7:0] ram_31; // @[vga.scala 14:20]
  reg [7:0] ram_32; // @[vga.scala 14:20]
  reg [7:0] ram_33; // @[vga.scala 14:20]
  reg [7:0] ram_34; // @[vga.scala 14:20]
  reg [7:0] ram_35; // @[vga.scala 14:20]
  reg [7:0] ram_36; // @[vga.scala 14:20]
  reg [7:0] ram_37; // @[vga.scala 14:20]
  reg [7:0] ram_38; // @[vga.scala 14:20]
  reg [7:0] ram_39; // @[vga.scala 14:20]
  reg [7:0] ram_40; // @[vga.scala 14:20]
  reg [7:0] ram_41; // @[vga.scala 14:20]
  reg [7:0] ram_42; // @[vga.scala 14:20]
  reg [7:0] ram_43; // @[vga.scala 14:20]
  reg [7:0] ram_44; // @[vga.scala 14:20]
  reg [7:0] ram_45; // @[vga.scala 14:20]
  reg [7:0] ram_46; // @[vga.scala 14:20]
  reg [7:0] ram_47; // @[vga.scala 14:20]
  reg [7:0] ram_48; // @[vga.scala 14:20]
  reg [7:0] ram_49; // @[vga.scala 14:20]
  reg [7:0] ram_50; // @[vga.scala 14:20]
  reg [7:0] ram_51; // @[vga.scala 14:20]
  reg [7:0] ram_52; // @[vga.scala 14:20]
  reg [7:0] ram_53; // @[vga.scala 14:20]
  reg [7:0] ram_54; // @[vga.scala 14:20]
  reg [7:0] ram_55; // @[vga.scala 14:20]
  reg [7:0] ram_56; // @[vga.scala 14:20]
  reg [7:0] ram_57; // @[vga.scala 14:20]
  reg [7:0] ram_58; // @[vga.scala 14:20]
  reg [7:0] ram_59; // @[vga.scala 14:20]
  reg [7:0] ram_60; // @[vga.scala 14:20]
  reg [7:0] ram_61; // @[vga.scala 14:20]
  reg [7:0] ram_62; // @[vga.scala 14:20]
  reg [7:0] ram_63; // @[vga.scala 14:20]
  reg [7:0] ram_64; // @[vga.scala 14:20]
  reg [7:0] ram_65; // @[vga.scala 14:20]
  reg [7:0] ram_66; // @[vga.scala 14:20]
  reg [7:0] ram_67; // @[vga.scala 14:20]
  reg [7:0] ram_68; // @[vga.scala 14:20]
  reg [7:0] ram_69; // @[vga.scala 14:20]
  reg [7:0] ram_70; // @[vga.scala 14:20]
  reg [7:0] ram_71; // @[vga.scala 14:20]
  reg [7:0] ram_72; // @[vga.scala 14:20]
  reg [7:0] ram_73; // @[vga.scala 14:20]
  reg [7:0] ram_74; // @[vga.scala 14:20]
  reg [7:0] ram_75; // @[vga.scala 14:20]
  reg [7:0] ram_76; // @[vga.scala 14:20]
  reg [7:0] ram_77; // @[vga.scala 14:20]
  reg [7:0] ram_78; // @[vga.scala 14:20]
  reg [7:0] ram_79; // @[vga.scala 14:20]
  reg [7:0] ram_80; // @[vga.scala 14:20]
  reg [7:0] ram_81; // @[vga.scala 14:20]
  reg [7:0] ram_82; // @[vga.scala 14:20]
  reg [7:0] ram_83; // @[vga.scala 14:20]
  reg [7:0] ram_84; // @[vga.scala 14:20]
  reg [7:0] ram_85; // @[vga.scala 14:20]
  reg [7:0] ram_86; // @[vga.scala 14:20]
  reg [7:0] ram_87; // @[vga.scala 14:20]
  reg [7:0] ram_88; // @[vga.scala 14:20]
  reg [7:0] ram_89; // @[vga.scala 14:20]
  reg [7:0] ram_90; // @[vga.scala 14:20]
  reg [7:0] ram_91; // @[vga.scala 14:20]
  reg [7:0] ram_92; // @[vga.scala 14:20]
  reg [7:0] ram_93; // @[vga.scala 14:20]
  reg [7:0] ram_94; // @[vga.scala 14:20]
  reg [7:0] ram_95; // @[vga.scala 14:20]
  reg [7:0] ram_96; // @[vga.scala 14:20]
  reg [7:0] ram_97; // @[vga.scala 14:20]
  reg [7:0] ram_98; // @[vga.scala 14:20]
  reg [7:0] ram_99; // @[vga.scala 14:20]
  reg [7:0] ram_100; // @[vga.scala 14:20]
  reg [7:0] ram_101; // @[vga.scala 14:20]
  reg [7:0] ram_102; // @[vga.scala 14:20]
  reg [7:0] ram_103; // @[vga.scala 14:20]
  reg [7:0] ram_104; // @[vga.scala 14:20]
  reg [7:0] ram_105; // @[vga.scala 14:20]
  reg [7:0] ram_106; // @[vga.scala 14:20]
  reg [7:0] ram_107; // @[vga.scala 14:20]
  reg [7:0] ram_108; // @[vga.scala 14:20]
  reg [7:0] ram_109; // @[vga.scala 14:20]
  reg [7:0] ram_110; // @[vga.scala 14:20]
  reg [7:0] ram_111; // @[vga.scala 14:20]
  reg [7:0] ram_112; // @[vga.scala 14:20]
  reg [7:0] ram_113; // @[vga.scala 14:20]
  reg [7:0] ram_114; // @[vga.scala 14:20]
  reg [7:0] ram_115; // @[vga.scala 14:20]
  reg [7:0] ram_116; // @[vga.scala 14:20]
  reg [7:0] ram_117; // @[vga.scala 14:20]
  reg [7:0] ram_118; // @[vga.scala 14:20]
  reg [7:0] ram_119; // @[vga.scala 14:20]
  reg [7:0] ram_120; // @[vga.scala 14:20]
  reg [7:0] ram_121; // @[vga.scala 14:20]
  reg [7:0] ram_122; // @[vga.scala 14:20]
  reg [7:0] ram_123; // @[vga.scala 14:20]
  reg [7:0] ram_124; // @[vga.scala 14:20]
  reg [7:0] ram_125; // @[vga.scala 14:20]
  reg [7:0] ram_126; // @[vga.scala 14:20]
  reg [7:0] ram_127; // @[vga.scala 14:20]
  reg [7:0] ram_128; // @[vga.scala 14:20]
  reg [7:0] ram_129; // @[vga.scala 14:20]
  reg [7:0] ram_130; // @[vga.scala 14:20]
  reg [7:0] ram_131; // @[vga.scala 14:20]
  reg [7:0] ram_132; // @[vga.scala 14:20]
  reg [7:0] ram_133; // @[vga.scala 14:20]
  reg [7:0] ram_134; // @[vga.scala 14:20]
  reg [7:0] ram_135; // @[vga.scala 14:20]
  reg [7:0] ram_136; // @[vga.scala 14:20]
  reg [7:0] ram_137; // @[vga.scala 14:20]
  reg [7:0] ram_138; // @[vga.scala 14:20]
  reg [7:0] ram_139; // @[vga.scala 14:20]
  reg [7:0] ram_140; // @[vga.scala 14:20]
  reg [7:0] ram_141; // @[vga.scala 14:20]
  reg [7:0] ram_142; // @[vga.scala 14:20]
  reg [7:0] ram_143; // @[vga.scala 14:20]
  reg [7:0] ram_144; // @[vga.scala 14:20]
  reg [7:0] ram_145; // @[vga.scala 14:20]
  reg [7:0] ram_146; // @[vga.scala 14:20]
  reg [7:0] ram_147; // @[vga.scala 14:20]
  reg [7:0] ram_148; // @[vga.scala 14:20]
  reg [7:0] ram_149; // @[vga.scala 14:20]
  reg [7:0] ram_150; // @[vga.scala 14:20]
  reg [7:0] ram_151; // @[vga.scala 14:20]
  reg [7:0] ram_152; // @[vga.scala 14:20]
  reg [7:0] ram_153; // @[vga.scala 14:20]
  reg [7:0] ram_154; // @[vga.scala 14:20]
  reg [7:0] ram_155; // @[vga.scala 14:20]
  reg [7:0] ram_156; // @[vga.scala 14:20]
  reg [7:0] ram_157; // @[vga.scala 14:20]
  reg [7:0] ram_158; // @[vga.scala 14:20]
  reg [7:0] ram_159; // @[vga.scala 14:20]
  reg [7:0] ram_160; // @[vga.scala 14:20]
  reg [7:0] ram_161; // @[vga.scala 14:20]
  reg [7:0] ram_162; // @[vga.scala 14:20]
  reg [7:0] ram_163; // @[vga.scala 14:20]
  reg [7:0] ram_164; // @[vga.scala 14:20]
  reg [7:0] ram_165; // @[vga.scala 14:20]
  reg [7:0] ram_166; // @[vga.scala 14:20]
  reg [7:0] ram_167; // @[vga.scala 14:20]
  reg [7:0] ram_168; // @[vga.scala 14:20]
  reg [7:0] ram_169; // @[vga.scala 14:20]
  reg [7:0] ram_170; // @[vga.scala 14:20]
  reg [7:0] ram_171; // @[vga.scala 14:20]
  reg [7:0] ram_172; // @[vga.scala 14:20]
  reg [7:0] ram_173; // @[vga.scala 14:20]
  reg [7:0] ram_174; // @[vga.scala 14:20]
  reg [7:0] ram_175; // @[vga.scala 14:20]
  reg [7:0] ram_176; // @[vga.scala 14:20]
  reg [7:0] ram_177; // @[vga.scala 14:20]
  reg [7:0] ram_178; // @[vga.scala 14:20]
  reg [7:0] ram_179; // @[vga.scala 14:20]
  reg [7:0] ram_180; // @[vga.scala 14:20]
  reg [7:0] ram_181; // @[vga.scala 14:20]
  reg [7:0] ram_182; // @[vga.scala 14:20]
  reg [7:0] ram_183; // @[vga.scala 14:20]
  reg [7:0] ram_184; // @[vga.scala 14:20]
  reg [7:0] ram_185; // @[vga.scala 14:20]
  reg [7:0] ram_186; // @[vga.scala 14:20]
  reg [7:0] ram_187; // @[vga.scala 14:20]
  reg [7:0] ram_188; // @[vga.scala 14:20]
  reg [7:0] ram_189; // @[vga.scala 14:20]
  reg [7:0] ram_190; // @[vga.scala 14:20]
  reg [7:0] ram_191; // @[vga.scala 14:20]
  reg [7:0] ram_192; // @[vga.scala 14:20]
  reg [7:0] ram_193; // @[vga.scala 14:20]
  reg [7:0] ram_194; // @[vga.scala 14:20]
  reg [7:0] ram_195; // @[vga.scala 14:20]
  reg [7:0] ram_196; // @[vga.scala 14:20]
  reg [7:0] ram_197; // @[vga.scala 14:20]
  reg [7:0] ram_198; // @[vga.scala 14:20]
  reg [7:0] ram_199; // @[vga.scala 14:20]
  reg [7:0] ram_200; // @[vga.scala 14:20]
  reg [7:0] ram_201; // @[vga.scala 14:20]
  reg [7:0] ram_202; // @[vga.scala 14:20]
  reg [7:0] ram_203; // @[vga.scala 14:20]
  reg [7:0] ram_204; // @[vga.scala 14:20]
  reg [7:0] ram_205; // @[vga.scala 14:20]
  reg [7:0] ram_206; // @[vga.scala 14:20]
  reg [7:0] ram_207; // @[vga.scala 14:20]
  reg [7:0] ram_208; // @[vga.scala 14:20]
  reg [7:0] ram_209; // @[vga.scala 14:20]
  reg [7:0] ram_210; // @[vga.scala 14:20]
  reg [7:0] ram_211; // @[vga.scala 14:20]
  reg [7:0] ram_212; // @[vga.scala 14:20]
  reg [7:0] ram_213; // @[vga.scala 14:20]
  reg [7:0] ram_214; // @[vga.scala 14:20]
  reg [7:0] ram_215; // @[vga.scala 14:20]
  reg [7:0] ram_216; // @[vga.scala 14:20]
  reg [7:0] ram_217; // @[vga.scala 14:20]
  reg [7:0] ram_218; // @[vga.scala 14:20]
  reg [7:0] ram_219; // @[vga.scala 14:20]
  reg [7:0] ram_220; // @[vga.scala 14:20]
  reg [7:0] ram_221; // @[vga.scala 14:20]
  reg [7:0] ram_222; // @[vga.scala 14:20]
  reg [7:0] ram_223; // @[vga.scala 14:20]
  reg [7:0] ram_224; // @[vga.scala 14:20]
  reg [7:0] ram_225; // @[vga.scala 14:20]
  reg [7:0] ram_226; // @[vga.scala 14:20]
  reg [7:0] ram_227; // @[vga.scala 14:20]
  reg [7:0] ram_228; // @[vga.scala 14:20]
  reg [7:0] ram_229; // @[vga.scala 14:20]
  reg [7:0] ram_230; // @[vga.scala 14:20]
  reg [7:0] ram_231; // @[vga.scala 14:20]
  reg [7:0] ram_232; // @[vga.scala 14:20]
  reg [7:0] ram_233; // @[vga.scala 14:20]
  reg [7:0] ram_234; // @[vga.scala 14:20]
  reg [7:0] ram_235; // @[vga.scala 14:20]
  reg [7:0] ram_236; // @[vga.scala 14:20]
  reg [7:0] ram_237; // @[vga.scala 14:20]
  reg [7:0] ram_238; // @[vga.scala 14:20]
  reg [7:0] ram_239; // @[vga.scala 14:20]
  reg [7:0] ram_240; // @[vga.scala 14:20]
  reg [7:0] ram_241; // @[vga.scala 14:20]
  reg [7:0] ram_242; // @[vga.scala 14:20]
  reg [7:0] ram_243; // @[vga.scala 14:20]
  reg [7:0] ram_244; // @[vga.scala 14:20]
  reg [7:0] ram_245; // @[vga.scala 14:20]
  reg [7:0] ram_246; // @[vga.scala 14:20]
  reg [7:0] ram_247; // @[vga.scala 14:20]
  reg [7:0] ram_248; // @[vga.scala 14:20]
  reg [7:0] ram_249; // @[vga.scala 14:20]
  reg [7:0] ram_250; // @[vga.scala 14:20]
  reg [7:0] ram_251; // @[vga.scala 14:20]
  reg [7:0] ram_252; // @[vga.scala 14:20]
  reg [7:0] ram_253; // @[vga.scala 14:20]
  reg [7:0] ram_254; // @[vga.scala 14:20]
  reg [7:0] ram_255; // @[vga.scala 14:20]
  reg [7:0] ram_256; // @[vga.scala 14:20]
  reg [7:0] ram_257; // @[vga.scala 14:20]
  reg [7:0] ram_258; // @[vga.scala 14:20]
  reg [7:0] ram_259; // @[vga.scala 14:20]
  reg [7:0] ram_260; // @[vga.scala 14:20]
  reg [7:0] ram_261; // @[vga.scala 14:20]
  reg [7:0] ram_262; // @[vga.scala 14:20]
  reg [7:0] ram_263; // @[vga.scala 14:20]
  reg [7:0] ram_264; // @[vga.scala 14:20]
  reg [7:0] ram_265; // @[vga.scala 14:20]
  reg [7:0] ram_266; // @[vga.scala 14:20]
  reg [7:0] ram_267; // @[vga.scala 14:20]
  reg [7:0] ram_268; // @[vga.scala 14:20]
  reg [7:0] ram_269; // @[vga.scala 14:20]
  reg [7:0] ram_270; // @[vga.scala 14:20]
  reg [7:0] ram_271; // @[vga.scala 14:20]
  reg [7:0] ram_272; // @[vga.scala 14:20]
  reg [7:0] ram_273; // @[vga.scala 14:20]
  reg [7:0] ram_274; // @[vga.scala 14:20]
  reg [7:0] ram_275; // @[vga.scala 14:20]
  reg [7:0] ram_276; // @[vga.scala 14:20]
  reg [7:0] ram_277; // @[vga.scala 14:20]
  reg [7:0] ram_278; // @[vga.scala 14:20]
  reg [7:0] ram_279; // @[vga.scala 14:20]
  reg [7:0] ram_280; // @[vga.scala 14:20]
  reg [7:0] ram_281; // @[vga.scala 14:20]
  reg [7:0] ram_282; // @[vga.scala 14:20]
  reg [7:0] ram_283; // @[vga.scala 14:20]
  reg [7:0] ram_284; // @[vga.scala 14:20]
  reg [7:0] ram_285; // @[vga.scala 14:20]
  reg [7:0] ram_286; // @[vga.scala 14:20]
  reg [7:0] ram_287; // @[vga.scala 14:20]
  reg [7:0] ram_288; // @[vga.scala 14:20]
  reg [7:0] ram_289; // @[vga.scala 14:20]
  reg [7:0] ram_290; // @[vga.scala 14:20]
  reg [7:0] ram_291; // @[vga.scala 14:20]
  reg [7:0] ram_292; // @[vga.scala 14:20]
  reg [7:0] ram_293; // @[vga.scala 14:20]
  reg [7:0] ram_294; // @[vga.scala 14:20]
  reg [7:0] ram_295; // @[vga.scala 14:20]
  reg [7:0] ram_296; // @[vga.scala 14:20]
  reg [7:0] ram_297; // @[vga.scala 14:20]
  reg [7:0] ram_298; // @[vga.scala 14:20]
  reg [7:0] ram_299; // @[vga.scala 14:20]
  reg [7:0] ram_300; // @[vga.scala 14:20]
  reg [7:0] ram_301; // @[vga.scala 14:20]
  reg [7:0] ram_302; // @[vga.scala 14:20]
  reg [7:0] ram_303; // @[vga.scala 14:20]
  reg [7:0] ram_304; // @[vga.scala 14:20]
  reg [7:0] ram_305; // @[vga.scala 14:20]
  reg [7:0] ram_306; // @[vga.scala 14:20]
  reg [7:0] ram_307; // @[vga.scala 14:20]
  reg [7:0] ram_308; // @[vga.scala 14:20]
  reg [7:0] ram_309; // @[vga.scala 14:20]
  reg [7:0] ram_310; // @[vga.scala 14:20]
  reg [7:0] ram_311; // @[vga.scala 14:20]
  reg [7:0] ram_312; // @[vga.scala 14:20]
  reg [7:0] ram_313; // @[vga.scala 14:20]
  reg [7:0] ram_314; // @[vga.scala 14:20]
  reg [7:0] ram_315; // @[vga.scala 14:20]
  reg [7:0] ram_316; // @[vga.scala 14:20]
  reg [7:0] ram_317; // @[vga.scala 14:20]
  reg [7:0] ram_318; // @[vga.scala 14:20]
  reg [7:0] ram_319; // @[vga.scala 14:20]
  reg [7:0] ram_320; // @[vga.scala 14:20]
  reg [7:0] ram_321; // @[vga.scala 14:20]
  reg [7:0] ram_322; // @[vga.scala 14:20]
  reg [7:0] ram_323; // @[vga.scala 14:20]
  reg [7:0] ram_324; // @[vga.scala 14:20]
  reg [7:0] ram_325; // @[vga.scala 14:20]
  reg [7:0] ram_326; // @[vga.scala 14:20]
  reg [7:0] ram_327; // @[vga.scala 14:20]
  reg [7:0] ram_328; // @[vga.scala 14:20]
  reg [7:0] ram_329; // @[vga.scala 14:20]
  reg [7:0] ram_330; // @[vga.scala 14:20]
  reg [7:0] ram_331; // @[vga.scala 14:20]
  reg [7:0] ram_332; // @[vga.scala 14:20]
  reg [7:0] ram_333; // @[vga.scala 14:20]
  reg [7:0] ram_334; // @[vga.scala 14:20]
  reg [7:0] ram_335; // @[vga.scala 14:20]
  reg [7:0] ram_336; // @[vga.scala 14:20]
  reg [7:0] ram_337; // @[vga.scala 14:20]
  reg [7:0] ram_338; // @[vga.scala 14:20]
  reg [7:0] ram_339; // @[vga.scala 14:20]
  reg [7:0] ram_340; // @[vga.scala 14:20]
  reg [7:0] ram_341; // @[vga.scala 14:20]
  reg [7:0] ram_342; // @[vga.scala 14:20]
  reg [7:0] ram_343; // @[vga.scala 14:20]
  reg [7:0] ram_344; // @[vga.scala 14:20]
  reg [7:0] ram_345; // @[vga.scala 14:20]
  reg [7:0] ram_346; // @[vga.scala 14:20]
  reg [7:0] ram_347; // @[vga.scala 14:20]
  reg [7:0] ram_348; // @[vga.scala 14:20]
  reg [7:0] ram_349; // @[vga.scala 14:20]
  reg [7:0] ram_350; // @[vga.scala 14:20]
  reg [7:0] ram_351; // @[vga.scala 14:20]
  reg [7:0] ram_352; // @[vga.scala 14:20]
  reg [7:0] ram_353; // @[vga.scala 14:20]
  reg [7:0] ram_354; // @[vga.scala 14:20]
  reg [7:0] ram_355; // @[vga.scala 14:20]
  reg [7:0] ram_356; // @[vga.scala 14:20]
  reg [7:0] ram_357; // @[vga.scala 14:20]
  reg [7:0] ram_358; // @[vga.scala 14:20]
  reg [7:0] ram_359; // @[vga.scala 14:20]
  reg [7:0] ram_360; // @[vga.scala 14:20]
  reg [7:0] ram_361; // @[vga.scala 14:20]
  reg [7:0] ram_362; // @[vga.scala 14:20]
  reg [7:0] ram_363; // @[vga.scala 14:20]
  reg [7:0] ram_364; // @[vga.scala 14:20]
  reg [7:0] ram_365; // @[vga.scala 14:20]
  reg [7:0] ram_366; // @[vga.scala 14:20]
  reg [7:0] ram_367; // @[vga.scala 14:20]
  reg [7:0] ram_368; // @[vga.scala 14:20]
  reg [7:0] ram_369; // @[vga.scala 14:20]
  reg [7:0] ram_370; // @[vga.scala 14:20]
  reg [7:0] ram_371; // @[vga.scala 14:20]
  reg [7:0] ram_372; // @[vga.scala 14:20]
  reg [7:0] ram_373; // @[vga.scala 14:20]
  reg [7:0] ram_374; // @[vga.scala 14:20]
  reg [7:0] ram_375; // @[vga.scala 14:20]
  reg [7:0] ram_376; // @[vga.scala 14:20]
  reg [7:0] ram_377; // @[vga.scala 14:20]
  reg [7:0] ram_378; // @[vga.scala 14:20]
  reg [7:0] ram_379; // @[vga.scala 14:20]
  reg [7:0] ram_380; // @[vga.scala 14:20]
  reg [7:0] ram_381; // @[vga.scala 14:20]
  reg [7:0] ram_382; // @[vga.scala 14:20]
  reg [7:0] ram_383; // @[vga.scala 14:20]
  reg [7:0] ram_384; // @[vga.scala 14:20]
  reg [7:0] ram_385; // @[vga.scala 14:20]
  reg [7:0] ram_386; // @[vga.scala 14:20]
  reg [7:0] ram_387; // @[vga.scala 14:20]
  reg [7:0] ram_388; // @[vga.scala 14:20]
  reg [7:0] ram_389; // @[vga.scala 14:20]
  reg [7:0] ram_390; // @[vga.scala 14:20]
  reg [7:0] ram_391; // @[vga.scala 14:20]
  reg [7:0] ram_392; // @[vga.scala 14:20]
  reg [7:0] ram_393; // @[vga.scala 14:20]
  reg [7:0] ram_394; // @[vga.scala 14:20]
  reg [7:0] ram_395; // @[vga.scala 14:20]
  reg [7:0] ram_396; // @[vga.scala 14:20]
  reg [7:0] ram_397; // @[vga.scala 14:20]
  reg [7:0] ram_398; // @[vga.scala 14:20]
  reg [7:0] ram_399; // @[vga.scala 14:20]
  reg [7:0] ram_400; // @[vga.scala 14:20]
  reg [7:0] ram_401; // @[vga.scala 14:20]
  reg [7:0] ram_402; // @[vga.scala 14:20]
  reg [7:0] ram_403; // @[vga.scala 14:20]
  reg [7:0] ram_404; // @[vga.scala 14:20]
  reg [7:0] ram_405; // @[vga.scala 14:20]
  reg [7:0] ram_406; // @[vga.scala 14:20]
  reg [7:0] ram_407; // @[vga.scala 14:20]
  reg [7:0] ram_408; // @[vga.scala 14:20]
  reg [7:0] ram_409; // @[vga.scala 14:20]
  reg [7:0] ram_410; // @[vga.scala 14:20]
  reg [7:0] ram_411; // @[vga.scala 14:20]
  reg [7:0] ram_412; // @[vga.scala 14:20]
  reg [7:0] ram_413; // @[vga.scala 14:20]
  reg [7:0] ram_414; // @[vga.scala 14:20]
  reg [7:0] ram_415; // @[vga.scala 14:20]
  reg [7:0] ram_416; // @[vga.scala 14:20]
  reg [7:0] ram_417; // @[vga.scala 14:20]
  reg [7:0] ram_418; // @[vga.scala 14:20]
  reg [7:0] ram_419; // @[vga.scala 14:20]
  reg [7:0] ram_420; // @[vga.scala 14:20]
  reg [7:0] ram_421; // @[vga.scala 14:20]
  reg [7:0] ram_422; // @[vga.scala 14:20]
  reg [7:0] ram_423; // @[vga.scala 14:20]
  reg [7:0] ram_424; // @[vga.scala 14:20]
  reg [7:0] ram_425; // @[vga.scala 14:20]
  reg [7:0] ram_426; // @[vga.scala 14:20]
  reg [7:0] ram_427; // @[vga.scala 14:20]
  reg [7:0] ram_428; // @[vga.scala 14:20]
  reg [7:0] ram_429; // @[vga.scala 14:20]
  reg [7:0] ram_430; // @[vga.scala 14:20]
  reg [7:0] ram_431; // @[vga.scala 14:20]
  reg [7:0] ram_432; // @[vga.scala 14:20]
  reg [7:0] ram_433; // @[vga.scala 14:20]
  reg [7:0] ram_434; // @[vga.scala 14:20]
  reg [7:0] ram_435; // @[vga.scala 14:20]
  reg [7:0] ram_436; // @[vga.scala 14:20]
  reg [7:0] ram_437; // @[vga.scala 14:20]
  reg [7:0] ram_438; // @[vga.scala 14:20]
  reg [7:0] ram_439; // @[vga.scala 14:20]
  reg [7:0] ram_440; // @[vga.scala 14:20]
  reg [7:0] ram_441; // @[vga.scala 14:20]
  reg [7:0] ram_442; // @[vga.scala 14:20]
  reg [7:0] ram_443; // @[vga.scala 14:20]
  reg [7:0] ram_444; // @[vga.scala 14:20]
  reg [7:0] ram_445; // @[vga.scala 14:20]
  reg [7:0] ram_446; // @[vga.scala 14:20]
  reg [7:0] ram_447; // @[vga.scala 14:20]
  reg [7:0] ram_448; // @[vga.scala 14:20]
  reg [7:0] ram_449; // @[vga.scala 14:20]
  reg [7:0] ram_450; // @[vga.scala 14:20]
  reg [7:0] ram_451; // @[vga.scala 14:20]
  reg [7:0] ram_452; // @[vga.scala 14:20]
  reg [7:0] ram_453; // @[vga.scala 14:20]
  reg [7:0] ram_454; // @[vga.scala 14:20]
  reg [7:0] ram_455; // @[vga.scala 14:20]
  reg [7:0] ram_456; // @[vga.scala 14:20]
  reg [7:0] ram_457; // @[vga.scala 14:20]
  reg [7:0] ram_458; // @[vga.scala 14:20]
  reg [7:0] ram_459; // @[vga.scala 14:20]
  reg [7:0] ram_460; // @[vga.scala 14:20]
  reg [7:0] ram_461; // @[vga.scala 14:20]
  reg [7:0] ram_462; // @[vga.scala 14:20]
  reg [7:0] ram_463; // @[vga.scala 14:20]
  reg [7:0] ram_464; // @[vga.scala 14:20]
  reg [7:0] ram_465; // @[vga.scala 14:20]
  reg [7:0] ram_466; // @[vga.scala 14:20]
  reg [7:0] ram_467; // @[vga.scala 14:20]
  reg [7:0] ram_468; // @[vga.scala 14:20]
  reg [7:0] ram_469; // @[vga.scala 14:20]
  reg [7:0] ram_470; // @[vga.scala 14:20]
  reg [7:0] ram_471; // @[vga.scala 14:20]
  reg [7:0] ram_472; // @[vga.scala 14:20]
  reg [7:0] ram_473; // @[vga.scala 14:20]
  reg [7:0] ram_474; // @[vga.scala 14:20]
  reg [7:0] ram_475; // @[vga.scala 14:20]
  reg [7:0] ram_476; // @[vga.scala 14:20]
  reg [7:0] ram_477; // @[vga.scala 14:20]
  reg [7:0] ram_478; // @[vga.scala 14:20]
  reg [7:0] ram_479; // @[vga.scala 14:20]
  reg [7:0] ram_480; // @[vga.scala 14:20]
  reg [7:0] ram_481; // @[vga.scala 14:20]
  reg [7:0] ram_482; // @[vga.scala 14:20]
  reg [7:0] ram_483; // @[vga.scala 14:20]
  reg [7:0] ram_484; // @[vga.scala 14:20]
  reg [7:0] ram_485; // @[vga.scala 14:20]
  reg [7:0] ram_486; // @[vga.scala 14:20]
  reg [7:0] ram_487; // @[vga.scala 14:20]
  reg [7:0] ram_488; // @[vga.scala 14:20]
  reg [7:0] ram_489; // @[vga.scala 14:20]
  reg [7:0] ram_490; // @[vga.scala 14:20]
  reg [7:0] ram_491; // @[vga.scala 14:20]
  reg [7:0] ram_492; // @[vga.scala 14:20]
  reg [7:0] ram_493; // @[vga.scala 14:20]
  reg [7:0] ram_494; // @[vga.scala 14:20]
  reg [7:0] ram_495; // @[vga.scala 14:20]
  reg [7:0] ram_496; // @[vga.scala 14:20]
  reg [7:0] ram_497; // @[vga.scala 14:20]
  reg [7:0] ram_498; // @[vga.scala 14:20]
  reg [7:0] ram_499; // @[vga.scala 14:20]
  reg [7:0] ram_500; // @[vga.scala 14:20]
  reg [7:0] ram_501; // @[vga.scala 14:20]
  reg [7:0] ram_502; // @[vga.scala 14:20]
  reg [7:0] ram_503; // @[vga.scala 14:20]
  reg [7:0] ram_504; // @[vga.scala 14:20]
  reg [7:0] ram_505; // @[vga.scala 14:20]
  reg [7:0] ram_506; // @[vga.scala 14:20]
  reg [7:0] ram_507; // @[vga.scala 14:20]
  reg [7:0] ram_508; // @[vga.scala 14:20]
  reg [7:0] ram_509; // @[vga.scala 14:20]
  reg [7:0] ram_510; // @[vga.scala 14:20]
  reg [7:0] ram_511; // @[vga.scala 14:20]
  reg [7:0] ram_512; // @[vga.scala 14:20]
  reg [7:0] ram_513; // @[vga.scala 14:20]
  reg [7:0] ram_514; // @[vga.scala 14:20]
  reg [7:0] ram_515; // @[vga.scala 14:20]
  reg [7:0] ram_516; // @[vga.scala 14:20]
  reg [7:0] ram_517; // @[vga.scala 14:20]
  reg [7:0] ram_518; // @[vga.scala 14:20]
  reg [7:0] ram_519; // @[vga.scala 14:20]
  reg [7:0] ram_520; // @[vga.scala 14:20]
  reg [7:0] ram_521; // @[vga.scala 14:20]
  reg [7:0] ram_522; // @[vga.scala 14:20]
  reg [7:0] ram_523; // @[vga.scala 14:20]
  reg [7:0] ram_524; // @[vga.scala 14:20]
  reg [7:0] ram_525; // @[vga.scala 14:20]
  reg [7:0] ram_526; // @[vga.scala 14:20]
  reg [7:0] ram_527; // @[vga.scala 14:20]
  reg [7:0] ram_528; // @[vga.scala 14:20]
  reg [7:0] ram_529; // @[vga.scala 14:20]
  reg [7:0] ram_530; // @[vga.scala 14:20]
  reg [7:0] ram_531; // @[vga.scala 14:20]
  reg [7:0] ram_532; // @[vga.scala 14:20]
  reg [7:0] ram_533; // @[vga.scala 14:20]
  reg [7:0] ram_534; // @[vga.scala 14:20]
  reg [7:0] ram_535; // @[vga.scala 14:20]
  reg [7:0] ram_536; // @[vga.scala 14:20]
  reg [7:0] ram_537; // @[vga.scala 14:20]
  reg [7:0] ram_538; // @[vga.scala 14:20]
  reg [7:0] ram_539; // @[vga.scala 14:20]
  reg [7:0] ram_540; // @[vga.scala 14:20]
  reg [7:0] ram_541; // @[vga.scala 14:20]
  reg [7:0] ram_542; // @[vga.scala 14:20]
  reg [7:0] ram_543; // @[vga.scala 14:20]
  reg [7:0] ram_544; // @[vga.scala 14:20]
  reg [7:0] ram_545; // @[vga.scala 14:20]
  reg [7:0] ram_546; // @[vga.scala 14:20]
  reg [7:0] ram_547; // @[vga.scala 14:20]
  reg [7:0] ram_548; // @[vga.scala 14:20]
  reg [7:0] ram_549; // @[vga.scala 14:20]
  reg [7:0] ram_550; // @[vga.scala 14:20]
  reg [7:0] ram_551; // @[vga.scala 14:20]
  reg [7:0] ram_552; // @[vga.scala 14:20]
  reg [7:0] ram_553; // @[vga.scala 14:20]
  reg [7:0] ram_554; // @[vga.scala 14:20]
  reg [7:0] ram_555; // @[vga.scala 14:20]
  reg [7:0] ram_556; // @[vga.scala 14:20]
  reg [7:0] ram_557; // @[vga.scala 14:20]
  reg [7:0] ram_558; // @[vga.scala 14:20]
  reg [7:0] ram_559; // @[vga.scala 14:20]
  reg [7:0] ram_560; // @[vga.scala 14:20]
  reg [7:0] ram_561; // @[vga.scala 14:20]
  reg [7:0] ram_562; // @[vga.scala 14:20]
  reg [7:0] ram_563; // @[vga.scala 14:20]
  reg [7:0] ram_564; // @[vga.scala 14:20]
  reg [7:0] ram_565; // @[vga.scala 14:20]
  reg [7:0] ram_566; // @[vga.scala 14:20]
  reg [7:0] ram_567; // @[vga.scala 14:20]
  reg [7:0] ram_568; // @[vga.scala 14:20]
  reg [7:0] ram_569; // @[vga.scala 14:20]
  reg [7:0] ram_570; // @[vga.scala 14:20]
  reg [7:0] ram_571; // @[vga.scala 14:20]
  reg [7:0] ram_572; // @[vga.scala 14:20]
  reg [7:0] ram_573; // @[vga.scala 14:20]
  reg [7:0] ram_574; // @[vga.scala 14:20]
  reg [7:0] ram_575; // @[vga.scala 14:20]
  reg [7:0] ram_576; // @[vga.scala 14:20]
  reg [7:0] ram_577; // @[vga.scala 14:20]
  reg [7:0] ram_578; // @[vga.scala 14:20]
  reg [7:0] ram_579; // @[vga.scala 14:20]
  reg [7:0] ram_580; // @[vga.scala 14:20]
  reg [7:0] ram_581; // @[vga.scala 14:20]
  reg [7:0] ram_582; // @[vga.scala 14:20]
  reg [7:0] ram_583; // @[vga.scala 14:20]
  reg [7:0] ram_584; // @[vga.scala 14:20]
  reg [7:0] ram_585; // @[vga.scala 14:20]
  reg [7:0] ram_586; // @[vga.scala 14:20]
  reg [7:0] ram_587; // @[vga.scala 14:20]
  reg [7:0] ram_588; // @[vga.scala 14:20]
  reg [7:0] ram_589; // @[vga.scala 14:20]
  reg [7:0] ram_590; // @[vga.scala 14:20]
  reg [7:0] ram_591; // @[vga.scala 14:20]
  reg [7:0] ram_592; // @[vga.scala 14:20]
  reg [7:0] ram_593; // @[vga.scala 14:20]
  reg [7:0] ram_594; // @[vga.scala 14:20]
  reg [7:0] ram_595; // @[vga.scala 14:20]
  reg [7:0] ram_596; // @[vga.scala 14:20]
  reg [7:0] ram_597; // @[vga.scala 14:20]
  reg [7:0] ram_598; // @[vga.scala 14:20]
  reg [7:0] ram_599; // @[vga.scala 14:20]
  reg [7:0] ram_600; // @[vga.scala 14:20]
  reg [7:0] ram_601; // @[vga.scala 14:20]
  reg [7:0] ram_602; // @[vga.scala 14:20]
  reg [7:0] ram_603; // @[vga.scala 14:20]
  reg [7:0] ram_604; // @[vga.scala 14:20]
  reg [7:0] ram_605; // @[vga.scala 14:20]
  reg [7:0] ram_606; // @[vga.scala 14:20]
  reg [7:0] ram_607; // @[vga.scala 14:20]
  reg [7:0] ram_608; // @[vga.scala 14:20]
  reg [7:0] ram_609; // @[vga.scala 14:20]
  reg [7:0] ram_610; // @[vga.scala 14:20]
  reg [7:0] ram_611; // @[vga.scala 14:20]
  reg [7:0] ram_612; // @[vga.scala 14:20]
  reg [7:0] ram_613; // @[vga.scala 14:20]
  reg [7:0] ram_614; // @[vga.scala 14:20]
  reg [7:0] ram_615; // @[vga.scala 14:20]
  reg [7:0] ram_616; // @[vga.scala 14:20]
  reg [7:0] ram_617; // @[vga.scala 14:20]
  reg [7:0] ram_618; // @[vga.scala 14:20]
  reg [7:0] ram_619; // @[vga.scala 14:20]
  reg [7:0] ram_620; // @[vga.scala 14:20]
  reg [7:0] ram_621; // @[vga.scala 14:20]
  reg [7:0] ram_622; // @[vga.scala 14:20]
  reg [7:0] ram_623; // @[vga.scala 14:20]
  reg [7:0] ram_624; // @[vga.scala 14:20]
  reg [7:0] ram_625; // @[vga.scala 14:20]
  reg [7:0] ram_626; // @[vga.scala 14:20]
  reg [7:0] ram_627; // @[vga.scala 14:20]
  reg [7:0] ram_628; // @[vga.scala 14:20]
  reg [7:0] ram_629; // @[vga.scala 14:20]
  reg [7:0] ram_630; // @[vga.scala 14:20]
  reg [7:0] ram_631; // @[vga.scala 14:20]
  reg [7:0] ram_632; // @[vga.scala 14:20]
  reg [7:0] ram_633; // @[vga.scala 14:20]
  reg [7:0] ram_634; // @[vga.scala 14:20]
  reg [7:0] ram_635; // @[vga.scala 14:20]
  reg [7:0] ram_636; // @[vga.scala 14:20]
  reg [7:0] ram_637; // @[vga.scala 14:20]
  reg [7:0] ram_638; // @[vga.scala 14:20]
  reg [7:0] ram_639; // @[vga.scala 14:20]
  reg [7:0] ram_640; // @[vga.scala 14:20]
  reg [7:0] ram_641; // @[vga.scala 14:20]
  reg [7:0] ram_642; // @[vga.scala 14:20]
  reg [7:0] ram_643; // @[vga.scala 14:20]
  reg [7:0] ram_644; // @[vga.scala 14:20]
  reg [7:0] ram_645; // @[vga.scala 14:20]
  reg [7:0] ram_646; // @[vga.scala 14:20]
  reg [7:0] ram_647; // @[vga.scala 14:20]
  reg [7:0] ram_648; // @[vga.scala 14:20]
  reg [7:0] ram_649; // @[vga.scala 14:20]
  reg [7:0] ram_650; // @[vga.scala 14:20]
  reg [7:0] ram_651; // @[vga.scala 14:20]
  reg [7:0] ram_652; // @[vga.scala 14:20]
  reg [7:0] ram_653; // @[vga.scala 14:20]
  reg [7:0] ram_654; // @[vga.scala 14:20]
  reg [7:0] ram_655; // @[vga.scala 14:20]
  reg [7:0] ram_656; // @[vga.scala 14:20]
  reg [7:0] ram_657; // @[vga.scala 14:20]
  reg [7:0] ram_658; // @[vga.scala 14:20]
  reg [7:0] ram_659; // @[vga.scala 14:20]
  reg [7:0] ram_660; // @[vga.scala 14:20]
  reg [7:0] ram_661; // @[vga.scala 14:20]
  reg [7:0] ram_662; // @[vga.scala 14:20]
  reg [7:0] ram_663; // @[vga.scala 14:20]
  reg [7:0] ram_664; // @[vga.scala 14:20]
  reg [7:0] ram_665; // @[vga.scala 14:20]
  reg [7:0] ram_666; // @[vga.scala 14:20]
  reg [7:0] ram_667; // @[vga.scala 14:20]
  reg [7:0] ram_668; // @[vga.scala 14:20]
  reg [7:0] ram_669; // @[vga.scala 14:20]
  reg [7:0] ram_670; // @[vga.scala 14:20]
  reg [7:0] ram_671; // @[vga.scala 14:20]
  reg [7:0] ram_672; // @[vga.scala 14:20]
  reg [7:0] ram_673; // @[vga.scala 14:20]
  reg [7:0] ram_674; // @[vga.scala 14:20]
  reg [7:0] ram_675; // @[vga.scala 14:20]
  reg [7:0] ram_676; // @[vga.scala 14:20]
  reg [7:0] ram_677; // @[vga.scala 14:20]
  reg [7:0] ram_678; // @[vga.scala 14:20]
  reg [7:0] ram_679; // @[vga.scala 14:20]
  reg [7:0] ram_680; // @[vga.scala 14:20]
  reg [7:0] ram_681; // @[vga.scala 14:20]
  reg [7:0] ram_682; // @[vga.scala 14:20]
  reg [7:0] ram_683; // @[vga.scala 14:20]
  reg [7:0] ram_684; // @[vga.scala 14:20]
  reg [7:0] ram_685; // @[vga.scala 14:20]
  reg [7:0] ram_686; // @[vga.scala 14:20]
  reg [7:0] ram_687; // @[vga.scala 14:20]
  reg [7:0] ram_688; // @[vga.scala 14:20]
  reg [7:0] ram_689; // @[vga.scala 14:20]
  reg [7:0] ram_690; // @[vga.scala 14:20]
  reg [7:0] ram_691; // @[vga.scala 14:20]
  reg [7:0] ram_692; // @[vga.scala 14:20]
  reg [7:0] ram_693; // @[vga.scala 14:20]
  reg [7:0] ram_694; // @[vga.scala 14:20]
  reg [7:0] ram_695; // @[vga.scala 14:20]
  reg [7:0] ram_696; // @[vga.scala 14:20]
  reg [7:0] ram_697; // @[vga.scala 14:20]
  reg [7:0] ram_698; // @[vga.scala 14:20]
  reg [7:0] ram_699; // @[vga.scala 14:20]
  reg [7:0] ram_700; // @[vga.scala 14:20]
  reg [7:0] ram_701; // @[vga.scala 14:20]
  reg [7:0] ram_702; // @[vga.scala 14:20]
  reg [7:0] ram_703; // @[vga.scala 14:20]
  reg [7:0] ram_704; // @[vga.scala 14:20]
  reg [7:0] ram_705; // @[vga.scala 14:20]
  reg [7:0] ram_706; // @[vga.scala 14:20]
  reg [7:0] ram_707; // @[vga.scala 14:20]
  reg [7:0] ram_708; // @[vga.scala 14:20]
  reg [7:0] ram_709; // @[vga.scala 14:20]
  reg [7:0] ram_710; // @[vga.scala 14:20]
  reg [7:0] ram_711; // @[vga.scala 14:20]
  reg [7:0] ram_712; // @[vga.scala 14:20]
  reg [7:0] ram_713; // @[vga.scala 14:20]
  reg [7:0] ram_714; // @[vga.scala 14:20]
  reg [7:0] ram_715; // @[vga.scala 14:20]
  reg [7:0] ram_716; // @[vga.scala 14:20]
  reg [7:0] ram_717; // @[vga.scala 14:20]
  reg [7:0] ram_718; // @[vga.scala 14:20]
  reg [7:0] ram_719; // @[vga.scala 14:20]
  reg [7:0] ram_720; // @[vga.scala 14:20]
  reg [7:0] ram_721; // @[vga.scala 14:20]
  reg [7:0] ram_722; // @[vga.scala 14:20]
  reg [7:0] ram_723; // @[vga.scala 14:20]
  reg [7:0] ram_724; // @[vga.scala 14:20]
  reg [7:0] ram_725; // @[vga.scala 14:20]
  reg [7:0] ram_726; // @[vga.scala 14:20]
  reg [7:0] ram_727; // @[vga.scala 14:20]
  reg [7:0] ram_728; // @[vga.scala 14:20]
  reg [7:0] ram_729; // @[vga.scala 14:20]
  reg [7:0] ram_730; // @[vga.scala 14:20]
  reg [7:0] ram_731; // @[vga.scala 14:20]
  reg [7:0] ram_732; // @[vga.scala 14:20]
  reg [7:0] ram_733; // @[vga.scala 14:20]
  reg [7:0] ram_734; // @[vga.scala 14:20]
  reg [7:0] ram_735; // @[vga.scala 14:20]
  reg [7:0] ram_736; // @[vga.scala 14:20]
  reg [7:0] ram_737; // @[vga.scala 14:20]
  reg [7:0] ram_738; // @[vga.scala 14:20]
  reg [7:0] ram_739; // @[vga.scala 14:20]
  reg [7:0] ram_740; // @[vga.scala 14:20]
  reg [7:0] ram_741; // @[vga.scala 14:20]
  reg [7:0] ram_742; // @[vga.scala 14:20]
  reg [7:0] ram_743; // @[vga.scala 14:20]
  reg [7:0] ram_744; // @[vga.scala 14:20]
  reg [7:0] ram_745; // @[vga.scala 14:20]
  reg [7:0] ram_746; // @[vga.scala 14:20]
  reg [7:0] ram_747; // @[vga.scala 14:20]
  reg [7:0] ram_748; // @[vga.scala 14:20]
  reg [7:0] ram_749; // @[vga.scala 14:20]
  reg [7:0] ram_750; // @[vga.scala 14:20]
  reg [7:0] ram_751; // @[vga.scala 14:20]
  reg [7:0] ram_752; // @[vga.scala 14:20]
  reg [7:0] ram_753; // @[vga.scala 14:20]
  reg [7:0] ram_754; // @[vga.scala 14:20]
  reg [7:0] ram_755; // @[vga.scala 14:20]
  reg [7:0] ram_756; // @[vga.scala 14:20]
  reg [7:0] ram_757; // @[vga.scala 14:20]
  reg [7:0] ram_758; // @[vga.scala 14:20]
  reg [7:0] ram_759; // @[vga.scala 14:20]
  reg [7:0] ram_760; // @[vga.scala 14:20]
  reg [7:0] ram_761; // @[vga.scala 14:20]
  reg [7:0] ram_762; // @[vga.scala 14:20]
  reg [7:0] ram_763; // @[vga.scala 14:20]
  reg [7:0] ram_764; // @[vga.scala 14:20]
  reg [7:0] ram_765; // @[vga.scala 14:20]
  reg [7:0] ram_766; // @[vga.scala 14:20]
  reg [7:0] ram_767; // @[vga.scala 14:20]
  reg [7:0] ram_768; // @[vga.scala 14:20]
  reg [7:0] ram_769; // @[vga.scala 14:20]
  reg [7:0] ram_770; // @[vga.scala 14:20]
  reg [7:0] ram_771; // @[vga.scala 14:20]
  reg [7:0] ram_772; // @[vga.scala 14:20]
  reg [7:0] ram_773; // @[vga.scala 14:20]
  reg [7:0] ram_774; // @[vga.scala 14:20]
  reg [7:0] ram_775; // @[vga.scala 14:20]
  reg [7:0] ram_776; // @[vga.scala 14:20]
  reg [7:0] ram_777; // @[vga.scala 14:20]
  reg [7:0] ram_778; // @[vga.scala 14:20]
  reg [7:0] ram_779; // @[vga.scala 14:20]
  reg [7:0] ram_780; // @[vga.scala 14:20]
  reg [7:0] ram_781; // @[vga.scala 14:20]
  reg [7:0] ram_782; // @[vga.scala 14:20]
  reg [7:0] ram_783; // @[vga.scala 14:20]
  reg [7:0] ram_784; // @[vga.scala 14:20]
  reg [7:0] ram_785; // @[vga.scala 14:20]
  reg [7:0] ram_786; // @[vga.scala 14:20]
  reg [7:0] ram_787; // @[vga.scala 14:20]
  reg [7:0] ram_788; // @[vga.scala 14:20]
  reg [7:0] ram_789; // @[vga.scala 14:20]
  reg [7:0] ram_790; // @[vga.scala 14:20]
  reg [7:0] ram_791; // @[vga.scala 14:20]
  reg [7:0] ram_792; // @[vga.scala 14:20]
  reg [7:0] ram_793; // @[vga.scala 14:20]
  reg [7:0] ram_794; // @[vga.scala 14:20]
  reg [7:0] ram_795; // @[vga.scala 14:20]
  reg [7:0] ram_796; // @[vga.scala 14:20]
  reg [7:0] ram_797; // @[vga.scala 14:20]
  reg [7:0] ram_798; // @[vga.scala 14:20]
  reg [7:0] ram_799; // @[vga.scala 14:20]
  reg [7:0] ram_800; // @[vga.scala 14:20]
  reg [7:0] ram_801; // @[vga.scala 14:20]
  reg [7:0] ram_802; // @[vga.scala 14:20]
  reg [7:0] ram_803; // @[vga.scala 14:20]
  reg [7:0] ram_804; // @[vga.scala 14:20]
  reg [7:0] ram_805; // @[vga.scala 14:20]
  reg [7:0] ram_806; // @[vga.scala 14:20]
  reg [7:0] ram_807; // @[vga.scala 14:20]
  reg [7:0] ram_808; // @[vga.scala 14:20]
  reg [7:0] ram_809; // @[vga.scala 14:20]
  reg [7:0] ram_810; // @[vga.scala 14:20]
  reg [7:0] ram_811; // @[vga.scala 14:20]
  reg [7:0] ram_812; // @[vga.scala 14:20]
  reg [7:0] ram_813; // @[vga.scala 14:20]
  reg [7:0] ram_814; // @[vga.scala 14:20]
  reg [7:0] ram_815; // @[vga.scala 14:20]
  reg [7:0] ram_816; // @[vga.scala 14:20]
  reg [7:0] ram_817; // @[vga.scala 14:20]
  reg [7:0] ram_818; // @[vga.scala 14:20]
  reg [7:0] ram_819; // @[vga.scala 14:20]
  reg [7:0] ram_820; // @[vga.scala 14:20]
  reg [7:0] ram_821; // @[vga.scala 14:20]
  reg [7:0] ram_822; // @[vga.scala 14:20]
  reg [7:0] ram_823; // @[vga.scala 14:20]
  reg [7:0] ram_824; // @[vga.scala 14:20]
  reg [7:0] ram_825; // @[vga.scala 14:20]
  reg [7:0] ram_826; // @[vga.scala 14:20]
  reg [7:0] ram_827; // @[vga.scala 14:20]
  reg [7:0] ram_828; // @[vga.scala 14:20]
  reg [7:0] ram_829; // @[vga.scala 14:20]
  reg [7:0] ram_830; // @[vga.scala 14:20]
  reg [7:0] ram_831; // @[vga.scala 14:20]
  reg [7:0] ram_832; // @[vga.scala 14:20]
  reg [7:0] ram_833; // @[vga.scala 14:20]
  reg [7:0] ram_834; // @[vga.scala 14:20]
  reg [7:0] ram_835; // @[vga.scala 14:20]
  reg [7:0] ram_836; // @[vga.scala 14:20]
  reg [7:0] ram_837; // @[vga.scala 14:20]
  reg [7:0] ram_838; // @[vga.scala 14:20]
  reg [7:0] ram_839; // @[vga.scala 14:20]
  reg [7:0] ram_840; // @[vga.scala 14:20]
  reg [7:0] ram_841; // @[vga.scala 14:20]
  reg [7:0] ram_842; // @[vga.scala 14:20]
  reg [7:0] ram_843; // @[vga.scala 14:20]
  reg [7:0] ram_844; // @[vga.scala 14:20]
  reg [7:0] ram_845; // @[vga.scala 14:20]
  reg [7:0] ram_846; // @[vga.scala 14:20]
  reg [7:0] ram_847; // @[vga.scala 14:20]
  reg [7:0] ram_848; // @[vga.scala 14:20]
  reg [7:0] ram_849; // @[vga.scala 14:20]
  reg [7:0] ram_850; // @[vga.scala 14:20]
  reg [7:0] ram_851; // @[vga.scala 14:20]
  reg [7:0] ram_852; // @[vga.scala 14:20]
  reg [7:0] ram_853; // @[vga.scala 14:20]
  reg [7:0] ram_854; // @[vga.scala 14:20]
  reg [7:0] ram_855; // @[vga.scala 14:20]
  reg [7:0] ram_856; // @[vga.scala 14:20]
  reg [7:0] ram_857; // @[vga.scala 14:20]
  reg [7:0] ram_858; // @[vga.scala 14:20]
  reg [7:0] ram_859; // @[vga.scala 14:20]
  reg [7:0] ram_860; // @[vga.scala 14:20]
  reg [7:0] ram_861; // @[vga.scala 14:20]
  reg [7:0] ram_862; // @[vga.scala 14:20]
  reg [7:0] ram_863; // @[vga.scala 14:20]
  reg [7:0] ram_864; // @[vga.scala 14:20]
  reg [7:0] ram_865; // @[vga.scala 14:20]
  reg [7:0] ram_866; // @[vga.scala 14:20]
  reg [7:0] ram_867; // @[vga.scala 14:20]
  reg [7:0] ram_868; // @[vga.scala 14:20]
  reg [7:0] ram_869; // @[vga.scala 14:20]
  reg [7:0] ram_870; // @[vga.scala 14:20]
  reg [7:0] ram_871; // @[vga.scala 14:20]
  reg [7:0] ram_872; // @[vga.scala 14:20]
  reg [7:0] ram_873; // @[vga.scala 14:20]
  reg [7:0] ram_874; // @[vga.scala 14:20]
  reg [7:0] ram_875; // @[vga.scala 14:20]
  reg [7:0] ram_876; // @[vga.scala 14:20]
  reg [7:0] ram_877; // @[vga.scala 14:20]
  reg [7:0] ram_878; // @[vga.scala 14:20]
  reg [7:0] ram_879; // @[vga.scala 14:20]
  reg [7:0] ram_880; // @[vga.scala 14:20]
  reg [7:0] ram_881; // @[vga.scala 14:20]
  reg [7:0] ram_882; // @[vga.scala 14:20]
  reg [7:0] ram_883; // @[vga.scala 14:20]
  reg [7:0] ram_884; // @[vga.scala 14:20]
  reg [7:0] ram_885; // @[vga.scala 14:20]
  reg [7:0] ram_886; // @[vga.scala 14:20]
  reg [7:0] ram_887; // @[vga.scala 14:20]
  reg [7:0] ram_888; // @[vga.scala 14:20]
  reg [7:0] ram_889; // @[vga.scala 14:20]
  reg [7:0] ram_890; // @[vga.scala 14:20]
  reg [7:0] ram_891; // @[vga.scala 14:20]
  reg [7:0] ram_892; // @[vga.scala 14:20]
  reg [7:0] ram_893; // @[vga.scala 14:20]
  reg [7:0] ram_894; // @[vga.scala 14:20]
  reg [7:0] ram_895; // @[vga.scala 14:20]
  reg [7:0] ram_896; // @[vga.scala 14:20]
  reg [7:0] ram_897; // @[vga.scala 14:20]
  reg [7:0] ram_898; // @[vga.scala 14:20]
  reg [7:0] ram_899; // @[vga.scala 14:20]
  reg [7:0] ram_900; // @[vga.scala 14:20]
  reg [7:0] ram_901; // @[vga.scala 14:20]
  reg [7:0] ram_902; // @[vga.scala 14:20]
  reg [7:0] ram_903; // @[vga.scala 14:20]
  reg [7:0] ram_904; // @[vga.scala 14:20]
  reg [7:0] ram_905; // @[vga.scala 14:20]
  reg [7:0] ram_906; // @[vga.scala 14:20]
  reg [7:0] ram_907; // @[vga.scala 14:20]
  reg [7:0] ram_908; // @[vga.scala 14:20]
  reg [7:0] ram_909; // @[vga.scala 14:20]
  reg [7:0] ram_910; // @[vga.scala 14:20]
  reg [7:0] ram_911; // @[vga.scala 14:20]
  reg [7:0] ram_912; // @[vga.scala 14:20]
  reg [7:0] ram_913; // @[vga.scala 14:20]
  reg [7:0] ram_914; // @[vga.scala 14:20]
  reg [7:0] ram_915; // @[vga.scala 14:20]
  reg [7:0] ram_916; // @[vga.scala 14:20]
  reg [7:0] ram_917; // @[vga.scala 14:20]
  reg [7:0] ram_918; // @[vga.scala 14:20]
  reg [7:0] ram_919; // @[vga.scala 14:20]
  reg [7:0] ram_920; // @[vga.scala 14:20]
  reg [7:0] ram_921; // @[vga.scala 14:20]
  reg [7:0] ram_922; // @[vga.scala 14:20]
  reg [7:0] ram_923; // @[vga.scala 14:20]
  reg [7:0] ram_924; // @[vga.scala 14:20]
  reg [7:0] ram_925; // @[vga.scala 14:20]
  reg [7:0] ram_926; // @[vga.scala 14:20]
  reg [7:0] ram_927; // @[vga.scala 14:20]
  reg [7:0] ram_928; // @[vga.scala 14:20]
  reg [7:0] ram_929; // @[vga.scala 14:20]
  reg [7:0] ram_930; // @[vga.scala 14:20]
  reg [7:0] ram_931; // @[vga.scala 14:20]
  reg [7:0] ram_932; // @[vga.scala 14:20]
  reg [7:0] ram_933; // @[vga.scala 14:20]
  reg [7:0] ram_934; // @[vga.scala 14:20]
  reg [7:0] ram_935; // @[vga.scala 14:20]
  reg [7:0] ram_936; // @[vga.scala 14:20]
  reg [7:0] ram_937; // @[vga.scala 14:20]
  reg [7:0] ram_938; // @[vga.scala 14:20]
  reg [7:0] ram_939; // @[vga.scala 14:20]
  reg [7:0] ram_940; // @[vga.scala 14:20]
  reg [7:0] ram_941; // @[vga.scala 14:20]
  reg [7:0] ram_942; // @[vga.scala 14:20]
  reg [7:0] ram_943; // @[vga.scala 14:20]
  reg [7:0] ram_944; // @[vga.scala 14:20]
  reg [7:0] ram_945; // @[vga.scala 14:20]
  reg [7:0] ram_946; // @[vga.scala 14:20]
  reg [7:0] ram_947; // @[vga.scala 14:20]
  reg [7:0] ram_948; // @[vga.scala 14:20]
  reg [7:0] ram_949; // @[vga.scala 14:20]
  reg [7:0] ram_950; // @[vga.scala 14:20]
  reg [7:0] ram_951; // @[vga.scala 14:20]
  reg [7:0] ram_952; // @[vga.scala 14:20]
  reg [7:0] ram_953; // @[vga.scala 14:20]
  reg [7:0] ram_954; // @[vga.scala 14:20]
  reg [7:0] ram_955; // @[vga.scala 14:20]
  reg [7:0] ram_956; // @[vga.scala 14:20]
  reg [7:0] ram_957; // @[vga.scala 14:20]
  reg [7:0] ram_958; // @[vga.scala 14:20]
  reg [7:0] ram_959; // @[vga.scala 14:20]
  reg [7:0] ram_960; // @[vga.scala 14:20]
  reg [7:0] ram_961; // @[vga.scala 14:20]
  reg [7:0] ram_962; // @[vga.scala 14:20]
  reg [7:0] ram_963; // @[vga.scala 14:20]
  reg [7:0] ram_964; // @[vga.scala 14:20]
  reg [7:0] ram_965; // @[vga.scala 14:20]
  reg [7:0] ram_966; // @[vga.scala 14:20]
  reg [7:0] ram_967; // @[vga.scala 14:20]
  reg [7:0] ram_968; // @[vga.scala 14:20]
  reg [7:0] ram_969; // @[vga.scala 14:20]
  reg [7:0] ram_970; // @[vga.scala 14:20]
  reg [7:0] ram_971; // @[vga.scala 14:20]
  reg [7:0] ram_972; // @[vga.scala 14:20]
  reg [7:0] ram_973; // @[vga.scala 14:20]
  reg [7:0] ram_974; // @[vga.scala 14:20]
  reg [7:0] ram_975; // @[vga.scala 14:20]
  reg [7:0] ram_976; // @[vga.scala 14:20]
  reg [7:0] ram_977; // @[vga.scala 14:20]
  reg [7:0] ram_978; // @[vga.scala 14:20]
  reg [7:0] ram_979; // @[vga.scala 14:20]
  reg [7:0] ram_980; // @[vga.scala 14:20]
  reg [7:0] ram_981; // @[vga.scala 14:20]
  reg [7:0] ram_982; // @[vga.scala 14:20]
  reg [7:0] ram_983; // @[vga.scala 14:20]
  reg [7:0] ram_984; // @[vga.scala 14:20]
  reg [7:0] ram_985; // @[vga.scala 14:20]
  reg [7:0] ram_986; // @[vga.scala 14:20]
  reg [7:0] ram_987; // @[vga.scala 14:20]
  reg [7:0] ram_988; // @[vga.scala 14:20]
  reg [7:0] ram_989; // @[vga.scala 14:20]
  reg [7:0] ram_990; // @[vga.scala 14:20]
  reg [7:0] ram_991; // @[vga.scala 14:20]
  reg [7:0] ram_992; // @[vga.scala 14:20]
  reg [7:0] ram_993; // @[vga.scala 14:20]
  reg [7:0] ram_994; // @[vga.scala 14:20]
  reg [7:0] ram_995; // @[vga.scala 14:20]
  reg [7:0] ram_996; // @[vga.scala 14:20]
  reg [7:0] ram_997; // @[vga.scala 14:20]
  reg [7:0] ram_998; // @[vga.scala 14:20]
  reg [7:0] ram_999; // @[vga.scala 14:20]
  reg [7:0] ram_1000; // @[vga.scala 14:20]
  reg [7:0] ram_1001; // @[vga.scala 14:20]
  reg [7:0] ram_1002; // @[vga.scala 14:20]
  reg [7:0] ram_1003; // @[vga.scala 14:20]
  reg [7:0] ram_1004; // @[vga.scala 14:20]
  reg [7:0] ram_1005; // @[vga.scala 14:20]
  reg [7:0] ram_1006; // @[vga.scala 14:20]
  reg [7:0] ram_1007; // @[vga.scala 14:20]
  reg [7:0] ram_1008; // @[vga.scala 14:20]
  reg [7:0] ram_1009; // @[vga.scala 14:20]
  reg [7:0] ram_1010; // @[vga.scala 14:20]
  reg [7:0] ram_1011; // @[vga.scala 14:20]
  reg [7:0] ram_1012; // @[vga.scala 14:20]
  reg [7:0] ram_1013; // @[vga.scala 14:20]
  reg [7:0] ram_1014; // @[vga.scala 14:20]
  reg [7:0] ram_1015; // @[vga.scala 14:20]
  reg [7:0] ram_1016; // @[vga.scala 14:20]
  reg [7:0] ram_1017; // @[vga.scala 14:20]
  reg [7:0] ram_1018; // @[vga.scala 14:20]
  reg [7:0] ram_1019; // @[vga.scala 14:20]
  reg [7:0] ram_1020; // @[vga.scala 14:20]
  reg [7:0] ram_1021; // @[vga.scala 14:20]
  reg [7:0] ram_1022; // @[vga.scala 14:20]
  reg [7:0] ram_1023; // @[vga.scala 14:20]
  reg [7:0] ram_1024; // @[vga.scala 14:20]
  reg [7:0] ram_1025; // @[vga.scala 14:20]
  reg [7:0] ram_1026; // @[vga.scala 14:20]
  reg [7:0] ram_1027; // @[vga.scala 14:20]
  reg [7:0] ram_1028; // @[vga.scala 14:20]
  reg [7:0] ram_1029; // @[vga.scala 14:20]
  reg [7:0] ram_1030; // @[vga.scala 14:20]
  reg [7:0] ram_1031; // @[vga.scala 14:20]
  reg [7:0] ram_1032; // @[vga.scala 14:20]
  reg [7:0] ram_1033; // @[vga.scala 14:20]
  reg [7:0] ram_1034; // @[vga.scala 14:20]
  reg [7:0] ram_1035; // @[vga.scala 14:20]
  reg [7:0] ram_1036; // @[vga.scala 14:20]
  reg [7:0] ram_1037; // @[vga.scala 14:20]
  reg [7:0] ram_1038; // @[vga.scala 14:20]
  reg [7:0] ram_1039; // @[vga.scala 14:20]
  reg [7:0] ram_1040; // @[vga.scala 14:20]
  reg [7:0] ram_1041; // @[vga.scala 14:20]
  reg [7:0] ram_1042; // @[vga.scala 14:20]
  reg [7:0] ram_1043; // @[vga.scala 14:20]
  reg [7:0] ram_1044; // @[vga.scala 14:20]
  reg [7:0] ram_1045; // @[vga.scala 14:20]
  reg [7:0] ram_1046; // @[vga.scala 14:20]
  reg [7:0] ram_1047; // @[vga.scala 14:20]
  reg [7:0] ram_1048; // @[vga.scala 14:20]
  reg [7:0] ram_1049; // @[vga.scala 14:20]
  reg [7:0] ram_1050; // @[vga.scala 14:20]
  reg [7:0] ram_1051; // @[vga.scala 14:20]
  reg [7:0] ram_1052; // @[vga.scala 14:20]
  reg [7:0] ram_1053; // @[vga.scala 14:20]
  reg [7:0] ram_1054; // @[vga.scala 14:20]
  reg [7:0] ram_1055; // @[vga.scala 14:20]
  reg [7:0] ram_1056; // @[vga.scala 14:20]
  reg [7:0] ram_1057; // @[vga.scala 14:20]
  reg [7:0] ram_1058; // @[vga.scala 14:20]
  reg [7:0] ram_1059; // @[vga.scala 14:20]
  reg [7:0] ram_1060; // @[vga.scala 14:20]
  reg [7:0] ram_1061; // @[vga.scala 14:20]
  reg [7:0] ram_1062; // @[vga.scala 14:20]
  reg [7:0] ram_1063; // @[vga.scala 14:20]
  reg [7:0] ram_1064; // @[vga.scala 14:20]
  reg [7:0] ram_1065; // @[vga.scala 14:20]
  reg [7:0] ram_1066; // @[vga.scala 14:20]
  reg [7:0] ram_1067; // @[vga.scala 14:20]
  reg [7:0] ram_1068; // @[vga.scala 14:20]
  reg [7:0] ram_1069; // @[vga.scala 14:20]
  reg [7:0] ram_1070; // @[vga.scala 14:20]
  reg [7:0] ram_1071; // @[vga.scala 14:20]
  reg [7:0] ram_1072; // @[vga.scala 14:20]
  reg [7:0] ram_1073; // @[vga.scala 14:20]
  reg [7:0] ram_1074; // @[vga.scala 14:20]
  reg [7:0] ram_1075; // @[vga.scala 14:20]
  reg [7:0] ram_1076; // @[vga.scala 14:20]
  reg [7:0] ram_1077; // @[vga.scala 14:20]
  reg [7:0] ram_1078; // @[vga.scala 14:20]
  reg [7:0] ram_1079; // @[vga.scala 14:20]
  reg [7:0] ram_1080; // @[vga.scala 14:20]
  reg [7:0] ram_1081; // @[vga.scala 14:20]
  reg [7:0] ram_1082; // @[vga.scala 14:20]
  reg [7:0] ram_1083; // @[vga.scala 14:20]
  reg [7:0] ram_1084; // @[vga.scala 14:20]
  reg [7:0] ram_1085; // @[vga.scala 14:20]
  reg [7:0] ram_1086; // @[vga.scala 14:20]
  reg [7:0] ram_1087; // @[vga.scala 14:20]
  reg [7:0] ram_1088; // @[vga.scala 14:20]
  reg [7:0] ram_1089; // @[vga.scala 14:20]
  reg [7:0] ram_1090; // @[vga.scala 14:20]
  reg [7:0] ram_1091; // @[vga.scala 14:20]
  reg [7:0] ram_1092; // @[vga.scala 14:20]
  reg [7:0] ram_1093; // @[vga.scala 14:20]
  reg [7:0] ram_1094; // @[vga.scala 14:20]
  reg [7:0] ram_1095; // @[vga.scala 14:20]
  reg [7:0] ram_1096; // @[vga.scala 14:20]
  reg [7:0] ram_1097; // @[vga.scala 14:20]
  reg [7:0] ram_1098; // @[vga.scala 14:20]
  reg [7:0] ram_1099; // @[vga.scala 14:20]
  reg [7:0] ram_1100; // @[vga.scala 14:20]
  reg [7:0] ram_1101; // @[vga.scala 14:20]
  reg [7:0] ram_1102; // @[vga.scala 14:20]
  reg [7:0] ram_1103; // @[vga.scala 14:20]
  reg [7:0] ram_1104; // @[vga.scala 14:20]
  reg [7:0] ram_1105; // @[vga.scala 14:20]
  reg [7:0] ram_1106; // @[vga.scala 14:20]
  reg [7:0] ram_1107; // @[vga.scala 14:20]
  reg [7:0] ram_1108; // @[vga.scala 14:20]
  reg [7:0] ram_1109; // @[vga.scala 14:20]
  reg [7:0] ram_1110; // @[vga.scala 14:20]
  reg [7:0] ram_1111; // @[vga.scala 14:20]
  reg [7:0] ram_1112; // @[vga.scala 14:20]
  reg [7:0] ram_1113; // @[vga.scala 14:20]
  reg [7:0] ram_1114; // @[vga.scala 14:20]
  reg [7:0] ram_1115; // @[vga.scala 14:20]
  reg [7:0] ram_1116; // @[vga.scala 14:20]
  reg [7:0] ram_1117; // @[vga.scala 14:20]
  reg [7:0] ram_1118; // @[vga.scala 14:20]
  reg [7:0] ram_1119; // @[vga.scala 14:20]
  reg [7:0] ram_1120; // @[vga.scala 14:20]
  reg [7:0] ram_1121; // @[vga.scala 14:20]
  reg [7:0] ram_1122; // @[vga.scala 14:20]
  reg [7:0] ram_1123; // @[vga.scala 14:20]
  reg [7:0] ram_1124; // @[vga.scala 14:20]
  reg [7:0] ram_1125; // @[vga.scala 14:20]
  reg [7:0] ram_1126; // @[vga.scala 14:20]
  reg [7:0] ram_1127; // @[vga.scala 14:20]
  reg [7:0] ram_1128; // @[vga.scala 14:20]
  reg [7:0] ram_1129; // @[vga.scala 14:20]
  reg [7:0] ram_1130; // @[vga.scala 14:20]
  reg [7:0] ram_1131; // @[vga.scala 14:20]
  reg [7:0] ram_1132; // @[vga.scala 14:20]
  reg [7:0] ram_1133; // @[vga.scala 14:20]
  reg [7:0] ram_1134; // @[vga.scala 14:20]
  reg [7:0] ram_1135; // @[vga.scala 14:20]
  reg [7:0] ram_1136; // @[vga.scala 14:20]
  reg [7:0] ram_1137; // @[vga.scala 14:20]
  reg [7:0] ram_1138; // @[vga.scala 14:20]
  reg [7:0] ram_1139; // @[vga.scala 14:20]
  reg [7:0] ram_1140; // @[vga.scala 14:20]
  reg [7:0] ram_1141; // @[vga.scala 14:20]
  reg [7:0] ram_1142; // @[vga.scala 14:20]
  reg [7:0] ram_1143; // @[vga.scala 14:20]
  reg [7:0] ram_1144; // @[vga.scala 14:20]
  reg [7:0] ram_1145; // @[vga.scala 14:20]
  reg [7:0] ram_1146; // @[vga.scala 14:20]
  reg [7:0] ram_1147; // @[vga.scala 14:20]
  reg [7:0] ram_1148; // @[vga.scala 14:20]
  reg [7:0] ram_1149; // @[vga.scala 14:20]
  reg [7:0] ram_1150; // @[vga.scala 14:20]
  reg [7:0] ram_1151; // @[vga.scala 14:20]
  reg [7:0] ram_1152; // @[vga.scala 14:20]
  reg [7:0] ram_1153; // @[vga.scala 14:20]
  reg [7:0] ram_1154; // @[vga.scala 14:20]
  reg [7:0] ram_1155; // @[vga.scala 14:20]
  reg [7:0] ram_1156; // @[vga.scala 14:20]
  reg [7:0] ram_1157; // @[vga.scala 14:20]
  reg [7:0] ram_1158; // @[vga.scala 14:20]
  reg [7:0] ram_1159; // @[vga.scala 14:20]
  reg [7:0] ram_1160; // @[vga.scala 14:20]
  reg [7:0] ram_1161; // @[vga.scala 14:20]
  reg [7:0] ram_1162; // @[vga.scala 14:20]
  reg [7:0] ram_1163; // @[vga.scala 14:20]
  reg [7:0] ram_1164; // @[vga.scala 14:20]
  reg [7:0] ram_1165; // @[vga.scala 14:20]
  reg [7:0] ram_1166; // @[vga.scala 14:20]
  reg [7:0] ram_1167; // @[vga.scala 14:20]
  reg [7:0] ram_1168; // @[vga.scala 14:20]
  reg [7:0] ram_1169; // @[vga.scala 14:20]
  reg [7:0] ram_1170; // @[vga.scala 14:20]
  reg [7:0] ram_1171; // @[vga.scala 14:20]
  reg [7:0] ram_1172; // @[vga.scala 14:20]
  reg [7:0] ram_1173; // @[vga.scala 14:20]
  reg [7:0] ram_1174; // @[vga.scala 14:20]
  reg [7:0] ram_1175; // @[vga.scala 14:20]
  reg [7:0] ram_1176; // @[vga.scala 14:20]
  reg [7:0] ram_1177; // @[vga.scala 14:20]
  reg [7:0] ram_1178; // @[vga.scala 14:20]
  reg [7:0] ram_1179; // @[vga.scala 14:20]
  reg [7:0] ram_1180; // @[vga.scala 14:20]
  reg [7:0] ram_1181; // @[vga.scala 14:20]
  reg [7:0] ram_1182; // @[vga.scala 14:20]
  reg [7:0] ram_1183; // @[vga.scala 14:20]
  reg [7:0] ram_1184; // @[vga.scala 14:20]
  reg [7:0] ram_1185; // @[vga.scala 14:20]
  reg [7:0] ram_1186; // @[vga.scala 14:20]
  reg [7:0] ram_1187; // @[vga.scala 14:20]
  reg [7:0] ram_1188; // @[vga.scala 14:20]
  reg [7:0] ram_1189; // @[vga.scala 14:20]
  reg [7:0] ram_1190; // @[vga.scala 14:20]
  reg [7:0] ram_1191; // @[vga.scala 14:20]
  reg [7:0] ram_1192; // @[vga.scala 14:20]
  reg [7:0] ram_1193; // @[vga.scala 14:20]
  reg [7:0] ram_1194; // @[vga.scala 14:20]
  reg [7:0] ram_1195; // @[vga.scala 14:20]
  reg [7:0] ram_1196; // @[vga.scala 14:20]
  reg [7:0] ram_1197; // @[vga.scala 14:20]
  reg [7:0] ram_1198; // @[vga.scala 14:20]
  reg [7:0] ram_1199; // @[vga.scala 14:20]
  reg [7:0] ram_1200; // @[vga.scala 14:20]
  reg [7:0] ram_1201; // @[vga.scala 14:20]
  reg [7:0] ram_1202; // @[vga.scala 14:20]
  reg [7:0] ram_1203; // @[vga.scala 14:20]
  reg [7:0] ram_1204; // @[vga.scala 14:20]
  reg [7:0] ram_1205; // @[vga.scala 14:20]
  reg [7:0] ram_1206; // @[vga.scala 14:20]
  reg [7:0] ram_1207; // @[vga.scala 14:20]
  reg [7:0] ram_1208; // @[vga.scala 14:20]
  reg [7:0] ram_1209; // @[vga.scala 14:20]
  reg [7:0] ram_1210; // @[vga.scala 14:20]
  reg [7:0] ram_1211; // @[vga.scala 14:20]
  reg [7:0] ram_1212; // @[vga.scala 14:20]
  reg [7:0] ram_1213; // @[vga.scala 14:20]
  reg [7:0] ram_1214; // @[vga.scala 14:20]
  reg [7:0] ram_1215; // @[vga.scala 14:20]
  reg [7:0] ram_1216; // @[vga.scala 14:20]
  reg [7:0] ram_1217; // @[vga.scala 14:20]
  reg [7:0] ram_1218; // @[vga.scala 14:20]
  reg [7:0] ram_1219; // @[vga.scala 14:20]
  reg [7:0] ram_1220; // @[vga.scala 14:20]
  reg [7:0] ram_1221; // @[vga.scala 14:20]
  reg [7:0] ram_1222; // @[vga.scala 14:20]
  reg [7:0] ram_1223; // @[vga.scala 14:20]
  reg [7:0] ram_1224; // @[vga.scala 14:20]
  reg [7:0] ram_1225; // @[vga.scala 14:20]
  reg [7:0] ram_1226; // @[vga.scala 14:20]
  reg [7:0] ram_1227; // @[vga.scala 14:20]
  reg [7:0] ram_1228; // @[vga.scala 14:20]
  reg [7:0] ram_1229; // @[vga.scala 14:20]
  reg [7:0] ram_1230; // @[vga.scala 14:20]
  reg [7:0] ram_1231; // @[vga.scala 14:20]
  reg [7:0] ram_1232; // @[vga.scala 14:20]
  reg [7:0] ram_1233; // @[vga.scala 14:20]
  reg [7:0] ram_1234; // @[vga.scala 14:20]
  reg [7:0] ram_1235; // @[vga.scala 14:20]
  reg [7:0] ram_1236; // @[vga.scala 14:20]
  reg [7:0] ram_1237; // @[vga.scala 14:20]
  reg [7:0] ram_1238; // @[vga.scala 14:20]
  reg [7:0] ram_1239; // @[vga.scala 14:20]
  reg [7:0] ram_1240; // @[vga.scala 14:20]
  reg [7:0] ram_1241; // @[vga.scala 14:20]
  reg [7:0] ram_1242; // @[vga.scala 14:20]
  reg [7:0] ram_1243; // @[vga.scala 14:20]
  reg [7:0] ram_1244; // @[vga.scala 14:20]
  reg [7:0] ram_1245; // @[vga.scala 14:20]
  reg [7:0] ram_1246; // @[vga.scala 14:20]
  reg [7:0] ram_1247; // @[vga.scala 14:20]
  reg [7:0] ram_1248; // @[vga.scala 14:20]
  reg [7:0] ram_1249; // @[vga.scala 14:20]
  reg [7:0] ram_1250; // @[vga.scala 14:20]
  reg [7:0] ram_1251; // @[vga.scala 14:20]
  reg [7:0] ram_1252; // @[vga.scala 14:20]
  reg [7:0] ram_1253; // @[vga.scala 14:20]
  reg [7:0] ram_1254; // @[vga.scala 14:20]
  reg [7:0] ram_1255; // @[vga.scala 14:20]
  reg [7:0] ram_1256; // @[vga.scala 14:20]
  reg [7:0] ram_1257; // @[vga.scala 14:20]
  reg [7:0] ram_1258; // @[vga.scala 14:20]
  reg [7:0] ram_1259; // @[vga.scala 14:20]
  reg [7:0] ram_1260; // @[vga.scala 14:20]
  reg [7:0] ram_1261; // @[vga.scala 14:20]
  reg [7:0] ram_1262; // @[vga.scala 14:20]
  reg [7:0] ram_1263; // @[vga.scala 14:20]
  reg [7:0] ram_1264; // @[vga.scala 14:20]
  reg [7:0] ram_1265; // @[vga.scala 14:20]
  reg [7:0] ram_1266; // @[vga.scala 14:20]
  reg [7:0] ram_1267; // @[vga.scala 14:20]
  reg [7:0] ram_1268; // @[vga.scala 14:20]
  reg [7:0] ram_1269; // @[vga.scala 14:20]
  reg [7:0] ram_1270; // @[vga.scala 14:20]
  reg [7:0] ram_1271; // @[vga.scala 14:20]
  reg [7:0] ram_1272; // @[vga.scala 14:20]
  reg [7:0] ram_1273; // @[vga.scala 14:20]
  reg [7:0] ram_1274; // @[vga.scala 14:20]
  reg [7:0] ram_1275; // @[vga.scala 14:20]
  reg [7:0] ram_1276; // @[vga.scala 14:20]
  reg [7:0] ram_1277; // @[vga.scala 14:20]
  reg [7:0] ram_1278; // @[vga.scala 14:20]
  reg [7:0] ram_1279; // @[vga.scala 14:20]
  reg [7:0] ram_1280; // @[vga.scala 14:20]
  reg [7:0] ram_1281; // @[vga.scala 14:20]
  reg [7:0] ram_1282; // @[vga.scala 14:20]
  reg [7:0] ram_1283; // @[vga.scala 14:20]
  reg [7:0] ram_1284; // @[vga.scala 14:20]
  reg [7:0] ram_1285; // @[vga.scala 14:20]
  reg [7:0] ram_1286; // @[vga.scala 14:20]
  reg [7:0] ram_1287; // @[vga.scala 14:20]
  reg [7:0] ram_1288; // @[vga.scala 14:20]
  reg [7:0] ram_1289; // @[vga.scala 14:20]
  reg [7:0] ram_1290; // @[vga.scala 14:20]
  reg [7:0] ram_1291; // @[vga.scala 14:20]
  reg [7:0] ram_1292; // @[vga.scala 14:20]
  reg [7:0] ram_1293; // @[vga.scala 14:20]
  reg [7:0] ram_1294; // @[vga.scala 14:20]
  reg [7:0] ram_1295; // @[vga.scala 14:20]
  reg [7:0] ram_1296; // @[vga.scala 14:20]
  reg [7:0] ram_1297; // @[vga.scala 14:20]
  reg [7:0] ram_1298; // @[vga.scala 14:20]
  reg [7:0] ram_1299; // @[vga.scala 14:20]
  reg [7:0] ram_1300; // @[vga.scala 14:20]
  reg [7:0] ram_1301; // @[vga.scala 14:20]
  reg [7:0] ram_1302; // @[vga.scala 14:20]
  reg [7:0] ram_1303; // @[vga.scala 14:20]
  reg [7:0] ram_1304; // @[vga.scala 14:20]
  reg [7:0] ram_1305; // @[vga.scala 14:20]
  reg [7:0] ram_1306; // @[vga.scala 14:20]
  reg [7:0] ram_1307; // @[vga.scala 14:20]
  reg [7:0] ram_1308; // @[vga.scala 14:20]
  reg [7:0] ram_1309; // @[vga.scala 14:20]
  reg [7:0] ram_1310; // @[vga.scala 14:20]
  reg [7:0] ram_1311; // @[vga.scala 14:20]
  reg [7:0] ram_1312; // @[vga.scala 14:20]
  reg [7:0] ram_1313; // @[vga.scala 14:20]
  reg [7:0] ram_1314; // @[vga.scala 14:20]
  reg [7:0] ram_1315; // @[vga.scala 14:20]
  reg [7:0] ram_1316; // @[vga.scala 14:20]
  reg [7:0] ram_1317; // @[vga.scala 14:20]
  reg [7:0] ram_1318; // @[vga.scala 14:20]
  reg [7:0] ram_1319; // @[vga.scala 14:20]
  reg [7:0] ram_1320; // @[vga.scala 14:20]
  reg [7:0] ram_1321; // @[vga.scala 14:20]
  reg [7:0] ram_1322; // @[vga.scala 14:20]
  reg [7:0] ram_1323; // @[vga.scala 14:20]
  reg [7:0] ram_1324; // @[vga.scala 14:20]
  reg [7:0] ram_1325; // @[vga.scala 14:20]
  reg [7:0] ram_1326; // @[vga.scala 14:20]
  reg [7:0] ram_1327; // @[vga.scala 14:20]
  reg [7:0] ram_1328; // @[vga.scala 14:20]
  reg [7:0] ram_1329; // @[vga.scala 14:20]
  reg [7:0] ram_1330; // @[vga.scala 14:20]
  reg [7:0] ram_1331; // @[vga.scala 14:20]
  reg [7:0] ram_1332; // @[vga.scala 14:20]
  reg [7:0] ram_1333; // @[vga.scala 14:20]
  reg [7:0] ram_1334; // @[vga.scala 14:20]
  reg [7:0] ram_1335; // @[vga.scala 14:20]
  reg [7:0] ram_1336; // @[vga.scala 14:20]
  reg [7:0] ram_1337; // @[vga.scala 14:20]
  reg [7:0] ram_1338; // @[vga.scala 14:20]
  reg [7:0] ram_1339; // @[vga.scala 14:20]
  reg [7:0] ram_1340; // @[vga.scala 14:20]
  reg [7:0] ram_1341; // @[vga.scala 14:20]
  reg [7:0] ram_1342; // @[vga.scala 14:20]
  reg [7:0] ram_1343; // @[vga.scala 14:20]
  reg [7:0] ram_1344; // @[vga.scala 14:20]
  reg [7:0] ram_1345; // @[vga.scala 14:20]
  reg [7:0] ram_1346; // @[vga.scala 14:20]
  reg [7:0] ram_1347; // @[vga.scala 14:20]
  reg [7:0] ram_1348; // @[vga.scala 14:20]
  reg [7:0] ram_1349; // @[vga.scala 14:20]
  reg [7:0] ram_1350; // @[vga.scala 14:20]
  reg [7:0] ram_1351; // @[vga.scala 14:20]
  reg [7:0] ram_1352; // @[vga.scala 14:20]
  reg [7:0] ram_1353; // @[vga.scala 14:20]
  reg [7:0] ram_1354; // @[vga.scala 14:20]
  reg [7:0] ram_1355; // @[vga.scala 14:20]
  reg [7:0] ram_1356; // @[vga.scala 14:20]
  reg [7:0] ram_1357; // @[vga.scala 14:20]
  reg [7:0] ram_1358; // @[vga.scala 14:20]
  reg [7:0] ram_1359; // @[vga.scala 14:20]
  reg [7:0] ram_1360; // @[vga.scala 14:20]
  reg [7:0] ram_1361; // @[vga.scala 14:20]
  reg [7:0] ram_1362; // @[vga.scala 14:20]
  reg [7:0] ram_1363; // @[vga.scala 14:20]
  reg [7:0] ram_1364; // @[vga.scala 14:20]
  reg [7:0] ram_1365; // @[vga.scala 14:20]
  reg [7:0] ram_1366; // @[vga.scala 14:20]
  reg [7:0] ram_1367; // @[vga.scala 14:20]
  reg [7:0] ram_1368; // @[vga.scala 14:20]
  reg [7:0] ram_1369; // @[vga.scala 14:20]
  reg [7:0] ram_1370; // @[vga.scala 14:20]
  reg [7:0] ram_1371; // @[vga.scala 14:20]
  reg [7:0] ram_1372; // @[vga.scala 14:20]
  reg [7:0] ram_1373; // @[vga.scala 14:20]
  reg [7:0] ram_1374; // @[vga.scala 14:20]
  reg [7:0] ram_1375; // @[vga.scala 14:20]
  reg [7:0] ram_1376; // @[vga.scala 14:20]
  reg [7:0] ram_1377; // @[vga.scala 14:20]
  reg [7:0] ram_1378; // @[vga.scala 14:20]
  reg [7:0] ram_1379; // @[vga.scala 14:20]
  reg [7:0] ram_1380; // @[vga.scala 14:20]
  reg [7:0] ram_1381; // @[vga.scala 14:20]
  reg [7:0] ram_1382; // @[vga.scala 14:20]
  reg [7:0] ram_1383; // @[vga.scala 14:20]
  reg [7:0] ram_1384; // @[vga.scala 14:20]
  reg [7:0] ram_1385; // @[vga.scala 14:20]
  reg [7:0] ram_1386; // @[vga.scala 14:20]
  reg [7:0] ram_1387; // @[vga.scala 14:20]
  reg [7:0] ram_1388; // @[vga.scala 14:20]
  reg [7:0] ram_1389; // @[vga.scala 14:20]
  reg [7:0] ram_1390; // @[vga.scala 14:20]
  reg [7:0] ram_1391; // @[vga.scala 14:20]
  reg [7:0] ram_1392; // @[vga.scala 14:20]
  reg [7:0] ram_1393; // @[vga.scala 14:20]
  reg [7:0] ram_1394; // @[vga.scala 14:20]
  reg [7:0] ram_1395; // @[vga.scala 14:20]
  reg [7:0] ram_1396; // @[vga.scala 14:20]
  reg [7:0] ram_1397; // @[vga.scala 14:20]
  reg [7:0] ram_1398; // @[vga.scala 14:20]
  reg [7:0] ram_1399; // @[vga.scala 14:20]
  reg [7:0] ram_1400; // @[vga.scala 14:20]
  reg [7:0] ram_1401; // @[vga.scala 14:20]
  reg [7:0] ram_1402; // @[vga.scala 14:20]
  reg [7:0] ram_1403; // @[vga.scala 14:20]
  reg [7:0] ram_1404; // @[vga.scala 14:20]
  reg [7:0] ram_1405; // @[vga.scala 14:20]
  reg [7:0] ram_1406; // @[vga.scala 14:20]
  reg [7:0] ram_1407; // @[vga.scala 14:20]
  reg [7:0] ram_1408; // @[vga.scala 14:20]
  reg [7:0] ram_1409; // @[vga.scala 14:20]
  reg [7:0] ram_1410; // @[vga.scala 14:20]
  reg [7:0] ram_1411; // @[vga.scala 14:20]
  reg [7:0] ram_1412; // @[vga.scala 14:20]
  reg [7:0] ram_1413; // @[vga.scala 14:20]
  reg [7:0] ram_1414; // @[vga.scala 14:20]
  reg [7:0] ram_1415; // @[vga.scala 14:20]
  reg [7:0] ram_1416; // @[vga.scala 14:20]
  reg [7:0] ram_1417; // @[vga.scala 14:20]
  reg [7:0] ram_1418; // @[vga.scala 14:20]
  reg [7:0] ram_1419; // @[vga.scala 14:20]
  reg [7:0] ram_1420; // @[vga.scala 14:20]
  reg [7:0] ram_1421; // @[vga.scala 14:20]
  reg [7:0] ram_1422; // @[vga.scala 14:20]
  reg [7:0] ram_1423; // @[vga.scala 14:20]
  reg [7:0] ram_1424; // @[vga.scala 14:20]
  reg [7:0] ram_1425; // @[vga.scala 14:20]
  reg [7:0] ram_1426; // @[vga.scala 14:20]
  reg [7:0] ram_1427; // @[vga.scala 14:20]
  reg [7:0] ram_1428; // @[vga.scala 14:20]
  reg [7:0] ram_1429; // @[vga.scala 14:20]
  reg [7:0] ram_1430; // @[vga.scala 14:20]
  reg [7:0] ram_1431; // @[vga.scala 14:20]
  reg [7:0] ram_1432; // @[vga.scala 14:20]
  reg [7:0] ram_1433; // @[vga.scala 14:20]
  reg [7:0] ram_1434; // @[vga.scala 14:20]
  reg [7:0] ram_1435; // @[vga.scala 14:20]
  reg [7:0] ram_1436; // @[vga.scala 14:20]
  reg [7:0] ram_1437; // @[vga.scala 14:20]
  reg [7:0] ram_1438; // @[vga.scala 14:20]
  reg [7:0] ram_1439; // @[vga.scala 14:20]
  reg [7:0] ram_1440; // @[vga.scala 14:20]
  reg [7:0] ram_1441; // @[vga.scala 14:20]
  reg [7:0] ram_1442; // @[vga.scala 14:20]
  reg [7:0] ram_1443; // @[vga.scala 14:20]
  reg [7:0] ram_1444; // @[vga.scala 14:20]
  reg [7:0] ram_1445; // @[vga.scala 14:20]
  reg [7:0] ram_1446; // @[vga.scala 14:20]
  reg [7:0] ram_1447; // @[vga.scala 14:20]
  reg [7:0] ram_1448; // @[vga.scala 14:20]
  reg [7:0] ram_1449; // @[vga.scala 14:20]
  reg [7:0] ram_1450; // @[vga.scala 14:20]
  reg [7:0] ram_1451; // @[vga.scala 14:20]
  reg [7:0] ram_1452; // @[vga.scala 14:20]
  reg [7:0] ram_1453; // @[vga.scala 14:20]
  reg [7:0] ram_1454; // @[vga.scala 14:20]
  reg [7:0] ram_1455; // @[vga.scala 14:20]
  reg [7:0] ram_1456; // @[vga.scala 14:20]
  reg [7:0] ram_1457; // @[vga.scala 14:20]
  reg [7:0] ram_1458; // @[vga.scala 14:20]
  reg [7:0] ram_1459; // @[vga.scala 14:20]
  reg [7:0] ram_1460; // @[vga.scala 14:20]
  reg [7:0] ram_1461; // @[vga.scala 14:20]
  reg [7:0] ram_1462; // @[vga.scala 14:20]
  reg [7:0] ram_1463; // @[vga.scala 14:20]
  reg [7:0] ram_1464; // @[vga.scala 14:20]
  reg [7:0] ram_1465; // @[vga.scala 14:20]
  reg [7:0] ram_1466; // @[vga.scala 14:20]
  reg [7:0] ram_1467; // @[vga.scala 14:20]
  reg [7:0] ram_1468; // @[vga.scala 14:20]
  reg [7:0] ram_1469; // @[vga.scala 14:20]
  reg [7:0] ram_1470; // @[vga.scala 14:20]
  reg [7:0] ram_1471; // @[vga.scala 14:20]
  reg [7:0] ram_1472; // @[vga.scala 14:20]
  reg [7:0] ram_1473; // @[vga.scala 14:20]
  reg [7:0] ram_1474; // @[vga.scala 14:20]
  reg [7:0] ram_1475; // @[vga.scala 14:20]
  reg [7:0] ram_1476; // @[vga.scala 14:20]
  reg [7:0] ram_1477; // @[vga.scala 14:20]
  reg [7:0] ram_1478; // @[vga.scala 14:20]
  reg [7:0] ram_1479; // @[vga.scala 14:20]
  reg [7:0] ram_1480; // @[vga.scala 14:20]
  reg [7:0] ram_1481; // @[vga.scala 14:20]
  reg [7:0] ram_1482; // @[vga.scala 14:20]
  reg [7:0] ram_1483; // @[vga.scala 14:20]
  reg [7:0] ram_1484; // @[vga.scala 14:20]
  reg [7:0] ram_1485; // @[vga.scala 14:20]
  reg [7:0] ram_1486; // @[vga.scala 14:20]
  reg [7:0] ram_1487; // @[vga.scala 14:20]
  reg [7:0] ram_1488; // @[vga.scala 14:20]
  reg [7:0] ram_1489; // @[vga.scala 14:20]
  reg [7:0] ram_1490; // @[vga.scala 14:20]
  reg [7:0] ram_1491; // @[vga.scala 14:20]
  reg [7:0] ram_1492; // @[vga.scala 14:20]
  reg [7:0] ram_1493; // @[vga.scala 14:20]
  reg [7:0] ram_1494; // @[vga.scala 14:20]
  reg [7:0] ram_1495; // @[vga.scala 14:20]
  reg [7:0] ram_1496; // @[vga.scala 14:20]
  reg [7:0] ram_1497; // @[vga.scala 14:20]
  reg [7:0] ram_1498; // @[vga.scala 14:20]
  reg [7:0] ram_1499; // @[vga.scala 14:20]
  reg [7:0] ram_1500; // @[vga.scala 14:20]
  reg [7:0] ram_1501; // @[vga.scala 14:20]
  reg [7:0] ram_1502; // @[vga.scala 14:20]
  reg [7:0] ram_1503; // @[vga.scala 14:20]
  reg [7:0] ram_1504; // @[vga.scala 14:20]
  reg [7:0] ram_1505; // @[vga.scala 14:20]
  reg [7:0] ram_1506; // @[vga.scala 14:20]
  reg [7:0] ram_1507; // @[vga.scala 14:20]
  reg [7:0] ram_1508; // @[vga.scala 14:20]
  reg [7:0] ram_1509; // @[vga.scala 14:20]
  reg [7:0] ram_1510; // @[vga.scala 14:20]
  reg [7:0] ram_1511; // @[vga.scala 14:20]
  reg [7:0] ram_1512; // @[vga.scala 14:20]
  reg [7:0] ram_1513; // @[vga.scala 14:20]
  reg [7:0] ram_1514; // @[vga.scala 14:20]
  reg [7:0] ram_1515; // @[vga.scala 14:20]
  reg [7:0] ram_1516; // @[vga.scala 14:20]
  reg [7:0] ram_1517; // @[vga.scala 14:20]
  reg [7:0] ram_1518; // @[vga.scala 14:20]
  reg [7:0] ram_1519; // @[vga.scala 14:20]
  reg [7:0] ram_1520; // @[vga.scala 14:20]
  reg [7:0] ram_1521; // @[vga.scala 14:20]
  reg [7:0] ram_1522; // @[vga.scala 14:20]
  reg [7:0] ram_1523; // @[vga.scala 14:20]
  reg [7:0] ram_1524; // @[vga.scala 14:20]
  reg [7:0] ram_1525; // @[vga.scala 14:20]
  reg [7:0] ram_1526; // @[vga.scala 14:20]
  reg [7:0] ram_1527; // @[vga.scala 14:20]
  reg [7:0] ram_1528; // @[vga.scala 14:20]
  reg [7:0] ram_1529; // @[vga.scala 14:20]
  reg [7:0] ram_1530; // @[vga.scala 14:20]
  reg [7:0] ram_1531; // @[vga.scala 14:20]
  reg [7:0] ram_1532; // @[vga.scala 14:20]
  reg [7:0] ram_1533; // @[vga.scala 14:20]
  reg [7:0] ram_1534; // @[vga.scala 14:20]
  reg [7:0] ram_1535; // @[vga.scala 14:20]
  reg [7:0] ram_1536; // @[vga.scala 14:20]
  reg [7:0] ram_1537; // @[vga.scala 14:20]
  reg [7:0] ram_1538; // @[vga.scala 14:20]
  reg [7:0] ram_1539; // @[vga.scala 14:20]
  reg [7:0] ram_1540; // @[vga.scala 14:20]
  reg [7:0] ram_1541; // @[vga.scala 14:20]
  reg [7:0] ram_1542; // @[vga.scala 14:20]
  reg [7:0] ram_1543; // @[vga.scala 14:20]
  reg [7:0] ram_1544; // @[vga.scala 14:20]
  reg [7:0] ram_1545; // @[vga.scala 14:20]
  reg [7:0] ram_1546; // @[vga.scala 14:20]
  reg [7:0] ram_1547; // @[vga.scala 14:20]
  reg [7:0] ram_1548; // @[vga.scala 14:20]
  reg [7:0] ram_1549; // @[vga.scala 14:20]
  reg [7:0] ram_1550; // @[vga.scala 14:20]
  reg [7:0] ram_1551; // @[vga.scala 14:20]
  reg [7:0] ram_1552; // @[vga.scala 14:20]
  reg [7:0] ram_1553; // @[vga.scala 14:20]
  reg [7:0] ram_1554; // @[vga.scala 14:20]
  reg [7:0] ram_1555; // @[vga.scala 14:20]
  reg [7:0] ram_1556; // @[vga.scala 14:20]
  reg [7:0] ram_1557; // @[vga.scala 14:20]
  reg [7:0] ram_1558; // @[vga.scala 14:20]
  reg [7:0] ram_1559; // @[vga.scala 14:20]
  reg [7:0] ram_1560; // @[vga.scala 14:20]
  reg [7:0] ram_1561; // @[vga.scala 14:20]
  reg [7:0] ram_1562; // @[vga.scala 14:20]
  reg [7:0] ram_1563; // @[vga.scala 14:20]
  reg [7:0] ram_1564; // @[vga.scala 14:20]
  reg [7:0] ram_1565; // @[vga.scala 14:20]
  reg [7:0] ram_1566; // @[vga.scala 14:20]
  reg [7:0] ram_1567; // @[vga.scala 14:20]
  reg [7:0] ram_1568; // @[vga.scala 14:20]
  reg [7:0] ram_1569; // @[vga.scala 14:20]
  reg [7:0] ram_1570; // @[vga.scala 14:20]
  reg [7:0] ram_1571; // @[vga.scala 14:20]
  reg [7:0] ram_1572; // @[vga.scala 14:20]
  reg [7:0] ram_1573; // @[vga.scala 14:20]
  reg [7:0] ram_1574; // @[vga.scala 14:20]
  reg [7:0] ram_1575; // @[vga.scala 14:20]
  reg [7:0] ram_1576; // @[vga.scala 14:20]
  reg [7:0] ram_1577; // @[vga.scala 14:20]
  reg [7:0] ram_1578; // @[vga.scala 14:20]
  reg [7:0] ram_1579; // @[vga.scala 14:20]
  reg [7:0] ram_1580; // @[vga.scala 14:20]
  reg [7:0] ram_1581; // @[vga.scala 14:20]
  reg [7:0] ram_1582; // @[vga.scala 14:20]
  reg [7:0] ram_1583; // @[vga.scala 14:20]
  reg [7:0] ram_1584; // @[vga.scala 14:20]
  reg [7:0] ram_1585; // @[vga.scala 14:20]
  reg [7:0] ram_1586; // @[vga.scala 14:20]
  reg [7:0] ram_1587; // @[vga.scala 14:20]
  reg [7:0] ram_1588; // @[vga.scala 14:20]
  reg [7:0] ram_1589; // @[vga.scala 14:20]
  reg [7:0] ram_1590; // @[vga.scala 14:20]
  reg [7:0] ram_1591; // @[vga.scala 14:20]
  reg [7:0] ram_1592; // @[vga.scala 14:20]
  reg [7:0] ram_1593; // @[vga.scala 14:20]
  reg [7:0] ram_1594; // @[vga.scala 14:20]
  reg [7:0] ram_1595; // @[vga.scala 14:20]
  reg [7:0] ram_1596; // @[vga.scala 14:20]
  reg [7:0] ram_1597; // @[vga.scala 14:20]
  reg [7:0] ram_1598; // @[vga.scala 14:20]
  reg [7:0] ram_1599; // @[vga.scala 14:20]
  reg [7:0] ram_1600; // @[vga.scala 14:20]
  reg [7:0] ram_1601; // @[vga.scala 14:20]
  reg [7:0] ram_1602; // @[vga.scala 14:20]
  reg [7:0] ram_1603; // @[vga.scala 14:20]
  reg [7:0] ram_1604; // @[vga.scala 14:20]
  reg [7:0] ram_1605; // @[vga.scala 14:20]
  reg [7:0] ram_1606; // @[vga.scala 14:20]
  reg [7:0] ram_1607; // @[vga.scala 14:20]
  reg [7:0] ram_1608; // @[vga.scala 14:20]
  reg [7:0] ram_1609; // @[vga.scala 14:20]
  reg [7:0] ram_1610; // @[vga.scala 14:20]
  reg [7:0] ram_1611; // @[vga.scala 14:20]
  reg [7:0] ram_1612; // @[vga.scala 14:20]
  reg [7:0] ram_1613; // @[vga.scala 14:20]
  reg [7:0] ram_1614; // @[vga.scala 14:20]
  reg [7:0] ram_1615; // @[vga.scala 14:20]
  reg [7:0] ram_1616; // @[vga.scala 14:20]
  reg [7:0] ram_1617; // @[vga.scala 14:20]
  reg [7:0] ram_1618; // @[vga.scala 14:20]
  reg [7:0] ram_1619; // @[vga.scala 14:20]
  reg [7:0] ram_1620; // @[vga.scala 14:20]
  reg [7:0] ram_1621; // @[vga.scala 14:20]
  reg [7:0] ram_1622; // @[vga.scala 14:20]
  reg [7:0] ram_1623; // @[vga.scala 14:20]
  reg [7:0] ram_1624; // @[vga.scala 14:20]
  reg [7:0] ram_1625; // @[vga.scala 14:20]
  reg [7:0] ram_1626; // @[vga.scala 14:20]
  reg [7:0] ram_1627; // @[vga.scala 14:20]
  reg [7:0] ram_1628; // @[vga.scala 14:20]
  reg [7:0] ram_1629; // @[vga.scala 14:20]
  reg [7:0] ram_1630; // @[vga.scala 14:20]
  reg [7:0] ram_1631; // @[vga.scala 14:20]
  reg [7:0] ram_1632; // @[vga.scala 14:20]
  reg [7:0] ram_1633; // @[vga.scala 14:20]
  reg [7:0] ram_1634; // @[vga.scala 14:20]
  reg [7:0] ram_1635; // @[vga.scala 14:20]
  reg [7:0] ram_1636; // @[vga.scala 14:20]
  reg [7:0] ram_1637; // @[vga.scala 14:20]
  reg [7:0] ram_1638; // @[vga.scala 14:20]
  reg [7:0] ram_1639; // @[vga.scala 14:20]
  reg [7:0] ram_1640; // @[vga.scala 14:20]
  reg [7:0] ram_1641; // @[vga.scala 14:20]
  reg [7:0] ram_1642; // @[vga.scala 14:20]
  reg [7:0] ram_1643; // @[vga.scala 14:20]
  reg [7:0] ram_1644; // @[vga.scala 14:20]
  reg [7:0] ram_1645; // @[vga.scala 14:20]
  reg [7:0] ram_1646; // @[vga.scala 14:20]
  reg [7:0] ram_1647; // @[vga.scala 14:20]
  reg [7:0] ram_1648; // @[vga.scala 14:20]
  reg [7:0] ram_1649; // @[vga.scala 14:20]
  reg [7:0] ram_1650; // @[vga.scala 14:20]
  reg [7:0] ram_1651; // @[vga.scala 14:20]
  reg [7:0] ram_1652; // @[vga.scala 14:20]
  reg [7:0] ram_1653; // @[vga.scala 14:20]
  reg [7:0] ram_1654; // @[vga.scala 14:20]
  reg [7:0] ram_1655; // @[vga.scala 14:20]
  reg [7:0] ram_1656; // @[vga.scala 14:20]
  reg [7:0] ram_1657; // @[vga.scala 14:20]
  reg [7:0] ram_1658; // @[vga.scala 14:20]
  reg [7:0] ram_1659; // @[vga.scala 14:20]
  reg [7:0] ram_1660; // @[vga.scala 14:20]
  reg [7:0] ram_1661; // @[vga.scala 14:20]
  reg [7:0] ram_1662; // @[vga.scala 14:20]
  reg [7:0] ram_1663; // @[vga.scala 14:20]
  reg [7:0] ram_1664; // @[vga.scala 14:20]
  reg [7:0] ram_1665; // @[vga.scala 14:20]
  reg [7:0] ram_1666; // @[vga.scala 14:20]
  reg [7:0] ram_1667; // @[vga.scala 14:20]
  reg [7:0] ram_1668; // @[vga.scala 14:20]
  reg [7:0] ram_1669; // @[vga.scala 14:20]
  reg [7:0] ram_1670; // @[vga.scala 14:20]
  reg [7:0] ram_1671; // @[vga.scala 14:20]
  reg [7:0] ram_1672; // @[vga.scala 14:20]
  reg [7:0] ram_1673; // @[vga.scala 14:20]
  reg [7:0] ram_1674; // @[vga.scala 14:20]
  reg [7:0] ram_1675; // @[vga.scala 14:20]
  reg [7:0] ram_1676; // @[vga.scala 14:20]
  reg [7:0] ram_1677; // @[vga.scala 14:20]
  reg [7:0] ram_1678; // @[vga.scala 14:20]
  reg [7:0] ram_1679; // @[vga.scala 14:20]
  reg [7:0] ram_1680; // @[vga.scala 14:20]
  reg [7:0] ram_1681; // @[vga.scala 14:20]
  reg [7:0] ram_1682; // @[vga.scala 14:20]
  reg [7:0] ram_1683; // @[vga.scala 14:20]
  reg [7:0] ram_1684; // @[vga.scala 14:20]
  reg [7:0] ram_1685; // @[vga.scala 14:20]
  reg [7:0] ram_1686; // @[vga.scala 14:20]
  reg [7:0] ram_1687; // @[vga.scala 14:20]
  reg [7:0] ram_1688; // @[vga.scala 14:20]
  reg [7:0] ram_1689; // @[vga.scala 14:20]
  reg [7:0] ram_1690; // @[vga.scala 14:20]
  reg [7:0] ram_1691; // @[vga.scala 14:20]
  reg [7:0] ram_1692; // @[vga.scala 14:20]
  reg [7:0] ram_1693; // @[vga.scala 14:20]
  reg [7:0] ram_1694; // @[vga.scala 14:20]
  reg [7:0] ram_1695; // @[vga.scala 14:20]
  reg [7:0] ram_1696; // @[vga.scala 14:20]
  reg [7:0] ram_1697; // @[vga.scala 14:20]
  reg [7:0] ram_1698; // @[vga.scala 14:20]
  reg [7:0] ram_1699; // @[vga.scala 14:20]
  reg [7:0] ram_1700; // @[vga.scala 14:20]
  reg [7:0] ram_1701; // @[vga.scala 14:20]
  reg [7:0] ram_1702; // @[vga.scala 14:20]
  reg [7:0] ram_1703; // @[vga.scala 14:20]
  reg [7:0] ram_1704; // @[vga.scala 14:20]
  reg [7:0] ram_1705; // @[vga.scala 14:20]
  reg [7:0] ram_1706; // @[vga.scala 14:20]
  reg [7:0] ram_1707; // @[vga.scala 14:20]
  reg [7:0] ram_1708; // @[vga.scala 14:20]
  reg [7:0] ram_1709; // @[vga.scala 14:20]
  reg [7:0] ram_1710; // @[vga.scala 14:20]
  reg [7:0] ram_1711; // @[vga.scala 14:20]
  reg [7:0] ram_1712; // @[vga.scala 14:20]
  reg [7:0] ram_1713; // @[vga.scala 14:20]
  reg [7:0] ram_1714; // @[vga.scala 14:20]
  reg [7:0] ram_1715; // @[vga.scala 14:20]
  reg [7:0] ram_1716; // @[vga.scala 14:20]
  reg [7:0] ram_1717; // @[vga.scala 14:20]
  reg [7:0] ram_1718; // @[vga.scala 14:20]
  reg [7:0] ram_1719; // @[vga.scala 14:20]
  reg [7:0] ram_1720; // @[vga.scala 14:20]
  reg [7:0] ram_1721; // @[vga.scala 14:20]
  reg [7:0] ram_1722; // @[vga.scala 14:20]
  reg [7:0] ram_1723; // @[vga.scala 14:20]
  reg [7:0] ram_1724; // @[vga.scala 14:20]
  reg [7:0] ram_1725; // @[vga.scala 14:20]
  reg [7:0] ram_1726; // @[vga.scala 14:20]
  reg [7:0] ram_1727; // @[vga.scala 14:20]
  reg [7:0] ram_1728; // @[vga.scala 14:20]
  reg [7:0] ram_1729; // @[vga.scala 14:20]
  reg [7:0] ram_1730; // @[vga.scala 14:20]
  reg [7:0] ram_1731; // @[vga.scala 14:20]
  reg [7:0] ram_1732; // @[vga.scala 14:20]
  reg [7:0] ram_1733; // @[vga.scala 14:20]
  reg [7:0] ram_1734; // @[vga.scala 14:20]
  reg [7:0] ram_1735; // @[vga.scala 14:20]
  reg [7:0] ram_1736; // @[vga.scala 14:20]
  reg [7:0] ram_1737; // @[vga.scala 14:20]
  reg [7:0] ram_1738; // @[vga.scala 14:20]
  reg [7:0] ram_1739; // @[vga.scala 14:20]
  reg [7:0] ram_1740; // @[vga.scala 14:20]
  reg [7:0] ram_1741; // @[vga.scala 14:20]
  reg [7:0] ram_1742; // @[vga.scala 14:20]
  reg [7:0] ram_1743; // @[vga.scala 14:20]
  reg [7:0] ram_1744; // @[vga.scala 14:20]
  reg [7:0] ram_1745; // @[vga.scala 14:20]
  reg [7:0] ram_1746; // @[vga.scala 14:20]
  reg [7:0] ram_1747; // @[vga.scala 14:20]
  reg [7:0] ram_1748; // @[vga.scala 14:20]
  reg [7:0] ram_1749; // @[vga.scala 14:20]
  reg [7:0] ram_1750; // @[vga.scala 14:20]
  reg [7:0] ram_1751; // @[vga.scala 14:20]
  reg [7:0] ram_1752; // @[vga.scala 14:20]
  reg [7:0] ram_1753; // @[vga.scala 14:20]
  reg [7:0] ram_1754; // @[vga.scala 14:20]
  reg [7:0] ram_1755; // @[vga.scala 14:20]
  reg [7:0] ram_1756; // @[vga.scala 14:20]
  reg [7:0] ram_1757; // @[vga.scala 14:20]
  reg [7:0] ram_1758; // @[vga.scala 14:20]
  reg [7:0] ram_1759; // @[vga.scala 14:20]
  reg [7:0] ram_1760; // @[vga.scala 14:20]
  reg [7:0] ram_1761; // @[vga.scala 14:20]
  reg [7:0] ram_1762; // @[vga.scala 14:20]
  reg [7:0] ram_1763; // @[vga.scala 14:20]
  reg [7:0] ram_1764; // @[vga.scala 14:20]
  reg [7:0] ram_1765; // @[vga.scala 14:20]
  reg [7:0] ram_1766; // @[vga.scala 14:20]
  reg [7:0] ram_1767; // @[vga.scala 14:20]
  reg [7:0] ram_1768; // @[vga.scala 14:20]
  reg [7:0] ram_1769; // @[vga.scala 14:20]
  reg [7:0] ram_1770; // @[vga.scala 14:20]
  reg [7:0] ram_1771; // @[vga.scala 14:20]
  reg [7:0] ram_1772; // @[vga.scala 14:20]
  reg [7:0] ram_1773; // @[vga.scala 14:20]
  reg [7:0] ram_1774; // @[vga.scala 14:20]
  reg [7:0] ram_1775; // @[vga.scala 14:20]
  reg [7:0] ram_1776; // @[vga.scala 14:20]
  reg [7:0] ram_1777; // @[vga.scala 14:20]
  reg [7:0] ram_1778; // @[vga.scala 14:20]
  reg [7:0] ram_1779; // @[vga.scala 14:20]
  reg [7:0] ram_1780; // @[vga.scala 14:20]
  reg [7:0] ram_1781; // @[vga.scala 14:20]
  reg [7:0] ram_1782; // @[vga.scala 14:20]
  reg [7:0] ram_1783; // @[vga.scala 14:20]
  reg [7:0] ram_1784; // @[vga.scala 14:20]
  reg [7:0] ram_1785; // @[vga.scala 14:20]
  reg [7:0] ram_1786; // @[vga.scala 14:20]
  reg [7:0] ram_1787; // @[vga.scala 14:20]
  reg [7:0] ram_1788; // @[vga.scala 14:20]
  reg [7:0] ram_1789; // @[vga.scala 14:20]
  reg [7:0] ram_1790; // @[vga.scala 14:20]
  reg [7:0] ram_1791; // @[vga.scala 14:20]
  reg [7:0] ram_1792; // @[vga.scala 14:20]
  reg [7:0] ram_1793; // @[vga.scala 14:20]
  reg [7:0] ram_1794; // @[vga.scala 14:20]
  reg [7:0] ram_1795; // @[vga.scala 14:20]
  reg [7:0] ram_1796; // @[vga.scala 14:20]
  reg [7:0] ram_1797; // @[vga.scala 14:20]
  reg [7:0] ram_1798; // @[vga.scala 14:20]
  reg [7:0] ram_1799; // @[vga.scala 14:20]
  reg [7:0] ram_1800; // @[vga.scala 14:20]
  reg [7:0] ram_1801; // @[vga.scala 14:20]
  reg [7:0] ram_1802; // @[vga.scala 14:20]
  reg [7:0] ram_1803; // @[vga.scala 14:20]
  reg [7:0] ram_1804; // @[vga.scala 14:20]
  reg [7:0] ram_1805; // @[vga.scala 14:20]
  reg [7:0] ram_1806; // @[vga.scala 14:20]
  reg [7:0] ram_1807; // @[vga.scala 14:20]
  reg [7:0] ram_1808; // @[vga.scala 14:20]
  reg [7:0] ram_1809; // @[vga.scala 14:20]
  reg [7:0] ram_1810; // @[vga.scala 14:20]
  reg [7:0] ram_1811; // @[vga.scala 14:20]
  reg [7:0] ram_1812; // @[vga.scala 14:20]
  reg [7:0] ram_1813; // @[vga.scala 14:20]
  reg [7:0] ram_1814; // @[vga.scala 14:20]
  reg [7:0] ram_1815; // @[vga.scala 14:20]
  reg [7:0] ram_1816; // @[vga.scala 14:20]
  reg [7:0] ram_1817; // @[vga.scala 14:20]
  reg [7:0] ram_1818; // @[vga.scala 14:20]
  reg [7:0] ram_1819; // @[vga.scala 14:20]
  reg [7:0] ram_1820; // @[vga.scala 14:20]
  reg [7:0] ram_1821; // @[vga.scala 14:20]
  reg [7:0] ram_1822; // @[vga.scala 14:20]
  reg [7:0] ram_1823; // @[vga.scala 14:20]
  reg [7:0] ram_1824; // @[vga.scala 14:20]
  reg [7:0] ram_1825; // @[vga.scala 14:20]
  reg [7:0] ram_1826; // @[vga.scala 14:20]
  reg [7:0] ram_1827; // @[vga.scala 14:20]
  reg [7:0] ram_1828; // @[vga.scala 14:20]
  reg [7:0] ram_1829; // @[vga.scala 14:20]
  reg [7:0] ram_1830; // @[vga.scala 14:20]
  reg [7:0] ram_1831; // @[vga.scala 14:20]
  reg [7:0] ram_1832; // @[vga.scala 14:20]
  reg [7:0] ram_1833; // @[vga.scala 14:20]
  reg [7:0] ram_1834; // @[vga.scala 14:20]
  reg [7:0] ram_1835; // @[vga.scala 14:20]
  reg [7:0] ram_1836; // @[vga.scala 14:20]
  reg [7:0] ram_1837; // @[vga.scala 14:20]
  reg [7:0] ram_1838; // @[vga.scala 14:20]
  reg [7:0] ram_1839; // @[vga.scala 14:20]
  reg [7:0] ram_1840; // @[vga.scala 14:20]
  reg [7:0] ram_1841; // @[vga.scala 14:20]
  reg [7:0] ram_1842; // @[vga.scala 14:20]
  reg [7:0] ram_1843; // @[vga.scala 14:20]
  reg [7:0] ram_1844; // @[vga.scala 14:20]
  reg [7:0] ram_1845; // @[vga.scala 14:20]
  reg [7:0] ram_1846; // @[vga.scala 14:20]
  reg [7:0] ram_1847; // @[vga.scala 14:20]
  reg [7:0] ram_1848; // @[vga.scala 14:20]
  reg [7:0] ram_1849; // @[vga.scala 14:20]
  reg [7:0] ram_1850; // @[vga.scala 14:20]
  reg [7:0] ram_1851; // @[vga.scala 14:20]
  reg [7:0] ram_1852; // @[vga.scala 14:20]
  reg [7:0] ram_1853; // @[vga.scala 14:20]
  reg [7:0] ram_1854; // @[vga.scala 14:20]
  reg [7:0] ram_1855; // @[vga.scala 14:20]
  reg [7:0] ram_1856; // @[vga.scala 14:20]
  reg [7:0] ram_1857; // @[vga.scala 14:20]
  reg [7:0] ram_1858; // @[vga.scala 14:20]
  reg [7:0] ram_1859; // @[vga.scala 14:20]
  reg [7:0] ram_1860; // @[vga.scala 14:20]
  reg [7:0] ram_1861; // @[vga.scala 14:20]
  reg [7:0] ram_1862; // @[vga.scala 14:20]
  reg [7:0] ram_1863; // @[vga.scala 14:20]
  reg [7:0] ram_1864; // @[vga.scala 14:20]
  reg [7:0] ram_1865; // @[vga.scala 14:20]
  reg [7:0] ram_1866; // @[vga.scala 14:20]
  reg [7:0] ram_1867; // @[vga.scala 14:20]
  reg [7:0] ram_1868; // @[vga.scala 14:20]
  reg [7:0] ram_1869; // @[vga.scala 14:20]
  reg [7:0] ram_1870; // @[vga.scala 14:20]
  reg [7:0] ram_1871; // @[vga.scala 14:20]
  reg [7:0] ram_1872; // @[vga.scala 14:20]
  reg [7:0] ram_1873; // @[vga.scala 14:20]
  reg [7:0] ram_1874; // @[vga.scala 14:20]
  reg [7:0] ram_1875; // @[vga.scala 14:20]
  reg [7:0] ram_1876; // @[vga.scala 14:20]
  reg [7:0] ram_1877; // @[vga.scala 14:20]
  reg [7:0] ram_1878; // @[vga.scala 14:20]
  reg [7:0] ram_1879; // @[vga.scala 14:20]
  reg [7:0] ram_1880; // @[vga.scala 14:20]
  reg [7:0] ram_1881; // @[vga.scala 14:20]
  reg [7:0] ram_1882; // @[vga.scala 14:20]
  reg [7:0] ram_1883; // @[vga.scala 14:20]
  reg [7:0] ram_1884; // @[vga.scala 14:20]
  reg [7:0] ram_1885; // @[vga.scala 14:20]
  reg [7:0] ram_1886; // @[vga.scala 14:20]
  reg [7:0] ram_1887; // @[vga.scala 14:20]
  reg [7:0] ram_1888; // @[vga.scala 14:20]
  reg [7:0] ram_1889; // @[vga.scala 14:20]
  reg [7:0] ram_1890; // @[vga.scala 14:20]
  reg [7:0] ram_1891; // @[vga.scala 14:20]
  reg [7:0] ram_1892; // @[vga.scala 14:20]
  reg [7:0] ram_1893; // @[vga.scala 14:20]
  reg [7:0] ram_1894; // @[vga.scala 14:20]
  reg [7:0] ram_1895; // @[vga.scala 14:20]
  reg [7:0] ram_1896; // @[vga.scala 14:20]
  reg [7:0] ram_1897; // @[vga.scala 14:20]
  reg [7:0] ram_1898; // @[vga.scala 14:20]
  reg [7:0] ram_1899; // @[vga.scala 14:20]
  reg [7:0] ram_1900; // @[vga.scala 14:20]
  reg [7:0] ram_1901; // @[vga.scala 14:20]
  reg [7:0] ram_1902; // @[vga.scala 14:20]
  reg [7:0] ram_1903; // @[vga.scala 14:20]
  reg [7:0] ram_1904; // @[vga.scala 14:20]
  reg [7:0] ram_1905; // @[vga.scala 14:20]
  reg [7:0] ram_1906; // @[vga.scala 14:20]
  reg [7:0] ram_1907; // @[vga.scala 14:20]
  reg [7:0] ram_1908; // @[vga.scala 14:20]
  reg [7:0] ram_1909; // @[vga.scala 14:20]
  reg [7:0] ram_1910; // @[vga.scala 14:20]
  reg [7:0] ram_1911; // @[vga.scala 14:20]
  reg [7:0] ram_1912; // @[vga.scala 14:20]
  reg [7:0] ram_1913; // @[vga.scala 14:20]
  reg [7:0] ram_1914; // @[vga.scala 14:20]
  reg [7:0] ram_1915; // @[vga.scala 14:20]
  reg [7:0] ram_1916; // @[vga.scala 14:20]
  reg [7:0] ram_1917; // @[vga.scala 14:20]
  reg [7:0] ram_1918; // @[vga.scala 14:20]
  reg [7:0] ram_1919; // @[vga.scala 14:20]
  reg [7:0] ram_1920; // @[vga.scala 14:20]
  reg [7:0] ram_1921; // @[vga.scala 14:20]
  reg [7:0] ram_1922; // @[vga.scala 14:20]
  reg [7:0] ram_1923; // @[vga.scala 14:20]
  reg [7:0] ram_1924; // @[vga.scala 14:20]
  reg [7:0] ram_1925; // @[vga.scala 14:20]
  reg [7:0] ram_1926; // @[vga.scala 14:20]
  reg [7:0] ram_1927; // @[vga.scala 14:20]
  reg [7:0] ram_1928; // @[vga.scala 14:20]
  reg [7:0] ram_1929; // @[vga.scala 14:20]
  reg [7:0] ram_1930; // @[vga.scala 14:20]
  reg [7:0] ram_1931; // @[vga.scala 14:20]
  reg [7:0] ram_1932; // @[vga.scala 14:20]
  reg [7:0] ram_1933; // @[vga.scala 14:20]
  reg [7:0] ram_1934; // @[vga.scala 14:20]
  reg [7:0] ram_1935; // @[vga.scala 14:20]
  reg [7:0] ram_1936; // @[vga.scala 14:20]
  reg [7:0] ram_1937; // @[vga.scala 14:20]
  reg [7:0] ram_1938; // @[vga.scala 14:20]
  reg [7:0] ram_1939; // @[vga.scala 14:20]
  reg [7:0] ram_1940; // @[vga.scala 14:20]
  reg [7:0] ram_1941; // @[vga.scala 14:20]
  reg [7:0] ram_1942; // @[vga.scala 14:20]
  reg [7:0] ram_1943; // @[vga.scala 14:20]
  reg [7:0] ram_1944; // @[vga.scala 14:20]
  reg [7:0] ram_1945; // @[vga.scala 14:20]
  reg [7:0] ram_1946; // @[vga.scala 14:20]
  reg [7:0] ram_1947; // @[vga.scala 14:20]
  reg [7:0] ram_1948; // @[vga.scala 14:20]
  reg [7:0] ram_1949; // @[vga.scala 14:20]
  reg [7:0] ram_1950; // @[vga.scala 14:20]
  reg [7:0] ram_1951; // @[vga.scala 14:20]
  reg [7:0] ram_1952; // @[vga.scala 14:20]
  reg [7:0] ram_1953; // @[vga.scala 14:20]
  reg [7:0] ram_1954; // @[vga.scala 14:20]
  reg [7:0] ram_1955; // @[vga.scala 14:20]
  reg [7:0] ram_1956; // @[vga.scala 14:20]
  reg [7:0] ram_1957; // @[vga.scala 14:20]
  reg [7:0] ram_1958; // @[vga.scala 14:20]
  reg [7:0] ram_1959; // @[vga.scala 14:20]
  reg [7:0] ram_1960; // @[vga.scala 14:20]
  reg [7:0] ram_1961; // @[vga.scala 14:20]
  reg [7:0] ram_1962; // @[vga.scala 14:20]
  reg [7:0] ram_1963; // @[vga.scala 14:20]
  reg [7:0] ram_1964; // @[vga.scala 14:20]
  reg [7:0] ram_1965; // @[vga.scala 14:20]
  reg [7:0] ram_1966; // @[vga.scala 14:20]
  reg [7:0] ram_1967; // @[vga.scala 14:20]
  reg [7:0] ram_1968; // @[vga.scala 14:20]
  reg [7:0] ram_1969; // @[vga.scala 14:20]
  reg [7:0] ram_1970; // @[vga.scala 14:20]
  reg [7:0] ram_1971; // @[vga.scala 14:20]
  reg [7:0] ram_1972; // @[vga.scala 14:20]
  reg [7:0] ram_1973; // @[vga.scala 14:20]
  reg [7:0] ram_1974; // @[vga.scala 14:20]
  reg [7:0] ram_1975; // @[vga.scala 14:20]
  reg [7:0] ram_1976; // @[vga.scala 14:20]
  reg [7:0] ram_1977; // @[vga.scala 14:20]
  reg [7:0] ram_1978; // @[vga.scala 14:20]
  reg [7:0] ram_1979; // @[vga.scala 14:20]
  reg [7:0] ram_1980; // @[vga.scala 14:20]
  reg [7:0] ram_1981; // @[vga.scala 14:20]
  reg [7:0] ram_1982; // @[vga.scala 14:20]
  reg [7:0] ram_1983; // @[vga.scala 14:20]
  reg [7:0] ram_1984; // @[vga.scala 14:20]
  reg [7:0] ram_1985; // @[vga.scala 14:20]
  reg [7:0] ram_1986; // @[vga.scala 14:20]
  reg [7:0] ram_1987; // @[vga.scala 14:20]
  reg [7:0] ram_1988; // @[vga.scala 14:20]
  reg [7:0] ram_1989; // @[vga.scala 14:20]
  reg [7:0] ram_1990; // @[vga.scala 14:20]
  reg [7:0] ram_1991; // @[vga.scala 14:20]
  reg [7:0] ram_1992; // @[vga.scala 14:20]
  reg [7:0] ram_1993; // @[vga.scala 14:20]
  reg [7:0] ram_1994; // @[vga.scala 14:20]
  reg [7:0] ram_1995; // @[vga.scala 14:20]
  reg [7:0] ram_1996; // @[vga.scala 14:20]
  reg [7:0] ram_1997; // @[vga.scala 14:20]
  reg [7:0] ram_1998; // @[vga.scala 14:20]
  reg [7:0] ram_1999; // @[vga.scala 14:20]
  reg [7:0] ram_2000; // @[vga.scala 14:20]
  reg [7:0] ram_2001; // @[vga.scala 14:20]
  reg [7:0] ram_2002; // @[vga.scala 14:20]
  reg [7:0] ram_2003; // @[vga.scala 14:20]
  reg [7:0] ram_2004; // @[vga.scala 14:20]
  reg [7:0] ram_2005; // @[vga.scala 14:20]
  reg [7:0] ram_2006; // @[vga.scala 14:20]
  reg [7:0] ram_2007; // @[vga.scala 14:20]
  reg [7:0] ram_2008; // @[vga.scala 14:20]
  reg [7:0] ram_2009; // @[vga.scala 14:20]
  reg [7:0] ram_2010; // @[vga.scala 14:20]
  reg [7:0] ram_2011; // @[vga.scala 14:20]
  reg [7:0] ram_2012; // @[vga.scala 14:20]
  reg [7:0] ram_2013; // @[vga.scala 14:20]
  reg [7:0] ram_2014; // @[vga.scala 14:20]
  reg [7:0] ram_2015; // @[vga.scala 14:20]
  reg [7:0] ram_2016; // @[vga.scala 14:20]
  reg [7:0] ram_2017; // @[vga.scala 14:20]
  reg [7:0] ram_2018; // @[vga.scala 14:20]
  reg [7:0] ram_2019; // @[vga.scala 14:20]
  reg [7:0] ram_2020; // @[vga.scala 14:20]
  reg [7:0] ram_2021; // @[vga.scala 14:20]
  reg [7:0] ram_2022; // @[vga.scala 14:20]
  reg [7:0] ram_2023; // @[vga.scala 14:20]
  reg [7:0] ram_2024; // @[vga.scala 14:20]
  reg [7:0] ram_2025; // @[vga.scala 14:20]
  reg [7:0] ram_2026; // @[vga.scala 14:20]
  reg [7:0] ram_2027; // @[vga.scala 14:20]
  reg [7:0] ram_2028; // @[vga.scala 14:20]
  reg [7:0] ram_2029; // @[vga.scala 14:20]
  reg [7:0] ram_2030; // @[vga.scala 14:20]
  reg [7:0] ram_2031; // @[vga.scala 14:20]
  reg [7:0] ram_2032; // @[vga.scala 14:20]
  reg [7:0] ram_2033; // @[vga.scala 14:20]
  reg [7:0] ram_2034; // @[vga.scala 14:20]
  reg [7:0] ram_2035; // @[vga.scala 14:20]
  reg [7:0] ram_2036; // @[vga.scala 14:20]
  reg [7:0] ram_2037; // @[vga.scala 14:20]
  reg [7:0] ram_2038; // @[vga.scala 14:20]
  reg [7:0] ram_2039; // @[vga.scala 14:20]
  reg [7:0] ram_2040; // @[vga.scala 14:20]
  reg [7:0] ram_2041; // @[vga.scala 14:20]
  reg [7:0] ram_2042; // @[vga.scala 14:20]
  reg [7:0] ram_2043; // @[vga.scala 14:20]
  reg [7:0] ram_2044; // @[vga.scala 14:20]
  reg [7:0] ram_2045; // @[vga.scala 14:20]
  reg [7:0] ram_2046; // @[vga.scala 14:20]
  reg [7:0] ram_2047; // @[vga.scala 14:20]
  reg [7:0] ram_2048; // @[vga.scala 14:20]
  reg [7:0] ram_2049; // @[vga.scala 14:20]
  reg [7:0] ram_2050; // @[vga.scala 14:20]
  reg [7:0] ram_2051; // @[vga.scala 14:20]
  reg [7:0] ram_2052; // @[vga.scala 14:20]
  reg [7:0] ram_2053; // @[vga.scala 14:20]
  reg [7:0] ram_2054; // @[vga.scala 14:20]
  reg [7:0] ram_2055; // @[vga.scala 14:20]
  reg [7:0] ram_2056; // @[vga.scala 14:20]
  reg [7:0] ram_2057; // @[vga.scala 14:20]
  reg [7:0] ram_2058; // @[vga.scala 14:20]
  reg [7:0] ram_2059; // @[vga.scala 14:20]
  reg [7:0] ram_2060; // @[vga.scala 14:20]
  reg [7:0] ram_2061; // @[vga.scala 14:20]
  reg [7:0] ram_2062; // @[vga.scala 14:20]
  reg [7:0] ram_2063; // @[vga.scala 14:20]
  reg [7:0] ram_2064; // @[vga.scala 14:20]
  reg [7:0] ram_2065; // @[vga.scala 14:20]
  reg [7:0] ram_2066; // @[vga.scala 14:20]
  reg [7:0] ram_2067; // @[vga.scala 14:20]
  reg [7:0] ram_2068; // @[vga.scala 14:20]
  reg [7:0] ram_2069; // @[vga.scala 14:20]
  reg [7:0] ram_2070; // @[vga.scala 14:20]
  reg [7:0] ram_2071; // @[vga.scala 14:20]
  reg [7:0] ram_2072; // @[vga.scala 14:20]
  reg [7:0] ram_2073; // @[vga.scala 14:20]
  reg [7:0] ram_2074; // @[vga.scala 14:20]
  reg [7:0] ram_2075; // @[vga.scala 14:20]
  reg [7:0] ram_2076; // @[vga.scala 14:20]
  reg [7:0] ram_2077; // @[vga.scala 14:20]
  reg [7:0] ram_2078; // @[vga.scala 14:20]
  reg [7:0] ram_2079; // @[vga.scala 14:20]
  reg [7:0] ram_2080; // @[vga.scala 14:20]
  reg [7:0] ram_2081; // @[vga.scala 14:20]
  reg [7:0] ram_2082; // @[vga.scala 14:20]
  reg [7:0] ram_2083; // @[vga.scala 14:20]
  reg [7:0] ram_2084; // @[vga.scala 14:20]
  reg [7:0] ram_2085; // @[vga.scala 14:20]
  reg [7:0] ram_2086; // @[vga.scala 14:20]
  reg [7:0] ram_2087; // @[vga.scala 14:20]
  reg [7:0] ram_2088; // @[vga.scala 14:20]
  reg [7:0] ram_2089; // @[vga.scala 14:20]
  reg [7:0] ram_2090; // @[vga.scala 14:20]
  reg [7:0] ram_2091; // @[vga.scala 14:20]
  reg [7:0] ram_2092; // @[vga.scala 14:20]
  reg [7:0] ram_2093; // @[vga.scala 14:20]
  reg [7:0] ram_2094; // @[vga.scala 14:20]
  reg [7:0] ram_2095; // @[vga.scala 14:20]
  reg [7:0] ram_2096; // @[vga.scala 14:20]
  reg [7:0] ram_2097; // @[vga.scala 14:20]
  reg [7:0] ram_2098; // @[vga.scala 14:20]
  reg [7:0] ram_2099; // @[vga.scala 14:20]
  reg [7:0] ram_2100; // @[vga.scala 14:20]
  reg [7:0] ram_2101; // @[vga.scala 14:20]
  reg [7:0] ram_2102; // @[vga.scala 14:20]
  reg [7:0] ram_2103; // @[vga.scala 14:20]
  reg [7:0] ram_2104; // @[vga.scala 14:20]
  reg [7:0] ram_2105; // @[vga.scala 14:20]
  reg [7:0] ram_2106; // @[vga.scala 14:20]
  reg [7:0] ram_2107; // @[vga.scala 14:20]
  reg [7:0] ram_2108; // @[vga.scala 14:20]
  reg [7:0] ram_2109; // @[vga.scala 14:20]
  reg [7:0] ram_2110; // @[vga.scala 14:20]
  reg [7:0] ram_2111; // @[vga.scala 14:20]
  reg [7:0] ram_2112; // @[vga.scala 14:20]
  reg [7:0] ram_2113; // @[vga.scala 14:20]
  reg [7:0] ram_2114; // @[vga.scala 14:20]
  reg [7:0] ram_2115; // @[vga.scala 14:20]
  reg [7:0] ram_2116; // @[vga.scala 14:20]
  reg [7:0] ram_2117; // @[vga.scala 14:20]
  reg [7:0] ram_2118; // @[vga.scala 14:20]
  reg [7:0] ram_2119; // @[vga.scala 14:20]
  reg [7:0] ram_2120; // @[vga.scala 14:20]
  reg [7:0] ram_2121; // @[vga.scala 14:20]
  reg [7:0] ram_2122; // @[vga.scala 14:20]
  reg [7:0] ram_2123; // @[vga.scala 14:20]
  reg [7:0] ram_2124; // @[vga.scala 14:20]
  reg [7:0] ram_2125; // @[vga.scala 14:20]
  reg [7:0] ram_2126; // @[vga.scala 14:20]
  reg [7:0] ram_2127; // @[vga.scala 14:20]
  reg [7:0] ram_2128; // @[vga.scala 14:20]
  reg [7:0] ram_2129; // @[vga.scala 14:20]
  reg [7:0] ram_2130; // @[vga.scala 14:20]
  reg [7:0] ram_2131; // @[vga.scala 14:20]
  reg [7:0] ram_2132; // @[vga.scala 14:20]
  reg [7:0] ram_2133; // @[vga.scala 14:20]
  reg [7:0] ram_2134; // @[vga.scala 14:20]
  reg [7:0] ram_2135; // @[vga.scala 14:20]
  reg [7:0] ram_2136; // @[vga.scala 14:20]
  reg [7:0] ram_2137; // @[vga.scala 14:20]
  reg [7:0] ram_2138; // @[vga.scala 14:20]
  reg [7:0] ram_2139; // @[vga.scala 14:20]
  reg [7:0] ram_2140; // @[vga.scala 14:20]
  reg [7:0] ram_2141; // @[vga.scala 14:20]
  reg [7:0] ram_2142; // @[vga.scala 14:20]
  reg [7:0] ram_2143; // @[vga.scala 14:20]
  reg [7:0] ram_2144; // @[vga.scala 14:20]
  reg [7:0] ram_2145; // @[vga.scala 14:20]
  reg [7:0] ram_2146; // @[vga.scala 14:20]
  reg [7:0] ram_2147; // @[vga.scala 14:20]
  reg [7:0] ram_2148; // @[vga.scala 14:20]
  reg [7:0] ram_2149; // @[vga.scala 14:20]
  reg [7:0] ram_2150; // @[vga.scala 14:20]
  reg [7:0] ram_2151; // @[vga.scala 14:20]
  reg [7:0] ram_2152; // @[vga.scala 14:20]
  reg [7:0] ram_2153; // @[vga.scala 14:20]
  reg [7:0] ram_2154; // @[vga.scala 14:20]
  reg [7:0] ram_2155; // @[vga.scala 14:20]
  reg [7:0] ram_2156; // @[vga.scala 14:20]
  reg [7:0] ram_2157; // @[vga.scala 14:20]
  reg [7:0] ram_2158; // @[vga.scala 14:20]
  reg [7:0] ram_2159; // @[vga.scala 14:20]
  reg [7:0] ram_2160; // @[vga.scala 14:20]
  reg [7:0] index; // @[vga.scala 20:22]
  wire [7:0] _index_T_1 = index + 8'h47; // @[vga.scala 23:26]
  wire [7:0] _GEN_0 = _index_T_1 % 8'h47; // @[vga.scala 23:45]
  wire [6:0] _index_T_4 = _GEN_0[6:0]; // @[vga.scala 23:45]
  wire [7:0] _GEN_8647 = {{1'd0}, _index_T_4}; // @[vga.scala 23:32]
  wire [7:0] _index_T_6 = _index_T_1 - _GEN_8647; // @[vga.scala 23:32]
  wire [8:0] _GEN_8648 = {{1'd0}, index}; // @[vga.scala 25:23 vga.scala 25:23 vga.scala 14:20]
  wire [9:0] _GEN_8904 = {{2'd0}, index}; // @[vga.scala 25:23 vga.scala 25:23 vga.scala 14:20]
  wire [10:0] _GEN_9416 = {{3'd0}, index}; // @[vga.scala 25:23 vga.scala 25:23 vga.scala 14:20]
  wire [11:0] _GEN_10440 = {{4'd0}, index}; // @[vga.scala 25:23 vga.scala 25:23 vga.scala 14:20]
  wire [7:0] _index_T_8 = index + 8'h1; // @[vga.scala 26:25]
  wire [8:0] _T_2 = {{4'd0}, io_v_addr[8:4]}; // @[vga.scala 29:33]
  wire [15:0] _T_3 = _T_2 * 7'h47; // @[vga.scala 29:39]
  wire [9:0] _T_4 = io_h_addr / 10'h9; // @[vga.scala 29:54]
  wire [15:0] _GEN_10554 = {{6'd0}, _T_4}; // @[vga.scala 29:44]
  wire [15:0] _T_6 = _T_3 + _GEN_10554; // @[vga.scala 29:44]
  wire [7:0] _GEN_6486 = 12'h1 == _T_6[11:0] ? ram_1 : ram_0; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6487 = 12'h2 == _T_6[11:0] ? ram_2 : _GEN_6486; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6488 = 12'h3 == _T_6[11:0] ? ram_3 : _GEN_6487; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6489 = 12'h4 == _T_6[11:0] ? ram_4 : _GEN_6488; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6490 = 12'h5 == _T_6[11:0] ? ram_5 : _GEN_6489; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6491 = 12'h6 == _T_6[11:0] ? ram_6 : _GEN_6490; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6492 = 12'h7 == _T_6[11:0] ? ram_7 : _GEN_6491; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6493 = 12'h8 == _T_6[11:0] ? ram_8 : _GEN_6492; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6494 = 12'h9 == _T_6[11:0] ? ram_9 : _GEN_6493; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6495 = 12'ha == _T_6[11:0] ? ram_10 : _GEN_6494; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6496 = 12'hb == _T_6[11:0] ? ram_11 : _GEN_6495; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6497 = 12'hc == _T_6[11:0] ? ram_12 : _GEN_6496; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6498 = 12'hd == _T_6[11:0] ? ram_13 : _GEN_6497; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6499 = 12'he == _T_6[11:0] ? ram_14 : _GEN_6498; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6500 = 12'hf == _T_6[11:0] ? ram_15 : _GEN_6499; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6501 = 12'h10 == _T_6[11:0] ? ram_16 : _GEN_6500; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6502 = 12'h11 == _T_6[11:0] ? ram_17 : _GEN_6501; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6503 = 12'h12 == _T_6[11:0] ? ram_18 : _GEN_6502; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6504 = 12'h13 == _T_6[11:0] ? ram_19 : _GEN_6503; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6505 = 12'h14 == _T_6[11:0] ? ram_20 : _GEN_6504; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6506 = 12'h15 == _T_6[11:0] ? ram_21 : _GEN_6505; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6507 = 12'h16 == _T_6[11:0] ? ram_22 : _GEN_6506; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6508 = 12'h17 == _T_6[11:0] ? ram_23 : _GEN_6507; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6509 = 12'h18 == _T_6[11:0] ? ram_24 : _GEN_6508; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6510 = 12'h19 == _T_6[11:0] ? ram_25 : _GEN_6509; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6511 = 12'h1a == _T_6[11:0] ? ram_26 : _GEN_6510; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6512 = 12'h1b == _T_6[11:0] ? ram_27 : _GEN_6511; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6513 = 12'h1c == _T_6[11:0] ? ram_28 : _GEN_6512; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6514 = 12'h1d == _T_6[11:0] ? ram_29 : _GEN_6513; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6515 = 12'h1e == _T_6[11:0] ? ram_30 : _GEN_6514; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6516 = 12'h1f == _T_6[11:0] ? ram_31 : _GEN_6515; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6517 = 12'h20 == _T_6[11:0] ? ram_32 : _GEN_6516; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6518 = 12'h21 == _T_6[11:0] ? ram_33 : _GEN_6517; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6519 = 12'h22 == _T_6[11:0] ? ram_34 : _GEN_6518; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6520 = 12'h23 == _T_6[11:0] ? ram_35 : _GEN_6519; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6521 = 12'h24 == _T_6[11:0] ? ram_36 : _GEN_6520; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6522 = 12'h25 == _T_6[11:0] ? ram_37 : _GEN_6521; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6523 = 12'h26 == _T_6[11:0] ? ram_38 : _GEN_6522; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6524 = 12'h27 == _T_6[11:0] ? ram_39 : _GEN_6523; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6525 = 12'h28 == _T_6[11:0] ? ram_40 : _GEN_6524; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6526 = 12'h29 == _T_6[11:0] ? ram_41 : _GEN_6525; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6527 = 12'h2a == _T_6[11:0] ? ram_42 : _GEN_6526; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6528 = 12'h2b == _T_6[11:0] ? ram_43 : _GEN_6527; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6529 = 12'h2c == _T_6[11:0] ? ram_44 : _GEN_6528; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6530 = 12'h2d == _T_6[11:0] ? ram_45 : _GEN_6529; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6531 = 12'h2e == _T_6[11:0] ? ram_46 : _GEN_6530; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6532 = 12'h2f == _T_6[11:0] ? ram_47 : _GEN_6531; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6533 = 12'h30 == _T_6[11:0] ? ram_48 : _GEN_6532; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6534 = 12'h31 == _T_6[11:0] ? ram_49 : _GEN_6533; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6535 = 12'h32 == _T_6[11:0] ? ram_50 : _GEN_6534; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6536 = 12'h33 == _T_6[11:0] ? ram_51 : _GEN_6535; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6537 = 12'h34 == _T_6[11:0] ? ram_52 : _GEN_6536; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6538 = 12'h35 == _T_6[11:0] ? ram_53 : _GEN_6537; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6539 = 12'h36 == _T_6[11:0] ? ram_54 : _GEN_6538; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6540 = 12'h37 == _T_6[11:0] ? ram_55 : _GEN_6539; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6541 = 12'h38 == _T_6[11:0] ? ram_56 : _GEN_6540; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6542 = 12'h39 == _T_6[11:0] ? ram_57 : _GEN_6541; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6543 = 12'h3a == _T_6[11:0] ? ram_58 : _GEN_6542; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6544 = 12'h3b == _T_6[11:0] ? ram_59 : _GEN_6543; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6545 = 12'h3c == _T_6[11:0] ? ram_60 : _GEN_6544; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6546 = 12'h3d == _T_6[11:0] ? ram_61 : _GEN_6545; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6547 = 12'h3e == _T_6[11:0] ? ram_62 : _GEN_6546; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6548 = 12'h3f == _T_6[11:0] ? ram_63 : _GEN_6547; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6549 = 12'h40 == _T_6[11:0] ? ram_64 : _GEN_6548; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6550 = 12'h41 == _T_6[11:0] ? ram_65 : _GEN_6549; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6551 = 12'h42 == _T_6[11:0] ? ram_66 : _GEN_6550; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6552 = 12'h43 == _T_6[11:0] ? ram_67 : _GEN_6551; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6553 = 12'h44 == _T_6[11:0] ? ram_68 : _GEN_6552; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6554 = 12'h45 == _T_6[11:0] ? ram_69 : _GEN_6553; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6555 = 12'h46 == _T_6[11:0] ? ram_70 : _GEN_6554; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6556 = 12'h47 == _T_6[11:0] ? ram_71 : _GEN_6555; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6557 = 12'h48 == _T_6[11:0] ? ram_72 : _GEN_6556; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6558 = 12'h49 == _T_6[11:0] ? ram_73 : _GEN_6557; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6559 = 12'h4a == _T_6[11:0] ? ram_74 : _GEN_6558; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6560 = 12'h4b == _T_6[11:0] ? ram_75 : _GEN_6559; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6561 = 12'h4c == _T_6[11:0] ? ram_76 : _GEN_6560; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6562 = 12'h4d == _T_6[11:0] ? ram_77 : _GEN_6561; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6563 = 12'h4e == _T_6[11:0] ? ram_78 : _GEN_6562; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6564 = 12'h4f == _T_6[11:0] ? ram_79 : _GEN_6563; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6565 = 12'h50 == _T_6[11:0] ? ram_80 : _GEN_6564; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6566 = 12'h51 == _T_6[11:0] ? ram_81 : _GEN_6565; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6567 = 12'h52 == _T_6[11:0] ? ram_82 : _GEN_6566; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6568 = 12'h53 == _T_6[11:0] ? ram_83 : _GEN_6567; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6569 = 12'h54 == _T_6[11:0] ? ram_84 : _GEN_6568; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6570 = 12'h55 == _T_6[11:0] ? ram_85 : _GEN_6569; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6571 = 12'h56 == _T_6[11:0] ? ram_86 : _GEN_6570; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6572 = 12'h57 == _T_6[11:0] ? ram_87 : _GEN_6571; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6573 = 12'h58 == _T_6[11:0] ? ram_88 : _GEN_6572; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6574 = 12'h59 == _T_6[11:0] ? ram_89 : _GEN_6573; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6575 = 12'h5a == _T_6[11:0] ? ram_90 : _GEN_6574; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6576 = 12'h5b == _T_6[11:0] ? ram_91 : _GEN_6575; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6577 = 12'h5c == _T_6[11:0] ? ram_92 : _GEN_6576; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6578 = 12'h5d == _T_6[11:0] ? ram_93 : _GEN_6577; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6579 = 12'h5e == _T_6[11:0] ? ram_94 : _GEN_6578; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6580 = 12'h5f == _T_6[11:0] ? ram_95 : _GEN_6579; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6581 = 12'h60 == _T_6[11:0] ? ram_96 : _GEN_6580; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6582 = 12'h61 == _T_6[11:0] ? ram_97 : _GEN_6581; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6583 = 12'h62 == _T_6[11:0] ? ram_98 : _GEN_6582; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6584 = 12'h63 == _T_6[11:0] ? ram_99 : _GEN_6583; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6585 = 12'h64 == _T_6[11:0] ? ram_100 : _GEN_6584; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6586 = 12'h65 == _T_6[11:0] ? ram_101 : _GEN_6585; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6587 = 12'h66 == _T_6[11:0] ? ram_102 : _GEN_6586; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6588 = 12'h67 == _T_6[11:0] ? ram_103 : _GEN_6587; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6589 = 12'h68 == _T_6[11:0] ? ram_104 : _GEN_6588; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6590 = 12'h69 == _T_6[11:0] ? ram_105 : _GEN_6589; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6591 = 12'h6a == _T_6[11:0] ? ram_106 : _GEN_6590; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6592 = 12'h6b == _T_6[11:0] ? ram_107 : _GEN_6591; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6593 = 12'h6c == _T_6[11:0] ? ram_108 : _GEN_6592; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6594 = 12'h6d == _T_6[11:0] ? ram_109 : _GEN_6593; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6595 = 12'h6e == _T_6[11:0] ? ram_110 : _GEN_6594; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6596 = 12'h6f == _T_6[11:0] ? ram_111 : _GEN_6595; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6597 = 12'h70 == _T_6[11:0] ? ram_112 : _GEN_6596; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6598 = 12'h71 == _T_6[11:0] ? ram_113 : _GEN_6597; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6599 = 12'h72 == _T_6[11:0] ? ram_114 : _GEN_6598; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6600 = 12'h73 == _T_6[11:0] ? ram_115 : _GEN_6599; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6601 = 12'h74 == _T_6[11:0] ? ram_116 : _GEN_6600; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6602 = 12'h75 == _T_6[11:0] ? ram_117 : _GEN_6601; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6603 = 12'h76 == _T_6[11:0] ? ram_118 : _GEN_6602; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6604 = 12'h77 == _T_6[11:0] ? ram_119 : _GEN_6603; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6605 = 12'h78 == _T_6[11:0] ? ram_120 : _GEN_6604; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6606 = 12'h79 == _T_6[11:0] ? ram_121 : _GEN_6605; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6607 = 12'h7a == _T_6[11:0] ? ram_122 : _GEN_6606; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6608 = 12'h7b == _T_6[11:0] ? ram_123 : _GEN_6607; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6609 = 12'h7c == _T_6[11:0] ? ram_124 : _GEN_6608; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6610 = 12'h7d == _T_6[11:0] ? ram_125 : _GEN_6609; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6611 = 12'h7e == _T_6[11:0] ? ram_126 : _GEN_6610; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6612 = 12'h7f == _T_6[11:0] ? ram_127 : _GEN_6611; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6613 = 12'h80 == _T_6[11:0] ? ram_128 : _GEN_6612; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6614 = 12'h81 == _T_6[11:0] ? ram_129 : _GEN_6613; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6615 = 12'h82 == _T_6[11:0] ? ram_130 : _GEN_6614; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6616 = 12'h83 == _T_6[11:0] ? ram_131 : _GEN_6615; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6617 = 12'h84 == _T_6[11:0] ? ram_132 : _GEN_6616; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6618 = 12'h85 == _T_6[11:0] ? ram_133 : _GEN_6617; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6619 = 12'h86 == _T_6[11:0] ? ram_134 : _GEN_6618; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6620 = 12'h87 == _T_6[11:0] ? ram_135 : _GEN_6619; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6621 = 12'h88 == _T_6[11:0] ? ram_136 : _GEN_6620; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6622 = 12'h89 == _T_6[11:0] ? ram_137 : _GEN_6621; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6623 = 12'h8a == _T_6[11:0] ? ram_138 : _GEN_6622; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6624 = 12'h8b == _T_6[11:0] ? ram_139 : _GEN_6623; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6625 = 12'h8c == _T_6[11:0] ? ram_140 : _GEN_6624; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6626 = 12'h8d == _T_6[11:0] ? ram_141 : _GEN_6625; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6627 = 12'h8e == _T_6[11:0] ? ram_142 : _GEN_6626; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6628 = 12'h8f == _T_6[11:0] ? ram_143 : _GEN_6627; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6629 = 12'h90 == _T_6[11:0] ? ram_144 : _GEN_6628; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6630 = 12'h91 == _T_6[11:0] ? ram_145 : _GEN_6629; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6631 = 12'h92 == _T_6[11:0] ? ram_146 : _GEN_6630; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6632 = 12'h93 == _T_6[11:0] ? ram_147 : _GEN_6631; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6633 = 12'h94 == _T_6[11:0] ? ram_148 : _GEN_6632; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6634 = 12'h95 == _T_6[11:0] ? ram_149 : _GEN_6633; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6635 = 12'h96 == _T_6[11:0] ? ram_150 : _GEN_6634; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6636 = 12'h97 == _T_6[11:0] ? ram_151 : _GEN_6635; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6637 = 12'h98 == _T_6[11:0] ? ram_152 : _GEN_6636; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6638 = 12'h99 == _T_6[11:0] ? ram_153 : _GEN_6637; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6639 = 12'h9a == _T_6[11:0] ? ram_154 : _GEN_6638; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6640 = 12'h9b == _T_6[11:0] ? ram_155 : _GEN_6639; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6641 = 12'h9c == _T_6[11:0] ? ram_156 : _GEN_6640; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6642 = 12'h9d == _T_6[11:0] ? ram_157 : _GEN_6641; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6643 = 12'h9e == _T_6[11:0] ? ram_158 : _GEN_6642; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6644 = 12'h9f == _T_6[11:0] ? ram_159 : _GEN_6643; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6645 = 12'ha0 == _T_6[11:0] ? ram_160 : _GEN_6644; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6646 = 12'ha1 == _T_6[11:0] ? ram_161 : _GEN_6645; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6647 = 12'ha2 == _T_6[11:0] ? ram_162 : _GEN_6646; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6648 = 12'ha3 == _T_6[11:0] ? ram_163 : _GEN_6647; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6649 = 12'ha4 == _T_6[11:0] ? ram_164 : _GEN_6648; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6650 = 12'ha5 == _T_6[11:0] ? ram_165 : _GEN_6649; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6651 = 12'ha6 == _T_6[11:0] ? ram_166 : _GEN_6650; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6652 = 12'ha7 == _T_6[11:0] ? ram_167 : _GEN_6651; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6653 = 12'ha8 == _T_6[11:0] ? ram_168 : _GEN_6652; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6654 = 12'ha9 == _T_6[11:0] ? ram_169 : _GEN_6653; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6655 = 12'haa == _T_6[11:0] ? ram_170 : _GEN_6654; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6656 = 12'hab == _T_6[11:0] ? ram_171 : _GEN_6655; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6657 = 12'hac == _T_6[11:0] ? ram_172 : _GEN_6656; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6658 = 12'had == _T_6[11:0] ? ram_173 : _GEN_6657; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6659 = 12'hae == _T_6[11:0] ? ram_174 : _GEN_6658; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6660 = 12'haf == _T_6[11:0] ? ram_175 : _GEN_6659; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6661 = 12'hb0 == _T_6[11:0] ? ram_176 : _GEN_6660; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6662 = 12'hb1 == _T_6[11:0] ? ram_177 : _GEN_6661; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6663 = 12'hb2 == _T_6[11:0] ? ram_178 : _GEN_6662; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6664 = 12'hb3 == _T_6[11:0] ? ram_179 : _GEN_6663; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6665 = 12'hb4 == _T_6[11:0] ? ram_180 : _GEN_6664; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6666 = 12'hb5 == _T_6[11:0] ? ram_181 : _GEN_6665; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6667 = 12'hb6 == _T_6[11:0] ? ram_182 : _GEN_6666; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6668 = 12'hb7 == _T_6[11:0] ? ram_183 : _GEN_6667; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6669 = 12'hb8 == _T_6[11:0] ? ram_184 : _GEN_6668; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6670 = 12'hb9 == _T_6[11:0] ? ram_185 : _GEN_6669; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6671 = 12'hba == _T_6[11:0] ? ram_186 : _GEN_6670; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6672 = 12'hbb == _T_6[11:0] ? ram_187 : _GEN_6671; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6673 = 12'hbc == _T_6[11:0] ? ram_188 : _GEN_6672; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6674 = 12'hbd == _T_6[11:0] ? ram_189 : _GEN_6673; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6675 = 12'hbe == _T_6[11:0] ? ram_190 : _GEN_6674; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6676 = 12'hbf == _T_6[11:0] ? ram_191 : _GEN_6675; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6677 = 12'hc0 == _T_6[11:0] ? ram_192 : _GEN_6676; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6678 = 12'hc1 == _T_6[11:0] ? ram_193 : _GEN_6677; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6679 = 12'hc2 == _T_6[11:0] ? ram_194 : _GEN_6678; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6680 = 12'hc3 == _T_6[11:0] ? ram_195 : _GEN_6679; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6681 = 12'hc4 == _T_6[11:0] ? ram_196 : _GEN_6680; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6682 = 12'hc5 == _T_6[11:0] ? ram_197 : _GEN_6681; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6683 = 12'hc6 == _T_6[11:0] ? ram_198 : _GEN_6682; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6684 = 12'hc7 == _T_6[11:0] ? ram_199 : _GEN_6683; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6685 = 12'hc8 == _T_6[11:0] ? ram_200 : _GEN_6684; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6686 = 12'hc9 == _T_6[11:0] ? ram_201 : _GEN_6685; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6687 = 12'hca == _T_6[11:0] ? ram_202 : _GEN_6686; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6688 = 12'hcb == _T_6[11:0] ? ram_203 : _GEN_6687; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6689 = 12'hcc == _T_6[11:0] ? ram_204 : _GEN_6688; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6690 = 12'hcd == _T_6[11:0] ? ram_205 : _GEN_6689; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6691 = 12'hce == _T_6[11:0] ? ram_206 : _GEN_6690; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6692 = 12'hcf == _T_6[11:0] ? ram_207 : _GEN_6691; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6693 = 12'hd0 == _T_6[11:0] ? ram_208 : _GEN_6692; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6694 = 12'hd1 == _T_6[11:0] ? ram_209 : _GEN_6693; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6695 = 12'hd2 == _T_6[11:0] ? ram_210 : _GEN_6694; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6696 = 12'hd3 == _T_6[11:0] ? ram_211 : _GEN_6695; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6697 = 12'hd4 == _T_6[11:0] ? ram_212 : _GEN_6696; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6698 = 12'hd5 == _T_6[11:0] ? ram_213 : _GEN_6697; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6699 = 12'hd6 == _T_6[11:0] ? ram_214 : _GEN_6698; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6700 = 12'hd7 == _T_6[11:0] ? ram_215 : _GEN_6699; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6701 = 12'hd8 == _T_6[11:0] ? ram_216 : _GEN_6700; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6702 = 12'hd9 == _T_6[11:0] ? ram_217 : _GEN_6701; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6703 = 12'hda == _T_6[11:0] ? ram_218 : _GEN_6702; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6704 = 12'hdb == _T_6[11:0] ? ram_219 : _GEN_6703; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6705 = 12'hdc == _T_6[11:0] ? ram_220 : _GEN_6704; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6706 = 12'hdd == _T_6[11:0] ? ram_221 : _GEN_6705; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6707 = 12'hde == _T_6[11:0] ? ram_222 : _GEN_6706; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6708 = 12'hdf == _T_6[11:0] ? ram_223 : _GEN_6707; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6709 = 12'he0 == _T_6[11:0] ? ram_224 : _GEN_6708; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6710 = 12'he1 == _T_6[11:0] ? ram_225 : _GEN_6709; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6711 = 12'he2 == _T_6[11:0] ? ram_226 : _GEN_6710; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6712 = 12'he3 == _T_6[11:0] ? ram_227 : _GEN_6711; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6713 = 12'he4 == _T_6[11:0] ? ram_228 : _GEN_6712; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6714 = 12'he5 == _T_6[11:0] ? ram_229 : _GEN_6713; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6715 = 12'he6 == _T_6[11:0] ? ram_230 : _GEN_6714; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6716 = 12'he7 == _T_6[11:0] ? ram_231 : _GEN_6715; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6717 = 12'he8 == _T_6[11:0] ? ram_232 : _GEN_6716; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6718 = 12'he9 == _T_6[11:0] ? ram_233 : _GEN_6717; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6719 = 12'hea == _T_6[11:0] ? ram_234 : _GEN_6718; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6720 = 12'heb == _T_6[11:0] ? ram_235 : _GEN_6719; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6721 = 12'hec == _T_6[11:0] ? ram_236 : _GEN_6720; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6722 = 12'hed == _T_6[11:0] ? ram_237 : _GEN_6721; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6723 = 12'hee == _T_6[11:0] ? ram_238 : _GEN_6722; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6724 = 12'hef == _T_6[11:0] ? ram_239 : _GEN_6723; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6725 = 12'hf0 == _T_6[11:0] ? ram_240 : _GEN_6724; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6726 = 12'hf1 == _T_6[11:0] ? ram_241 : _GEN_6725; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6727 = 12'hf2 == _T_6[11:0] ? ram_242 : _GEN_6726; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6728 = 12'hf3 == _T_6[11:0] ? ram_243 : _GEN_6727; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6729 = 12'hf4 == _T_6[11:0] ? ram_244 : _GEN_6728; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6730 = 12'hf5 == _T_6[11:0] ? ram_245 : _GEN_6729; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6731 = 12'hf6 == _T_6[11:0] ? ram_246 : _GEN_6730; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6732 = 12'hf7 == _T_6[11:0] ? ram_247 : _GEN_6731; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6733 = 12'hf8 == _T_6[11:0] ? ram_248 : _GEN_6732; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6734 = 12'hf9 == _T_6[11:0] ? ram_249 : _GEN_6733; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6735 = 12'hfa == _T_6[11:0] ? ram_250 : _GEN_6734; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6736 = 12'hfb == _T_6[11:0] ? ram_251 : _GEN_6735; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6737 = 12'hfc == _T_6[11:0] ? ram_252 : _GEN_6736; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6738 = 12'hfd == _T_6[11:0] ? ram_253 : _GEN_6737; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6739 = 12'hfe == _T_6[11:0] ? ram_254 : _GEN_6738; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6740 = 12'hff == _T_6[11:0] ? ram_255 : _GEN_6739; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6741 = 12'h100 == _T_6[11:0] ? ram_256 : _GEN_6740; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6742 = 12'h101 == _T_6[11:0] ? ram_257 : _GEN_6741; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6743 = 12'h102 == _T_6[11:0] ? ram_258 : _GEN_6742; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6744 = 12'h103 == _T_6[11:0] ? ram_259 : _GEN_6743; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6745 = 12'h104 == _T_6[11:0] ? ram_260 : _GEN_6744; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6746 = 12'h105 == _T_6[11:0] ? ram_261 : _GEN_6745; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6747 = 12'h106 == _T_6[11:0] ? ram_262 : _GEN_6746; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6748 = 12'h107 == _T_6[11:0] ? ram_263 : _GEN_6747; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6749 = 12'h108 == _T_6[11:0] ? ram_264 : _GEN_6748; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6750 = 12'h109 == _T_6[11:0] ? ram_265 : _GEN_6749; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6751 = 12'h10a == _T_6[11:0] ? ram_266 : _GEN_6750; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6752 = 12'h10b == _T_6[11:0] ? ram_267 : _GEN_6751; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6753 = 12'h10c == _T_6[11:0] ? ram_268 : _GEN_6752; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6754 = 12'h10d == _T_6[11:0] ? ram_269 : _GEN_6753; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6755 = 12'h10e == _T_6[11:0] ? ram_270 : _GEN_6754; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6756 = 12'h10f == _T_6[11:0] ? ram_271 : _GEN_6755; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6757 = 12'h110 == _T_6[11:0] ? ram_272 : _GEN_6756; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6758 = 12'h111 == _T_6[11:0] ? ram_273 : _GEN_6757; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6759 = 12'h112 == _T_6[11:0] ? ram_274 : _GEN_6758; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6760 = 12'h113 == _T_6[11:0] ? ram_275 : _GEN_6759; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6761 = 12'h114 == _T_6[11:0] ? ram_276 : _GEN_6760; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6762 = 12'h115 == _T_6[11:0] ? ram_277 : _GEN_6761; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6763 = 12'h116 == _T_6[11:0] ? ram_278 : _GEN_6762; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6764 = 12'h117 == _T_6[11:0] ? ram_279 : _GEN_6763; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6765 = 12'h118 == _T_6[11:0] ? ram_280 : _GEN_6764; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6766 = 12'h119 == _T_6[11:0] ? ram_281 : _GEN_6765; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6767 = 12'h11a == _T_6[11:0] ? ram_282 : _GEN_6766; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6768 = 12'h11b == _T_6[11:0] ? ram_283 : _GEN_6767; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6769 = 12'h11c == _T_6[11:0] ? ram_284 : _GEN_6768; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6770 = 12'h11d == _T_6[11:0] ? ram_285 : _GEN_6769; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6771 = 12'h11e == _T_6[11:0] ? ram_286 : _GEN_6770; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6772 = 12'h11f == _T_6[11:0] ? ram_287 : _GEN_6771; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6773 = 12'h120 == _T_6[11:0] ? ram_288 : _GEN_6772; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6774 = 12'h121 == _T_6[11:0] ? ram_289 : _GEN_6773; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6775 = 12'h122 == _T_6[11:0] ? ram_290 : _GEN_6774; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6776 = 12'h123 == _T_6[11:0] ? ram_291 : _GEN_6775; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6777 = 12'h124 == _T_6[11:0] ? ram_292 : _GEN_6776; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6778 = 12'h125 == _T_6[11:0] ? ram_293 : _GEN_6777; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6779 = 12'h126 == _T_6[11:0] ? ram_294 : _GEN_6778; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6780 = 12'h127 == _T_6[11:0] ? ram_295 : _GEN_6779; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6781 = 12'h128 == _T_6[11:0] ? ram_296 : _GEN_6780; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6782 = 12'h129 == _T_6[11:0] ? ram_297 : _GEN_6781; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6783 = 12'h12a == _T_6[11:0] ? ram_298 : _GEN_6782; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6784 = 12'h12b == _T_6[11:0] ? ram_299 : _GEN_6783; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6785 = 12'h12c == _T_6[11:0] ? ram_300 : _GEN_6784; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6786 = 12'h12d == _T_6[11:0] ? ram_301 : _GEN_6785; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6787 = 12'h12e == _T_6[11:0] ? ram_302 : _GEN_6786; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6788 = 12'h12f == _T_6[11:0] ? ram_303 : _GEN_6787; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6789 = 12'h130 == _T_6[11:0] ? ram_304 : _GEN_6788; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6790 = 12'h131 == _T_6[11:0] ? ram_305 : _GEN_6789; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6791 = 12'h132 == _T_6[11:0] ? ram_306 : _GEN_6790; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6792 = 12'h133 == _T_6[11:0] ? ram_307 : _GEN_6791; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6793 = 12'h134 == _T_6[11:0] ? ram_308 : _GEN_6792; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6794 = 12'h135 == _T_6[11:0] ? ram_309 : _GEN_6793; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6795 = 12'h136 == _T_6[11:0] ? ram_310 : _GEN_6794; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6796 = 12'h137 == _T_6[11:0] ? ram_311 : _GEN_6795; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6797 = 12'h138 == _T_6[11:0] ? ram_312 : _GEN_6796; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6798 = 12'h139 == _T_6[11:0] ? ram_313 : _GEN_6797; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6799 = 12'h13a == _T_6[11:0] ? ram_314 : _GEN_6798; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6800 = 12'h13b == _T_6[11:0] ? ram_315 : _GEN_6799; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6801 = 12'h13c == _T_6[11:0] ? ram_316 : _GEN_6800; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6802 = 12'h13d == _T_6[11:0] ? ram_317 : _GEN_6801; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6803 = 12'h13e == _T_6[11:0] ? ram_318 : _GEN_6802; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6804 = 12'h13f == _T_6[11:0] ? ram_319 : _GEN_6803; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6805 = 12'h140 == _T_6[11:0] ? ram_320 : _GEN_6804; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6806 = 12'h141 == _T_6[11:0] ? ram_321 : _GEN_6805; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6807 = 12'h142 == _T_6[11:0] ? ram_322 : _GEN_6806; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6808 = 12'h143 == _T_6[11:0] ? ram_323 : _GEN_6807; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6809 = 12'h144 == _T_6[11:0] ? ram_324 : _GEN_6808; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6810 = 12'h145 == _T_6[11:0] ? ram_325 : _GEN_6809; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6811 = 12'h146 == _T_6[11:0] ? ram_326 : _GEN_6810; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6812 = 12'h147 == _T_6[11:0] ? ram_327 : _GEN_6811; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6813 = 12'h148 == _T_6[11:0] ? ram_328 : _GEN_6812; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6814 = 12'h149 == _T_6[11:0] ? ram_329 : _GEN_6813; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6815 = 12'h14a == _T_6[11:0] ? ram_330 : _GEN_6814; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6816 = 12'h14b == _T_6[11:0] ? ram_331 : _GEN_6815; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6817 = 12'h14c == _T_6[11:0] ? ram_332 : _GEN_6816; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6818 = 12'h14d == _T_6[11:0] ? ram_333 : _GEN_6817; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6819 = 12'h14e == _T_6[11:0] ? ram_334 : _GEN_6818; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6820 = 12'h14f == _T_6[11:0] ? ram_335 : _GEN_6819; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6821 = 12'h150 == _T_6[11:0] ? ram_336 : _GEN_6820; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6822 = 12'h151 == _T_6[11:0] ? ram_337 : _GEN_6821; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6823 = 12'h152 == _T_6[11:0] ? ram_338 : _GEN_6822; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6824 = 12'h153 == _T_6[11:0] ? ram_339 : _GEN_6823; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6825 = 12'h154 == _T_6[11:0] ? ram_340 : _GEN_6824; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6826 = 12'h155 == _T_6[11:0] ? ram_341 : _GEN_6825; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6827 = 12'h156 == _T_6[11:0] ? ram_342 : _GEN_6826; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6828 = 12'h157 == _T_6[11:0] ? ram_343 : _GEN_6827; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6829 = 12'h158 == _T_6[11:0] ? ram_344 : _GEN_6828; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6830 = 12'h159 == _T_6[11:0] ? ram_345 : _GEN_6829; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6831 = 12'h15a == _T_6[11:0] ? ram_346 : _GEN_6830; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6832 = 12'h15b == _T_6[11:0] ? ram_347 : _GEN_6831; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6833 = 12'h15c == _T_6[11:0] ? ram_348 : _GEN_6832; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6834 = 12'h15d == _T_6[11:0] ? ram_349 : _GEN_6833; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6835 = 12'h15e == _T_6[11:0] ? ram_350 : _GEN_6834; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6836 = 12'h15f == _T_6[11:0] ? ram_351 : _GEN_6835; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6837 = 12'h160 == _T_6[11:0] ? ram_352 : _GEN_6836; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6838 = 12'h161 == _T_6[11:0] ? ram_353 : _GEN_6837; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6839 = 12'h162 == _T_6[11:0] ? ram_354 : _GEN_6838; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6840 = 12'h163 == _T_6[11:0] ? ram_355 : _GEN_6839; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6841 = 12'h164 == _T_6[11:0] ? ram_356 : _GEN_6840; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6842 = 12'h165 == _T_6[11:0] ? ram_357 : _GEN_6841; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6843 = 12'h166 == _T_6[11:0] ? ram_358 : _GEN_6842; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6844 = 12'h167 == _T_6[11:0] ? ram_359 : _GEN_6843; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6845 = 12'h168 == _T_6[11:0] ? ram_360 : _GEN_6844; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6846 = 12'h169 == _T_6[11:0] ? ram_361 : _GEN_6845; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6847 = 12'h16a == _T_6[11:0] ? ram_362 : _GEN_6846; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6848 = 12'h16b == _T_6[11:0] ? ram_363 : _GEN_6847; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6849 = 12'h16c == _T_6[11:0] ? ram_364 : _GEN_6848; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6850 = 12'h16d == _T_6[11:0] ? ram_365 : _GEN_6849; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6851 = 12'h16e == _T_6[11:0] ? ram_366 : _GEN_6850; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6852 = 12'h16f == _T_6[11:0] ? ram_367 : _GEN_6851; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6853 = 12'h170 == _T_6[11:0] ? ram_368 : _GEN_6852; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6854 = 12'h171 == _T_6[11:0] ? ram_369 : _GEN_6853; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6855 = 12'h172 == _T_6[11:0] ? ram_370 : _GEN_6854; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6856 = 12'h173 == _T_6[11:0] ? ram_371 : _GEN_6855; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6857 = 12'h174 == _T_6[11:0] ? ram_372 : _GEN_6856; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6858 = 12'h175 == _T_6[11:0] ? ram_373 : _GEN_6857; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6859 = 12'h176 == _T_6[11:0] ? ram_374 : _GEN_6858; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6860 = 12'h177 == _T_6[11:0] ? ram_375 : _GEN_6859; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6861 = 12'h178 == _T_6[11:0] ? ram_376 : _GEN_6860; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6862 = 12'h179 == _T_6[11:0] ? ram_377 : _GEN_6861; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6863 = 12'h17a == _T_6[11:0] ? ram_378 : _GEN_6862; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6864 = 12'h17b == _T_6[11:0] ? ram_379 : _GEN_6863; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6865 = 12'h17c == _T_6[11:0] ? ram_380 : _GEN_6864; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6866 = 12'h17d == _T_6[11:0] ? ram_381 : _GEN_6865; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6867 = 12'h17e == _T_6[11:0] ? ram_382 : _GEN_6866; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6868 = 12'h17f == _T_6[11:0] ? ram_383 : _GEN_6867; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6869 = 12'h180 == _T_6[11:0] ? ram_384 : _GEN_6868; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6870 = 12'h181 == _T_6[11:0] ? ram_385 : _GEN_6869; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6871 = 12'h182 == _T_6[11:0] ? ram_386 : _GEN_6870; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6872 = 12'h183 == _T_6[11:0] ? ram_387 : _GEN_6871; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6873 = 12'h184 == _T_6[11:0] ? ram_388 : _GEN_6872; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6874 = 12'h185 == _T_6[11:0] ? ram_389 : _GEN_6873; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6875 = 12'h186 == _T_6[11:0] ? ram_390 : _GEN_6874; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6876 = 12'h187 == _T_6[11:0] ? ram_391 : _GEN_6875; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6877 = 12'h188 == _T_6[11:0] ? ram_392 : _GEN_6876; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6878 = 12'h189 == _T_6[11:0] ? ram_393 : _GEN_6877; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6879 = 12'h18a == _T_6[11:0] ? ram_394 : _GEN_6878; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6880 = 12'h18b == _T_6[11:0] ? ram_395 : _GEN_6879; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6881 = 12'h18c == _T_6[11:0] ? ram_396 : _GEN_6880; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6882 = 12'h18d == _T_6[11:0] ? ram_397 : _GEN_6881; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6883 = 12'h18e == _T_6[11:0] ? ram_398 : _GEN_6882; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6884 = 12'h18f == _T_6[11:0] ? ram_399 : _GEN_6883; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6885 = 12'h190 == _T_6[11:0] ? ram_400 : _GEN_6884; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6886 = 12'h191 == _T_6[11:0] ? ram_401 : _GEN_6885; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6887 = 12'h192 == _T_6[11:0] ? ram_402 : _GEN_6886; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6888 = 12'h193 == _T_6[11:0] ? ram_403 : _GEN_6887; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6889 = 12'h194 == _T_6[11:0] ? ram_404 : _GEN_6888; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6890 = 12'h195 == _T_6[11:0] ? ram_405 : _GEN_6889; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6891 = 12'h196 == _T_6[11:0] ? ram_406 : _GEN_6890; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6892 = 12'h197 == _T_6[11:0] ? ram_407 : _GEN_6891; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6893 = 12'h198 == _T_6[11:0] ? ram_408 : _GEN_6892; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6894 = 12'h199 == _T_6[11:0] ? ram_409 : _GEN_6893; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6895 = 12'h19a == _T_6[11:0] ? ram_410 : _GEN_6894; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6896 = 12'h19b == _T_6[11:0] ? ram_411 : _GEN_6895; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6897 = 12'h19c == _T_6[11:0] ? ram_412 : _GEN_6896; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6898 = 12'h19d == _T_6[11:0] ? ram_413 : _GEN_6897; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6899 = 12'h19e == _T_6[11:0] ? ram_414 : _GEN_6898; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6900 = 12'h19f == _T_6[11:0] ? ram_415 : _GEN_6899; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6901 = 12'h1a0 == _T_6[11:0] ? ram_416 : _GEN_6900; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6902 = 12'h1a1 == _T_6[11:0] ? ram_417 : _GEN_6901; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6903 = 12'h1a2 == _T_6[11:0] ? ram_418 : _GEN_6902; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6904 = 12'h1a3 == _T_6[11:0] ? ram_419 : _GEN_6903; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6905 = 12'h1a4 == _T_6[11:0] ? ram_420 : _GEN_6904; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6906 = 12'h1a5 == _T_6[11:0] ? ram_421 : _GEN_6905; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6907 = 12'h1a6 == _T_6[11:0] ? ram_422 : _GEN_6906; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6908 = 12'h1a7 == _T_6[11:0] ? ram_423 : _GEN_6907; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6909 = 12'h1a8 == _T_6[11:0] ? ram_424 : _GEN_6908; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6910 = 12'h1a9 == _T_6[11:0] ? ram_425 : _GEN_6909; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6911 = 12'h1aa == _T_6[11:0] ? ram_426 : _GEN_6910; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6912 = 12'h1ab == _T_6[11:0] ? ram_427 : _GEN_6911; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6913 = 12'h1ac == _T_6[11:0] ? ram_428 : _GEN_6912; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6914 = 12'h1ad == _T_6[11:0] ? ram_429 : _GEN_6913; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6915 = 12'h1ae == _T_6[11:0] ? ram_430 : _GEN_6914; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6916 = 12'h1af == _T_6[11:0] ? ram_431 : _GEN_6915; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6917 = 12'h1b0 == _T_6[11:0] ? ram_432 : _GEN_6916; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6918 = 12'h1b1 == _T_6[11:0] ? ram_433 : _GEN_6917; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6919 = 12'h1b2 == _T_6[11:0] ? ram_434 : _GEN_6918; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6920 = 12'h1b3 == _T_6[11:0] ? ram_435 : _GEN_6919; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6921 = 12'h1b4 == _T_6[11:0] ? ram_436 : _GEN_6920; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6922 = 12'h1b5 == _T_6[11:0] ? ram_437 : _GEN_6921; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6923 = 12'h1b6 == _T_6[11:0] ? ram_438 : _GEN_6922; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6924 = 12'h1b7 == _T_6[11:0] ? ram_439 : _GEN_6923; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6925 = 12'h1b8 == _T_6[11:0] ? ram_440 : _GEN_6924; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6926 = 12'h1b9 == _T_6[11:0] ? ram_441 : _GEN_6925; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6927 = 12'h1ba == _T_6[11:0] ? ram_442 : _GEN_6926; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6928 = 12'h1bb == _T_6[11:0] ? ram_443 : _GEN_6927; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6929 = 12'h1bc == _T_6[11:0] ? ram_444 : _GEN_6928; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6930 = 12'h1bd == _T_6[11:0] ? ram_445 : _GEN_6929; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6931 = 12'h1be == _T_6[11:0] ? ram_446 : _GEN_6930; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6932 = 12'h1bf == _T_6[11:0] ? ram_447 : _GEN_6931; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6933 = 12'h1c0 == _T_6[11:0] ? ram_448 : _GEN_6932; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6934 = 12'h1c1 == _T_6[11:0] ? ram_449 : _GEN_6933; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6935 = 12'h1c2 == _T_6[11:0] ? ram_450 : _GEN_6934; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6936 = 12'h1c3 == _T_6[11:0] ? ram_451 : _GEN_6935; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6937 = 12'h1c4 == _T_6[11:0] ? ram_452 : _GEN_6936; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6938 = 12'h1c5 == _T_6[11:0] ? ram_453 : _GEN_6937; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6939 = 12'h1c6 == _T_6[11:0] ? ram_454 : _GEN_6938; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6940 = 12'h1c7 == _T_6[11:0] ? ram_455 : _GEN_6939; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6941 = 12'h1c8 == _T_6[11:0] ? ram_456 : _GEN_6940; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6942 = 12'h1c9 == _T_6[11:0] ? ram_457 : _GEN_6941; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6943 = 12'h1ca == _T_6[11:0] ? ram_458 : _GEN_6942; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6944 = 12'h1cb == _T_6[11:0] ? ram_459 : _GEN_6943; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6945 = 12'h1cc == _T_6[11:0] ? ram_460 : _GEN_6944; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6946 = 12'h1cd == _T_6[11:0] ? ram_461 : _GEN_6945; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6947 = 12'h1ce == _T_6[11:0] ? ram_462 : _GEN_6946; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6948 = 12'h1cf == _T_6[11:0] ? ram_463 : _GEN_6947; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6949 = 12'h1d0 == _T_6[11:0] ? ram_464 : _GEN_6948; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6950 = 12'h1d1 == _T_6[11:0] ? ram_465 : _GEN_6949; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6951 = 12'h1d2 == _T_6[11:0] ? ram_466 : _GEN_6950; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6952 = 12'h1d3 == _T_6[11:0] ? ram_467 : _GEN_6951; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6953 = 12'h1d4 == _T_6[11:0] ? ram_468 : _GEN_6952; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6954 = 12'h1d5 == _T_6[11:0] ? ram_469 : _GEN_6953; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6955 = 12'h1d6 == _T_6[11:0] ? ram_470 : _GEN_6954; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6956 = 12'h1d7 == _T_6[11:0] ? ram_471 : _GEN_6955; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6957 = 12'h1d8 == _T_6[11:0] ? ram_472 : _GEN_6956; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6958 = 12'h1d9 == _T_6[11:0] ? ram_473 : _GEN_6957; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6959 = 12'h1da == _T_6[11:0] ? ram_474 : _GEN_6958; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6960 = 12'h1db == _T_6[11:0] ? ram_475 : _GEN_6959; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6961 = 12'h1dc == _T_6[11:0] ? ram_476 : _GEN_6960; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6962 = 12'h1dd == _T_6[11:0] ? ram_477 : _GEN_6961; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6963 = 12'h1de == _T_6[11:0] ? ram_478 : _GEN_6962; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6964 = 12'h1df == _T_6[11:0] ? ram_479 : _GEN_6963; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6965 = 12'h1e0 == _T_6[11:0] ? ram_480 : _GEN_6964; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6966 = 12'h1e1 == _T_6[11:0] ? ram_481 : _GEN_6965; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6967 = 12'h1e2 == _T_6[11:0] ? ram_482 : _GEN_6966; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6968 = 12'h1e3 == _T_6[11:0] ? ram_483 : _GEN_6967; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6969 = 12'h1e4 == _T_6[11:0] ? ram_484 : _GEN_6968; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6970 = 12'h1e5 == _T_6[11:0] ? ram_485 : _GEN_6969; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6971 = 12'h1e6 == _T_6[11:0] ? ram_486 : _GEN_6970; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6972 = 12'h1e7 == _T_6[11:0] ? ram_487 : _GEN_6971; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6973 = 12'h1e8 == _T_6[11:0] ? ram_488 : _GEN_6972; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6974 = 12'h1e9 == _T_6[11:0] ? ram_489 : _GEN_6973; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6975 = 12'h1ea == _T_6[11:0] ? ram_490 : _GEN_6974; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6976 = 12'h1eb == _T_6[11:0] ? ram_491 : _GEN_6975; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6977 = 12'h1ec == _T_6[11:0] ? ram_492 : _GEN_6976; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6978 = 12'h1ed == _T_6[11:0] ? ram_493 : _GEN_6977; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6979 = 12'h1ee == _T_6[11:0] ? ram_494 : _GEN_6978; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6980 = 12'h1ef == _T_6[11:0] ? ram_495 : _GEN_6979; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6981 = 12'h1f0 == _T_6[11:0] ? ram_496 : _GEN_6980; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6982 = 12'h1f1 == _T_6[11:0] ? ram_497 : _GEN_6981; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6983 = 12'h1f2 == _T_6[11:0] ? ram_498 : _GEN_6982; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6984 = 12'h1f3 == _T_6[11:0] ? ram_499 : _GEN_6983; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6985 = 12'h1f4 == _T_6[11:0] ? ram_500 : _GEN_6984; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6986 = 12'h1f5 == _T_6[11:0] ? ram_501 : _GEN_6985; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6987 = 12'h1f6 == _T_6[11:0] ? ram_502 : _GEN_6986; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6988 = 12'h1f7 == _T_6[11:0] ? ram_503 : _GEN_6987; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6989 = 12'h1f8 == _T_6[11:0] ? ram_504 : _GEN_6988; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6990 = 12'h1f9 == _T_6[11:0] ? ram_505 : _GEN_6989; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6991 = 12'h1fa == _T_6[11:0] ? ram_506 : _GEN_6990; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6992 = 12'h1fb == _T_6[11:0] ? ram_507 : _GEN_6991; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6993 = 12'h1fc == _T_6[11:0] ? ram_508 : _GEN_6992; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6994 = 12'h1fd == _T_6[11:0] ? ram_509 : _GEN_6993; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6995 = 12'h1fe == _T_6[11:0] ? ram_510 : _GEN_6994; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6996 = 12'h1ff == _T_6[11:0] ? ram_511 : _GEN_6995; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6997 = 12'h200 == _T_6[11:0] ? ram_512 : _GEN_6996; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6998 = 12'h201 == _T_6[11:0] ? ram_513 : _GEN_6997; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_6999 = 12'h202 == _T_6[11:0] ? ram_514 : _GEN_6998; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7000 = 12'h203 == _T_6[11:0] ? ram_515 : _GEN_6999; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7001 = 12'h204 == _T_6[11:0] ? ram_516 : _GEN_7000; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7002 = 12'h205 == _T_6[11:0] ? ram_517 : _GEN_7001; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7003 = 12'h206 == _T_6[11:0] ? ram_518 : _GEN_7002; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7004 = 12'h207 == _T_6[11:0] ? ram_519 : _GEN_7003; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7005 = 12'h208 == _T_6[11:0] ? ram_520 : _GEN_7004; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7006 = 12'h209 == _T_6[11:0] ? ram_521 : _GEN_7005; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7007 = 12'h20a == _T_6[11:0] ? ram_522 : _GEN_7006; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7008 = 12'h20b == _T_6[11:0] ? ram_523 : _GEN_7007; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7009 = 12'h20c == _T_6[11:0] ? ram_524 : _GEN_7008; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7010 = 12'h20d == _T_6[11:0] ? ram_525 : _GEN_7009; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7011 = 12'h20e == _T_6[11:0] ? ram_526 : _GEN_7010; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7012 = 12'h20f == _T_6[11:0] ? ram_527 : _GEN_7011; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7013 = 12'h210 == _T_6[11:0] ? ram_528 : _GEN_7012; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7014 = 12'h211 == _T_6[11:0] ? ram_529 : _GEN_7013; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7015 = 12'h212 == _T_6[11:0] ? ram_530 : _GEN_7014; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7016 = 12'h213 == _T_6[11:0] ? ram_531 : _GEN_7015; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7017 = 12'h214 == _T_6[11:0] ? ram_532 : _GEN_7016; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7018 = 12'h215 == _T_6[11:0] ? ram_533 : _GEN_7017; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7019 = 12'h216 == _T_6[11:0] ? ram_534 : _GEN_7018; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7020 = 12'h217 == _T_6[11:0] ? ram_535 : _GEN_7019; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7021 = 12'h218 == _T_6[11:0] ? ram_536 : _GEN_7020; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7022 = 12'h219 == _T_6[11:0] ? ram_537 : _GEN_7021; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7023 = 12'h21a == _T_6[11:0] ? ram_538 : _GEN_7022; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7024 = 12'h21b == _T_6[11:0] ? ram_539 : _GEN_7023; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7025 = 12'h21c == _T_6[11:0] ? ram_540 : _GEN_7024; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7026 = 12'h21d == _T_6[11:0] ? ram_541 : _GEN_7025; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7027 = 12'h21e == _T_6[11:0] ? ram_542 : _GEN_7026; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7028 = 12'h21f == _T_6[11:0] ? ram_543 : _GEN_7027; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7029 = 12'h220 == _T_6[11:0] ? ram_544 : _GEN_7028; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7030 = 12'h221 == _T_6[11:0] ? ram_545 : _GEN_7029; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7031 = 12'h222 == _T_6[11:0] ? ram_546 : _GEN_7030; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7032 = 12'h223 == _T_6[11:0] ? ram_547 : _GEN_7031; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7033 = 12'h224 == _T_6[11:0] ? ram_548 : _GEN_7032; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7034 = 12'h225 == _T_6[11:0] ? ram_549 : _GEN_7033; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7035 = 12'h226 == _T_6[11:0] ? ram_550 : _GEN_7034; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7036 = 12'h227 == _T_6[11:0] ? ram_551 : _GEN_7035; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7037 = 12'h228 == _T_6[11:0] ? ram_552 : _GEN_7036; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7038 = 12'h229 == _T_6[11:0] ? ram_553 : _GEN_7037; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7039 = 12'h22a == _T_6[11:0] ? ram_554 : _GEN_7038; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7040 = 12'h22b == _T_6[11:0] ? ram_555 : _GEN_7039; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7041 = 12'h22c == _T_6[11:0] ? ram_556 : _GEN_7040; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7042 = 12'h22d == _T_6[11:0] ? ram_557 : _GEN_7041; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7043 = 12'h22e == _T_6[11:0] ? ram_558 : _GEN_7042; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7044 = 12'h22f == _T_6[11:0] ? ram_559 : _GEN_7043; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7045 = 12'h230 == _T_6[11:0] ? ram_560 : _GEN_7044; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7046 = 12'h231 == _T_6[11:0] ? ram_561 : _GEN_7045; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7047 = 12'h232 == _T_6[11:0] ? ram_562 : _GEN_7046; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7048 = 12'h233 == _T_6[11:0] ? ram_563 : _GEN_7047; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7049 = 12'h234 == _T_6[11:0] ? ram_564 : _GEN_7048; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7050 = 12'h235 == _T_6[11:0] ? ram_565 : _GEN_7049; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7051 = 12'h236 == _T_6[11:0] ? ram_566 : _GEN_7050; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7052 = 12'h237 == _T_6[11:0] ? ram_567 : _GEN_7051; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7053 = 12'h238 == _T_6[11:0] ? ram_568 : _GEN_7052; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7054 = 12'h239 == _T_6[11:0] ? ram_569 : _GEN_7053; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7055 = 12'h23a == _T_6[11:0] ? ram_570 : _GEN_7054; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7056 = 12'h23b == _T_6[11:0] ? ram_571 : _GEN_7055; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7057 = 12'h23c == _T_6[11:0] ? ram_572 : _GEN_7056; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7058 = 12'h23d == _T_6[11:0] ? ram_573 : _GEN_7057; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7059 = 12'h23e == _T_6[11:0] ? ram_574 : _GEN_7058; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7060 = 12'h23f == _T_6[11:0] ? ram_575 : _GEN_7059; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7061 = 12'h240 == _T_6[11:0] ? ram_576 : _GEN_7060; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7062 = 12'h241 == _T_6[11:0] ? ram_577 : _GEN_7061; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7063 = 12'h242 == _T_6[11:0] ? ram_578 : _GEN_7062; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7064 = 12'h243 == _T_6[11:0] ? ram_579 : _GEN_7063; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7065 = 12'h244 == _T_6[11:0] ? ram_580 : _GEN_7064; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7066 = 12'h245 == _T_6[11:0] ? ram_581 : _GEN_7065; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7067 = 12'h246 == _T_6[11:0] ? ram_582 : _GEN_7066; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7068 = 12'h247 == _T_6[11:0] ? ram_583 : _GEN_7067; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7069 = 12'h248 == _T_6[11:0] ? ram_584 : _GEN_7068; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7070 = 12'h249 == _T_6[11:0] ? ram_585 : _GEN_7069; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7071 = 12'h24a == _T_6[11:0] ? ram_586 : _GEN_7070; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7072 = 12'h24b == _T_6[11:0] ? ram_587 : _GEN_7071; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7073 = 12'h24c == _T_6[11:0] ? ram_588 : _GEN_7072; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7074 = 12'h24d == _T_6[11:0] ? ram_589 : _GEN_7073; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7075 = 12'h24e == _T_6[11:0] ? ram_590 : _GEN_7074; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7076 = 12'h24f == _T_6[11:0] ? ram_591 : _GEN_7075; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7077 = 12'h250 == _T_6[11:0] ? ram_592 : _GEN_7076; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7078 = 12'h251 == _T_6[11:0] ? ram_593 : _GEN_7077; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7079 = 12'h252 == _T_6[11:0] ? ram_594 : _GEN_7078; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7080 = 12'h253 == _T_6[11:0] ? ram_595 : _GEN_7079; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7081 = 12'h254 == _T_6[11:0] ? ram_596 : _GEN_7080; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7082 = 12'h255 == _T_6[11:0] ? ram_597 : _GEN_7081; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7083 = 12'h256 == _T_6[11:0] ? ram_598 : _GEN_7082; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7084 = 12'h257 == _T_6[11:0] ? ram_599 : _GEN_7083; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7085 = 12'h258 == _T_6[11:0] ? ram_600 : _GEN_7084; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7086 = 12'h259 == _T_6[11:0] ? ram_601 : _GEN_7085; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7087 = 12'h25a == _T_6[11:0] ? ram_602 : _GEN_7086; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7088 = 12'h25b == _T_6[11:0] ? ram_603 : _GEN_7087; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7089 = 12'h25c == _T_6[11:0] ? ram_604 : _GEN_7088; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7090 = 12'h25d == _T_6[11:0] ? ram_605 : _GEN_7089; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7091 = 12'h25e == _T_6[11:0] ? ram_606 : _GEN_7090; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7092 = 12'h25f == _T_6[11:0] ? ram_607 : _GEN_7091; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7093 = 12'h260 == _T_6[11:0] ? ram_608 : _GEN_7092; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7094 = 12'h261 == _T_6[11:0] ? ram_609 : _GEN_7093; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7095 = 12'h262 == _T_6[11:0] ? ram_610 : _GEN_7094; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7096 = 12'h263 == _T_6[11:0] ? ram_611 : _GEN_7095; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7097 = 12'h264 == _T_6[11:0] ? ram_612 : _GEN_7096; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7098 = 12'h265 == _T_6[11:0] ? ram_613 : _GEN_7097; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7099 = 12'h266 == _T_6[11:0] ? ram_614 : _GEN_7098; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7100 = 12'h267 == _T_6[11:0] ? ram_615 : _GEN_7099; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7101 = 12'h268 == _T_6[11:0] ? ram_616 : _GEN_7100; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7102 = 12'h269 == _T_6[11:0] ? ram_617 : _GEN_7101; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7103 = 12'h26a == _T_6[11:0] ? ram_618 : _GEN_7102; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7104 = 12'h26b == _T_6[11:0] ? ram_619 : _GEN_7103; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7105 = 12'h26c == _T_6[11:0] ? ram_620 : _GEN_7104; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7106 = 12'h26d == _T_6[11:0] ? ram_621 : _GEN_7105; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7107 = 12'h26e == _T_6[11:0] ? ram_622 : _GEN_7106; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7108 = 12'h26f == _T_6[11:0] ? ram_623 : _GEN_7107; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7109 = 12'h270 == _T_6[11:0] ? ram_624 : _GEN_7108; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7110 = 12'h271 == _T_6[11:0] ? ram_625 : _GEN_7109; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7111 = 12'h272 == _T_6[11:0] ? ram_626 : _GEN_7110; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7112 = 12'h273 == _T_6[11:0] ? ram_627 : _GEN_7111; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7113 = 12'h274 == _T_6[11:0] ? ram_628 : _GEN_7112; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7114 = 12'h275 == _T_6[11:0] ? ram_629 : _GEN_7113; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7115 = 12'h276 == _T_6[11:0] ? ram_630 : _GEN_7114; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7116 = 12'h277 == _T_6[11:0] ? ram_631 : _GEN_7115; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7117 = 12'h278 == _T_6[11:0] ? ram_632 : _GEN_7116; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7118 = 12'h279 == _T_6[11:0] ? ram_633 : _GEN_7117; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7119 = 12'h27a == _T_6[11:0] ? ram_634 : _GEN_7118; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7120 = 12'h27b == _T_6[11:0] ? ram_635 : _GEN_7119; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7121 = 12'h27c == _T_6[11:0] ? ram_636 : _GEN_7120; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7122 = 12'h27d == _T_6[11:0] ? ram_637 : _GEN_7121; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7123 = 12'h27e == _T_6[11:0] ? ram_638 : _GEN_7122; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7124 = 12'h27f == _T_6[11:0] ? ram_639 : _GEN_7123; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7125 = 12'h280 == _T_6[11:0] ? ram_640 : _GEN_7124; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7126 = 12'h281 == _T_6[11:0] ? ram_641 : _GEN_7125; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7127 = 12'h282 == _T_6[11:0] ? ram_642 : _GEN_7126; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7128 = 12'h283 == _T_6[11:0] ? ram_643 : _GEN_7127; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7129 = 12'h284 == _T_6[11:0] ? ram_644 : _GEN_7128; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7130 = 12'h285 == _T_6[11:0] ? ram_645 : _GEN_7129; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7131 = 12'h286 == _T_6[11:0] ? ram_646 : _GEN_7130; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7132 = 12'h287 == _T_6[11:0] ? ram_647 : _GEN_7131; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7133 = 12'h288 == _T_6[11:0] ? ram_648 : _GEN_7132; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7134 = 12'h289 == _T_6[11:0] ? ram_649 : _GEN_7133; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7135 = 12'h28a == _T_6[11:0] ? ram_650 : _GEN_7134; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7136 = 12'h28b == _T_6[11:0] ? ram_651 : _GEN_7135; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7137 = 12'h28c == _T_6[11:0] ? ram_652 : _GEN_7136; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7138 = 12'h28d == _T_6[11:0] ? ram_653 : _GEN_7137; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7139 = 12'h28e == _T_6[11:0] ? ram_654 : _GEN_7138; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7140 = 12'h28f == _T_6[11:0] ? ram_655 : _GEN_7139; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7141 = 12'h290 == _T_6[11:0] ? ram_656 : _GEN_7140; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7142 = 12'h291 == _T_6[11:0] ? ram_657 : _GEN_7141; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7143 = 12'h292 == _T_6[11:0] ? ram_658 : _GEN_7142; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7144 = 12'h293 == _T_6[11:0] ? ram_659 : _GEN_7143; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7145 = 12'h294 == _T_6[11:0] ? ram_660 : _GEN_7144; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7146 = 12'h295 == _T_6[11:0] ? ram_661 : _GEN_7145; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7147 = 12'h296 == _T_6[11:0] ? ram_662 : _GEN_7146; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7148 = 12'h297 == _T_6[11:0] ? ram_663 : _GEN_7147; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7149 = 12'h298 == _T_6[11:0] ? ram_664 : _GEN_7148; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7150 = 12'h299 == _T_6[11:0] ? ram_665 : _GEN_7149; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7151 = 12'h29a == _T_6[11:0] ? ram_666 : _GEN_7150; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7152 = 12'h29b == _T_6[11:0] ? ram_667 : _GEN_7151; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7153 = 12'h29c == _T_6[11:0] ? ram_668 : _GEN_7152; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7154 = 12'h29d == _T_6[11:0] ? ram_669 : _GEN_7153; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7155 = 12'h29e == _T_6[11:0] ? ram_670 : _GEN_7154; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7156 = 12'h29f == _T_6[11:0] ? ram_671 : _GEN_7155; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7157 = 12'h2a0 == _T_6[11:0] ? ram_672 : _GEN_7156; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7158 = 12'h2a1 == _T_6[11:0] ? ram_673 : _GEN_7157; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7159 = 12'h2a2 == _T_6[11:0] ? ram_674 : _GEN_7158; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7160 = 12'h2a3 == _T_6[11:0] ? ram_675 : _GEN_7159; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7161 = 12'h2a4 == _T_6[11:0] ? ram_676 : _GEN_7160; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7162 = 12'h2a5 == _T_6[11:0] ? ram_677 : _GEN_7161; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7163 = 12'h2a6 == _T_6[11:0] ? ram_678 : _GEN_7162; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7164 = 12'h2a7 == _T_6[11:0] ? ram_679 : _GEN_7163; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7165 = 12'h2a8 == _T_6[11:0] ? ram_680 : _GEN_7164; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7166 = 12'h2a9 == _T_6[11:0] ? ram_681 : _GEN_7165; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7167 = 12'h2aa == _T_6[11:0] ? ram_682 : _GEN_7166; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7168 = 12'h2ab == _T_6[11:0] ? ram_683 : _GEN_7167; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7169 = 12'h2ac == _T_6[11:0] ? ram_684 : _GEN_7168; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7170 = 12'h2ad == _T_6[11:0] ? ram_685 : _GEN_7169; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7171 = 12'h2ae == _T_6[11:0] ? ram_686 : _GEN_7170; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7172 = 12'h2af == _T_6[11:0] ? ram_687 : _GEN_7171; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7173 = 12'h2b0 == _T_6[11:0] ? ram_688 : _GEN_7172; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7174 = 12'h2b1 == _T_6[11:0] ? ram_689 : _GEN_7173; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7175 = 12'h2b2 == _T_6[11:0] ? ram_690 : _GEN_7174; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7176 = 12'h2b3 == _T_6[11:0] ? ram_691 : _GEN_7175; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7177 = 12'h2b4 == _T_6[11:0] ? ram_692 : _GEN_7176; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7178 = 12'h2b5 == _T_6[11:0] ? ram_693 : _GEN_7177; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7179 = 12'h2b6 == _T_6[11:0] ? ram_694 : _GEN_7178; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7180 = 12'h2b7 == _T_6[11:0] ? ram_695 : _GEN_7179; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7181 = 12'h2b8 == _T_6[11:0] ? ram_696 : _GEN_7180; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7182 = 12'h2b9 == _T_6[11:0] ? ram_697 : _GEN_7181; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7183 = 12'h2ba == _T_6[11:0] ? ram_698 : _GEN_7182; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7184 = 12'h2bb == _T_6[11:0] ? ram_699 : _GEN_7183; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7185 = 12'h2bc == _T_6[11:0] ? ram_700 : _GEN_7184; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7186 = 12'h2bd == _T_6[11:0] ? ram_701 : _GEN_7185; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7187 = 12'h2be == _T_6[11:0] ? ram_702 : _GEN_7186; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7188 = 12'h2bf == _T_6[11:0] ? ram_703 : _GEN_7187; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7189 = 12'h2c0 == _T_6[11:0] ? ram_704 : _GEN_7188; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7190 = 12'h2c1 == _T_6[11:0] ? ram_705 : _GEN_7189; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7191 = 12'h2c2 == _T_6[11:0] ? ram_706 : _GEN_7190; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7192 = 12'h2c3 == _T_6[11:0] ? ram_707 : _GEN_7191; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7193 = 12'h2c4 == _T_6[11:0] ? ram_708 : _GEN_7192; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7194 = 12'h2c5 == _T_6[11:0] ? ram_709 : _GEN_7193; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7195 = 12'h2c6 == _T_6[11:0] ? ram_710 : _GEN_7194; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7196 = 12'h2c7 == _T_6[11:0] ? ram_711 : _GEN_7195; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7197 = 12'h2c8 == _T_6[11:0] ? ram_712 : _GEN_7196; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7198 = 12'h2c9 == _T_6[11:0] ? ram_713 : _GEN_7197; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7199 = 12'h2ca == _T_6[11:0] ? ram_714 : _GEN_7198; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7200 = 12'h2cb == _T_6[11:0] ? ram_715 : _GEN_7199; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7201 = 12'h2cc == _T_6[11:0] ? ram_716 : _GEN_7200; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7202 = 12'h2cd == _T_6[11:0] ? ram_717 : _GEN_7201; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7203 = 12'h2ce == _T_6[11:0] ? ram_718 : _GEN_7202; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7204 = 12'h2cf == _T_6[11:0] ? ram_719 : _GEN_7203; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7205 = 12'h2d0 == _T_6[11:0] ? ram_720 : _GEN_7204; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7206 = 12'h2d1 == _T_6[11:0] ? ram_721 : _GEN_7205; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7207 = 12'h2d2 == _T_6[11:0] ? ram_722 : _GEN_7206; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7208 = 12'h2d3 == _T_6[11:0] ? ram_723 : _GEN_7207; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7209 = 12'h2d4 == _T_6[11:0] ? ram_724 : _GEN_7208; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7210 = 12'h2d5 == _T_6[11:0] ? ram_725 : _GEN_7209; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7211 = 12'h2d6 == _T_6[11:0] ? ram_726 : _GEN_7210; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7212 = 12'h2d7 == _T_6[11:0] ? ram_727 : _GEN_7211; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7213 = 12'h2d8 == _T_6[11:0] ? ram_728 : _GEN_7212; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7214 = 12'h2d9 == _T_6[11:0] ? ram_729 : _GEN_7213; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7215 = 12'h2da == _T_6[11:0] ? ram_730 : _GEN_7214; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7216 = 12'h2db == _T_6[11:0] ? ram_731 : _GEN_7215; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7217 = 12'h2dc == _T_6[11:0] ? ram_732 : _GEN_7216; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7218 = 12'h2dd == _T_6[11:0] ? ram_733 : _GEN_7217; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7219 = 12'h2de == _T_6[11:0] ? ram_734 : _GEN_7218; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7220 = 12'h2df == _T_6[11:0] ? ram_735 : _GEN_7219; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7221 = 12'h2e0 == _T_6[11:0] ? ram_736 : _GEN_7220; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7222 = 12'h2e1 == _T_6[11:0] ? ram_737 : _GEN_7221; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7223 = 12'h2e2 == _T_6[11:0] ? ram_738 : _GEN_7222; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7224 = 12'h2e3 == _T_6[11:0] ? ram_739 : _GEN_7223; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7225 = 12'h2e4 == _T_6[11:0] ? ram_740 : _GEN_7224; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7226 = 12'h2e5 == _T_6[11:0] ? ram_741 : _GEN_7225; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7227 = 12'h2e6 == _T_6[11:0] ? ram_742 : _GEN_7226; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7228 = 12'h2e7 == _T_6[11:0] ? ram_743 : _GEN_7227; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7229 = 12'h2e8 == _T_6[11:0] ? ram_744 : _GEN_7228; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7230 = 12'h2e9 == _T_6[11:0] ? ram_745 : _GEN_7229; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7231 = 12'h2ea == _T_6[11:0] ? ram_746 : _GEN_7230; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7232 = 12'h2eb == _T_6[11:0] ? ram_747 : _GEN_7231; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7233 = 12'h2ec == _T_6[11:0] ? ram_748 : _GEN_7232; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7234 = 12'h2ed == _T_6[11:0] ? ram_749 : _GEN_7233; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7235 = 12'h2ee == _T_6[11:0] ? ram_750 : _GEN_7234; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7236 = 12'h2ef == _T_6[11:0] ? ram_751 : _GEN_7235; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7237 = 12'h2f0 == _T_6[11:0] ? ram_752 : _GEN_7236; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7238 = 12'h2f1 == _T_6[11:0] ? ram_753 : _GEN_7237; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7239 = 12'h2f2 == _T_6[11:0] ? ram_754 : _GEN_7238; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7240 = 12'h2f3 == _T_6[11:0] ? ram_755 : _GEN_7239; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7241 = 12'h2f4 == _T_6[11:0] ? ram_756 : _GEN_7240; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7242 = 12'h2f5 == _T_6[11:0] ? ram_757 : _GEN_7241; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7243 = 12'h2f6 == _T_6[11:0] ? ram_758 : _GEN_7242; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7244 = 12'h2f7 == _T_6[11:0] ? ram_759 : _GEN_7243; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7245 = 12'h2f8 == _T_6[11:0] ? ram_760 : _GEN_7244; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7246 = 12'h2f9 == _T_6[11:0] ? ram_761 : _GEN_7245; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7247 = 12'h2fa == _T_6[11:0] ? ram_762 : _GEN_7246; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7248 = 12'h2fb == _T_6[11:0] ? ram_763 : _GEN_7247; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7249 = 12'h2fc == _T_6[11:0] ? ram_764 : _GEN_7248; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7250 = 12'h2fd == _T_6[11:0] ? ram_765 : _GEN_7249; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7251 = 12'h2fe == _T_6[11:0] ? ram_766 : _GEN_7250; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7252 = 12'h2ff == _T_6[11:0] ? ram_767 : _GEN_7251; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7253 = 12'h300 == _T_6[11:0] ? ram_768 : _GEN_7252; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7254 = 12'h301 == _T_6[11:0] ? ram_769 : _GEN_7253; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7255 = 12'h302 == _T_6[11:0] ? ram_770 : _GEN_7254; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7256 = 12'h303 == _T_6[11:0] ? ram_771 : _GEN_7255; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7257 = 12'h304 == _T_6[11:0] ? ram_772 : _GEN_7256; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7258 = 12'h305 == _T_6[11:0] ? ram_773 : _GEN_7257; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7259 = 12'h306 == _T_6[11:0] ? ram_774 : _GEN_7258; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7260 = 12'h307 == _T_6[11:0] ? ram_775 : _GEN_7259; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7261 = 12'h308 == _T_6[11:0] ? ram_776 : _GEN_7260; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7262 = 12'h309 == _T_6[11:0] ? ram_777 : _GEN_7261; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7263 = 12'h30a == _T_6[11:0] ? ram_778 : _GEN_7262; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7264 = 12'h30b == _T_6[11:0] ? ram_779 : _GEN_7263; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7265 = 12'h30c == _T_6[11:0] ? ram_780 : _GEN_7264; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7266 = 12'h30d == _T_6[11:0] ? ram_781 : _GEN_7265; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7267 = 12'h30e == _T_6[11:0] ? ram_782 : _GEN_7266; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7268 = 12'h30f == _T_6[11:0] ? ram_783 : _GEN_7267; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7269 = 12'h310 == _T_6[11:0] ? ram_784 : _GEN_7268; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7270 = 12'h311 == _T_6[11:0] ? ram_785 : _GEN_7269; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7271 = 12'h312 == _T_6[11:0] ? ram_786 : _GEN_7270; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7272 = 12'h313 == _T_6[11:0] ? ram_787 : _GEN_7271; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7273 = 12'h314 == _T_6[11:0] ? ram_788 : _GEN_7272; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7274 = 12'h315 == _T_6[11:0] ? ram_789 : _GEN_7273; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7275 = 12'h316 == _T_6[11:0] ? ram_790 : _GEN_7274; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7276 = 12'h317 == _T_6[11:0] ? ram_791 : _GEN_7275; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7277 = 12'h318 == _T_6[11:0] ? ram_792 : _GEN_7276; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7278 = 12'h319 == _T_6[11:0] ? ram_793 : _GEN_7277; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7279 = 12'h31a == _T_6[11:0] ? ram_794 : _GEN_7278; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7280 = 12'h31b == _T_6[11:0] ? ram_795 : _GEN_7279; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7281 = 12'h31c == _T_6[11:0] ? ram_796 : _GEN_7280; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7282 = 12'h31d == _T_6[11:0] ? ram_797 : _GEN_7281; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7283 = 12'h31e == _T_6[11:0] ? ram_798 : _GEN_7282; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7284 = 12'h31f == _T_6[11:0] ? ram_799 : _GEN_7283; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7285 = 12'h320 == _T_6[11:0] ? ram_800 : _GEN_7284; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7286 = 12'h321 == _T_6[11:0] ? ram_801 : _GEN_7285; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7287 = 12'h322 == _T_6[11:0] ? ram_802 : _GEN_7286; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7288 = 12'h323 == _T_6[11:0] ? ram_803 : _GEN_7287; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7289 = 12'h324 == _T_6[11:0] ? ram_804 : _GEN_7288; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7290 = 12'h325 == _T_6[11:0] ? ram_805 : _GEN_7289; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7291 = 12'h326 == _T_6[11:0] ? ram_806 : _GEN_7290; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7292 = 12'h327 == _T_6[11:0] ? ram_807 : _GEN_7291; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7293 = 12'h328 == _T_6[11:0] ? ram_808 : _GEN_7292; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7294 = 12'h329 == _T_6[11:0] ? ram_809 : _GEN_7293; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7295 = 12'h32a == _T_6[11:0] ? ram_810 : _GEN_7294; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7296 = 12'h32b == _T_6[11:0] ? ram_811 : _GEN_7295; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7297 = 12'h32c == _T_6[11:0] ? ram_812 : _GEN_7296; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7298 = 12'h32d == _T_6[11:0] ? ram_813 : _GEN_7297; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7299 = 12'h32e == _T_6[11:0] ? ram_814 : _GEN_7298; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7300 = 12'h32f == _T_6[11:0] ? ram_815 : _GEN_7299; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7301 = 12'h330 == _T_6[11:0] ? ram_816 : _GEN_7300; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7302 = 12'h331 == _T_6[11:0] ? ram_817 : _GEN_7301; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7303 = 12'h332 == _T_6[11:0] ? ram_818 : _GEN_7302; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7304 = 12'h333 == _T_6[11:0] ? ram_819 : _GEN_7303; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7305 = 12'h334 == _T_6[11:0] ? ram_820 : _GEN_7304; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7306 = 12'h335 == _T_6[11:0] ? ram_821 : _GEN_7305; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7307 = 12'h336 == _T_6[11:0] ? ram_822 : _GEN_7306; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7308 = 12'h337 == _T_6[11:0] ? ram_823 : _GEN_7307; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7309 = 12'h338 == _T_6[11:0] ? ram_824 : _GEN_7308; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7310 = 12'h339 == _T_6[11:0] ? ram_825 : _GEN_7309; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7311 = 12'h33a == _T_6[11:0] ? ram_826 : _GEN_7310; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7312 = 12'h33b == _T_6[11:0] ? ram_827 : _GEN_7311; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7313 = 12'h33c == _T_6[11:0] ? ram_828 : _GEN_7312; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7314 = 12'h33d == _T_6[11:0] ? ram_829 : _GEN_7313; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7315 = 12'h33e == _T_6[11:0] ? ram_830 : _GEN_7314; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7316 = 12'h33f == _T_6[11:0] ? ram_831 : _GEN_7315; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7317 = 12'h340 == _T_6[11:0] ? ram_832 : _GEN_7316; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7318 = 12'h341 == _T_6[11:0] ? ram_833 : _GEN_7317; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7319 = 12'h342 == _T_6[11:0] ? ram_834 : _GEN_7318; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7320 = 12'h343 == _T_6[11:0] ? ram_835 : _GEN_7319; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7321 = 12'h344 == _T_6[11:0] ? ram_836 : _GEN_7320; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7322 = 12'h345 == _T_6[11:0] ? ram_837 : _GEN_7321; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7323 = 12'h346 == _T_6[11:0] ? ram_838 : _GEN_7322; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7324 = 12'h347 == _T_6[11:0] ? ram_839 : _GEN_7323; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7325 = 12'h348 == _T_6[11:0] ? ram_840 : _GEN_7324; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7326 = 12'h349 == _T_6[11:0] ? ram_841 : _GEN_7325; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7327 = 12'h34a == _T_6[11:0] ? ram_842 : _GEN_7326; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7328 = 12'h34b == _T_6[11:0] ? ram_843 : _GEN_7327; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7329 = 12'h34c == _T_6[11:0] ? ram_844 : _GEN_7328; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7330 = 12'h34d == _T_6[11:0] ? ram_845 : _GEN_7329; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7331 = 12'h34e == _T_6[11:0] ? ram_846 : _GEN_7330; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7332 = 12'h34f == _T_6[11:0] ? ram_847 : _GEN_7331; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7333 = 12'h350 == _T_6[11:0] ? ram_848 : _GEN_7332; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7334 = 12'h351 == _T_6[11:0] ? ram_849 : _GEN_7333; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7335 = 12'h352 == _T_6[11:0] ? ram_850 : _GEN_7334; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7336 = 12'h353 == _T_6[11:0] ? ram_851 : _GEN_7335; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7337 = 12'h354 == _T_6[11:0] ? ram_852 : _GEN_7336; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7338 = 12'h355 == _T_6[11:0] ? ram_853 : _GEN_7337; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7339 = 12'h356 == _T_6[11:0] ? ram_854 : _GEN_7338; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7340 = 12'h357 == _T_6[11:0] ? ram_855 : _GEN_7339; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7341 = 12'h358 == _T_6[11:0] ? ram_856 : _GEN_7340; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7342 = 12'h359 == _T_6[11:0] ? ram_857 : _GEN_7341; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7343 = 12'h35a == _T_6[11:0] ? ram_858 : _GEN_7342; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7344 = 12'h35b == _T_6[11:0] ? ram_859 : _GEN_7343; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7345 = 12'h35c == _T_6[11:0] ? ram_860 : _GEN_7344; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7346 = 12'h35d == _T_6[11:0] ? ram_861 : _GEN_7345; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7347 = 12'h35e == _T_6[11:0] ? ram_862 : _GEN_7346; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7348 = 12'h35f == _T_6[11:0] ? ram_863 : _GEN_7347; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7349 = 12'h360 == _T_6[11:0] ? ram_864 : _GEN_7348; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7350 = 12'h361 == _T_6[11:0] ? ram_865 : _GEN_7349; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7351 = 12'h362 == _T_6[11:0] ? ram_866 : _GEN_7350; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7352 = 12'h363 == _T_6[11:0] ? ram_867 : _GEN_7351; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7353 = 12'h364 == _T_6[11:0] ? ram_868 : _GEN_7352; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7354 = 12'h365 == _T_6[11:0] ? ram_869 : _GEN_7353; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7355 = 12'h366 == _T_6[11:0] ? ram_870 : _GEN_7354; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7356 = 12'h367 == _T_6[11:0] ? ram_871 : _GEN_7355; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7357 = 12'h368 == _T_6[11:0] ? ram_872 : _GEN_7356; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7358 = 12'h369 == _T_6[11:0] ? ram_873 : _GEN_7357; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7359 = 12'h36a == _T_6[11:0] ? ram_874 : _GEN_7358; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7360 = 12'h36b == _T_6[11:0] ? ram_875 : _GEN_7359; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7361 = 12'h36c == _T_6[11:0] ? ram_876 : _GEN_7360; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7362 = 12'h36d == _T_6[11:0] ? ram_877 : _GEN_7361; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7363 = 12'h36e == _T_6[11:0] ? ram_878 : _GEN_7362; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7364 = 12'h36f == _T_6[11:0] ? ram_879 : _GEN_7363; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7365 = 12'h370 == _T_6[11:0] ? ram_880 : _GEN_7364; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7366 = 12'h371 == _T_6[11:0] ? ram_881 : _GEN_7365; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7367 = 12'h372 == _T_6[11:0] ? ram_882 : _GEN_7366; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7368 = 12'h373 == _T_6[11:0] ? ram_883 : _GEN_7367; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7369 = 12'h374 == _T_6[11:0] ? ram_884 : _GEN_7368; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7370 = 12'h375 == _T_6[11:0] ? ram_885 : _GEN_7369; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7371 = 12'h376 == _T_6[11:0] ? ram_886 : _GEN_7370; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7372 = 12'h377 == _T_6[11:0] ? ram_887 : _GEN_7371; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7373 = 12'h378 == _T_6[11:0] ? ram_888 : _GEN_7372; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7374 = 12'h379 == _T_6[11:0] ? ram_889 : _GEN_7373; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7375 = 12'h37a == _T_6[11:0] ? ram_890 : _GEN_7374; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7376 = 12'h37b == _T_6[11:0] ? ram_891 : _GEN_7375; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7377 = 12'h37c == _T_6[11:0] ? ram_892 : _GEN_7376; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7378 = 12'h37d == _T_6[11:0] ? ram_893 : _GEN_7377; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7379 = 12'h37e == _T_6[11:0] ? ram_894 : _GEN_7378; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7380 = 12'h37f == _T_6[11:0] ? ram_895 : _GEN_7379; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7381 = 12'h380 == _T_6[11:0] ? ram_896 : _GEN_7380; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7382 = 12'h381 == _T_6[11:0] ? ram_897 : _GEN_7381; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7383 = 12'h382 == _T_6[11:0] ? ram_898 : _GEN_7382; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7384 = 12'h383 == _T_6[11:0] ? ram_899 : _GEN_7383; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7385 = 12'h384 == _T_6[11:0] ? ram_900 : _GEN_7384; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7386 = 12'h385 == _T_6[11:0] ? ram_901 : _GEN_7385; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7387 = 12'h386 == _T_6[11:0] ? ram_902 : _GEN_7386; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7388 = 12'h387 == _T_6[11:0] ? ram_903 : _GEN_7387; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7389 = 12'h388 == _T_6[11:0] ? ram_904 : _GEN_7388; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7390 = 12'h389 == _T_6[11:0] ? ram_905 : _GEN_7389; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7391 = 12'h38a == _T_6[11:0] ? ram_906 : _GEN_7390; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7392 = 12'h38b == _T_6[11:0] ? ram_907 : _GEN_7391; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7393 = 12'h38c == _T_6[11:0] ? ram_908 : _GEN_7392; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7394 = 12'h38d == _T_6[11:0] ? ram_909 : _GEN_7393; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7395 = 12'h38e == _T_6[11:0] ? ram_910 : _GEN_7394; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7396 = 12'h38f == _T_6[11:0] ? ram_911 : _GEN_7395; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7397 = 12'h390 == _T_6[11:0] ? ram_912 : _GEN_7396; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7398 = 12'h391 == _T_6[11:0] ? ram_913 : _GEN_7397; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7399 = 12'h392 == _T_6[11:0] ? ram_914 : _GEN_7398; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7400 = 12'h393 == _T_6[11:0] ? ram_915 : _GEN_7399; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7401 = 12'h394 == _T_6[11:0] ? ram_916 : _GEN_7400; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7402 = 12'h395 == _T_6[11:0] ? ram_917 : _GEN_7401; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7403 = 12'h396 == _T_6[11:0] ? ram_918 : _GEN_7402; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7404 = 12'h397 == _T_6[11:0] ? ram_919 : _GEN_7403; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7405 = 12'h398 == _T_6[11:0] ? ram_920 : _GEN_7404; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7406 = 12'h399 == _T_6[11:0] ? ram_921 : _GEN_7405; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7407 = 12'h39a == _T_6[11:0] ? ram_922 : _GEN_7406; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7408 = 12'h39b == _T_6[11:0] ? ram_923 : _GEN_7407; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7409 = 12'h39c == _T_6[11:0] ? ram_924 : _GEN_7408; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7410 = 12'h39d == _T_6[11:0] ? ram_925 : _GEN_7409; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7411 = 12'h39e == _T_6[11:0] ? ram_926 : _GEN_7410; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7412 = 12'h39f == _T_6[11:0] ? ram_927 : _GEN_7411; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7413 = 12'h3a0 == _T_6[11:0] ? ram_928 : _GEN_7412; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7414 = 12'h3a1 == _T_6[11:0] ? ram_929 : _GEN_7413; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7415 = 12'h3a2 == _T_6[11:0] ? ram_930 : _GEN_7414; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7416 = 12'h3a3 == _T_6[11:0] ? ram_931 : _GEN_7415; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7417 = 12'h3a4 == _T_6[11:0] ? ram_932 : _GEN_7416; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7418 = 12'h3a5 == _T_6[11:0] ? ram_933 : _GEN_7417; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7419 = 12'h3a6 == _T_6[11:0] ? ram_934 : _GEN_7418; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7420 = 12'h3a7 == _T_6[11:0] ? ram_935 : _GEN_7419; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7421 = 12'h3a8 == _T_6[11:0] ? ram_936 : _GEN_7420; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7422 = 12'h3a9 == _T_6[11:0] ? ram_937 : _GEN_7421; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7423 = 12'h3aa == _T_6[11:0] ? ram_938 : _GEN_7422; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7424 = 12'h3ab == _T_6[11:0] ? ram_939 : _GEN_7423; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7425 = 12'h3ac == _T_6[11:0] ? ram_940 : _GEN_7424; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7426 = 12'h3ad == _T_6[11:0] ? ram_941 : _GEN_7425; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7427 = 12'h3ae == _T_6[11:0] ? ram_942 : _GEN_7426; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7428 = 12'h3af == _T_6[11:0] ? ram_943 : _GEN_7427; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7429 = 12'h3b0 == _T_6[11:0] ? ram_944 : _GEN_7428; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7430 = 12'h3b1 == _T_6[11:0] ? ram_945 : _GEN_7429; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7431 = 12'h3b2 == _T_6[11:0] ? ram_946 : _GEN_7430; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7432 = 12'h3b3 == _T_6[11:0] ? ram_947 : _GEN_7431; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7433 = 12'h3b4 == _T_6[11:0] ? ram_948 : _GEN_7432; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7434 = 12'h3b5 == _T_6[11:0] ? ram_949 : _GEN_7433; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7435 = 12'h3b6 == _T_6[11:0] ? ram_950 : _GEN_7434; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7436 = 12'h3b7 == _T_6[11:0] ? ram_951 : _GEN_7435; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7437 = 12'h3b8 == _T_6[11:0] ? ram_952 : _GEN_7436; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7438 = 12'h3b9 == _T_6[11:0] ? ram_953 : _GEN_7437; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7439 = 12'h3ba == _T_6[11:0] ? ram_954 : _GEN_7438; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7440 = 12'h3bb == _T_6[11:0] ? ram_955 : _GEN_7439; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7441 = 12'h3bc == _T_6[11:0] ? ram_956 : _GEN_7440; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7442 = 12'h3bd == _T_6[11:0] ? ram_957 : _GEN_7441; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7443 = 12'h3be == _T_6[11:0] ? ram_958 : _GEN_7442; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7444 = 12'h3bf == _T_6[11:0] ? ram_959 : _GEN_7443; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7445 = 12'h3c0 == _T_6[11:0] ? ram_960 : _GEN_7444; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7446 = 12'h3c1 == _T_6[11:0] ? ram_961 : _GEN_7445; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7447 = 12'h3c2 == _T_6[11:0] ? ram_962 : _GEN_7446; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7448 = 12'h3c3 == _T_6[11:0] ? ram_963 : _GEN_7447; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7449 = 12'h3c4 == _T_6[11:0] ? ram_964 : _GEN_7448; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7450 = 12'h3c5 == _T_6[11:0] ? ram_965 : _GEN_7449; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7451 = 12'h3c6 == _T_6[11:0] ? ram_966 : _GEN_7450; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7452 = 12'h3c7 == _T_6[11:0] ? ram_967 : _GEN_7451; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7453 = 12'h3c8 == _T_6[11:0] ? ram_968 : _GEN_7452; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7454 = 12'h3c9 == _T_6[11:0] ? ram_969 : _GEN_7453; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7455 = 12'h3ca == _T_6[11:0] ? ram_970 : _GEN_7454; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7456 = 12'h3cb == _T_6[11:0] ? ram_971 : _GEN_7455; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7457 = 12'h3cc == _T_6[11:0] ? ram_972 : _GEN_7456; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7458 = 12'h3cd == _T_6[11:0] ? ram_973 : _GEN_7457; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7459 = 12'h3ce == _T_6[11:0] ? ram_974 : _GEN_7458; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7460 = 12'h3cf == _T_6[11:0] ? ram_975 : _GEN_7459; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7461 = 12'h3d0 == _T_6[11:0] ? ram_976 : _GEN_7460; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7462 = 12'h3d1 == _T_6[11:0] ? ram_977 : _GEN_7461; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7463 = 12'h3d2 == _T_6[11:0] ? ram_978 : _GEN_7462; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7464 = 12'h3d3 == _T_6[11:0] ? ram_979 : _GEN_7463; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7465 = 12'h3d4 == _T_6[11:0] ? ram_980 : _GEN_7464; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7466 = 12'h3d5 == _T_6[11:0] ? ram_981 : _GEN_7465; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7467 = 12'h3d6 == _T_6[11:0] ? ram_982 : _GEN_7466; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7468 = 12'h3d7 == _T_6[11:0] ? ram_983 : _GEN_7467; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7469 = 12'h3d8 == _T_6[11:0] ? ram_984 : _GEN_7468; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7470 = 12'h3d9 == _T_6[11:0] ? ram_985 : _GEN_7469; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7471 = 12'h3da == _T_6[11:0] ? ram_986 : _GEN_7470; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7472 = 12'h3db == _T_6[11:0] ? ram_987 : _GEN_7471; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7473 = 12'h3dc == _T_6[11:0] ? ram_988 : _GEN_7472; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7474 = 12'h3dd == _T_6[11:0] ? ram_989 : _GEN_7473; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7475 = 12'h3de == _T_6[11:0] ? ram_990 : _GEN_7474; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7476 = 12'h3df == _T_6[11:0] ? ram_991 : _GEN_7475; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7477 = 12'h3e0 == _T_6[11:0] ? ram_992 : _GEN_7476; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7478 = 12'h3e1 == _T_6[11:0] ? ram_993 : _GEN_7477; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7479 = 12'h3e2 == _T_6[11:0] ? ram_994 : _GEN_7478; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7480 = 12'h3e3 == _T_6[11:0] ? ram_995 : _GEN_7479; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7481 = 12'h3e4 == _T_6[11:0] ? ram_996 : _GEN_7480; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7482 = 12'h3e5 == _T_6[11:0] ? ram_997 : _GEN_7481; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7483 = 12'h3e6 == _T_6[11:0] ? ram_998 : _GEN_7482; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7484 = 12'h3e7 == _T_6[11:0] ? ram_999 : _GEN_7483; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7485 = 12'h3e8 == _T_6[11:0] ? ram_1000 : _GEN_7484; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7486 = 12'h3e9 == _T_6[11:0] ? ram_1001 : _GEN_7485; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7487 = 12'h3ea == _T_6[11:0] ? ram_1002 : _GEN_7486; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7488 = 12'h3eb == _T_6[11:0] ? ram_1003 : _GEN_7487; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7489 = 12'h3ec == _T_6[11:0] ? ram_1004 : _GEN_7488; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7490 = 12'h3ed == _T_6[11:0] ? ram_1005 : _GEN_7489; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7491 = 12'h3ee == _T_6[11:0] ? ram_1006 : _GEN_7490; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7492 = 12'h3ef == _T_6[11:0] ? ram_1007 : _GEN_7491; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7493 = 12'h3f0 == _T_6[11:0] ? ram_1008 : _GEN_7492; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7494 = 12'h3f1 == _T_6[11:0] ? ram_1009 : _GEN_7493; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7495 = 12'h3f2 == _T_6[11:0] ? ram_1010 : _GEN_7494; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7496 = 12'h3f3 == _T_6[11:0] ? ram_1011 : _GEN_7495; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7497 = 12'h3f4 == _T_6[11:0] ? ram_1012 : _GEN_7496; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7498 = 12'h3f5 == _T_6[11:0] ? ram_1013 : _GEN_7497; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7499 = 12'h3f6 == _T_6[11:0] ? ram_1014 : _GEN_7498; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7500 = 12'h3f7 == _T_6[11:0] ? ram_1015 : _GEN_7499; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7501 = 12'h3f8 == _T_6[11:0] ? ram_1016 : _GEN_7500; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7502 = 12'h3f9 == _T_6[11:0] ? ram_1017 : _GEN_7501; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7503 = 12'h3fa == _T_6[11:0] ? ram_1018 : _GEN_7502; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7504 = 12'h3fb == _T_6[11:0] ? ram_1019 : _GEN_7503; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7505 = 12'h3fc == _T_6[11:0] ? ram_1020 : _GEN_7504; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7506 = 12'h3fd == _T_6[11:0] ? ram_1021 : _GEN_7505; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7507 = 12'h3fe == _T_6[11:0] ? ram_1022 : _GEN_7506; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7508 = 12'h3ff == _T_6[11:0] ? ram_1023 : _GEN_7507; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7509 = 12'h400 == _T_6[11:0] ? ram_1024 : _GEN_7508; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7510 = 12'h401 == _T_6[11:0] ? ram_1025 : _GEN_7509; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7511 = 12'h402 == _T_6[11:0] ? ram_1026 : _GEN_7510; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7512 = 12'h403 == _T_6[11:0] ? ram_1027 : _GEN_7511; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7513 = 12'h404 == _T_6[11:0] ? ram_1028 : _GEN_7512; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7514 = 12'h405 == _T_6[11:0] ? ram_1029 : _GEN_7513; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7515 = 12'h406 == _T_6[11:0] ? ram_1030 : _GEN_7514; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7516 = 12'h407 == _T_6[11:0] ? ram_1031 : _GEN_7515; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7517 = 12'h408 == _T_6[11:0] ? ram_1032 : _GEN_7516; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7518 = 12'h409 == _T_6[11:0] ? ram_1033 : _GEN_7517; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7519 = 12'h40a == _T_6[11:0] ? ram_1034 : _GEN_7518; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7520 = 12'h40b == _T_6[11:0] ? ram_1035 : _GEN_7519; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7521 = 12'h40c == _T_6[11:0] ? ram_1036 : _GEN_7520; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7522 = 12'h40d == _T_6[11:0] ? ram_1037 : _GEN_7521; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7523 = 12'h40e == _T_6[11:0] ? ram_1038 : _GEN_7522; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7524 = 12'h40f == _T_6[11:0] ? ram_1039 : _GEN_7523; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7525 = 12'h410 == _T_6[11:0] ? ram_1040 : _GEN_7524; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7526 = 12'h411 == _T_6[11:0] ? ram_1041 : _GEN_7525; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7527 = 12'h412 == _T_6[11:0] ? ram_1042 : _GEN_7526; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7528 = 12'h413 == _T_6[11:0] ? ram_1043 : _GEN_7527; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7529 = 12'h414 == _T_6[11:0] ? ram_1044 : _GEN_7528; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7530 = 12'h415 == _T_6[11:0] ? ram_1045 : _GEN_7529; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7531 = 12'h416 == _T_6[11:0] ? ram_1046 : _GEN_7530; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7532 = 12'h417 == _T_6[11:0] ? ram_1047 : _GEN_7531; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7533 = 12'h418 == _T_6[11:0] ? ram_1048 : _GEN_7532; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7534 = 12'h419 == _T_6[11:0] ? ram_1049 : _GEN_7533; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7535 = 12'h41a == _T_6[11:0] ? ram_1050 : _GEN_7534; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7536 = 12'h41b == _T_6[11:0] ? ram_1051 : _GEN_7535; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7537 = 12'h41c == _T_6[11:0] ? ram_1052 : _GEN_7536; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7538 = 12'h41d == _T_6[11:0] ? ram_1053 : _GEN_7537; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7539 = 12'h41e == _T_6[11:0] ? ram_1054 : _GEN_7538; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7540 = 12'h41f == _T_6[11:0] ? ram_1055 : _GEN_7539; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7541 = 12'h420 == _T_6[11:0] ? ram_1056 : _GEN_7540; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7542 = 12'h421 == _T_6[11:0] ? ram_1057 : _GEN_7541; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7543 = 12'h422 == _T_6[11:0] ? ram_1058 : _GEN_7542; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7544 = 12'h423 == _T_6[11:0] ? ram_1059 : _GEN_7543; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7545 = 12'h424 == _T_6[11:0] ? ram_1060 : _GEN_7544; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7546 = 12'h425 == _T_6[11:0] ? ram_1061 : _GEN_7545; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7547 = 12'h426 == _T_6[11:0] ? ram_1062 : _GEN_7546; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7548 = 12'h427 == _T_6[11:0] ? ram_1063 : _GEN_7547; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7549 = 12'h428 == _T_6[11:0] ? ram_1064 : _GEN_7548; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7550 = 12'h429 == _T_6[11:0] ? ram_1065 : _GEN_7549; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7551 = 12'h42a == _T_6[11:0] ? ram_1066 : _GEN_7550; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7552 = 12'h42b == _T_6[11:0] ? ram_1067 : _GEN_7551; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7553 = 12'h42c == _T_6[11:0] ? ram_1068 : _GEN_7552; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7554 = 12'h42d == _T_6[11:0] ? ram_1069 : _GEN_7553; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7555 = 12'h42e == _T_6[11:0] ? ram_1070 : _GEN_7554; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7556 = 12'h42f == _T_6[11:0] ? ram_1071 : _GEN_7555; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7557 = 12'h430 == _T_6[11:0] ? ram_1072 : _GEN_7556; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7558 = 12'h431 == _T_6[11:0] ? ram_1073 : _GEN_7557; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7559 = 12'h432 == _T_6[11:0] ? ram_1074 : _GEN_7558; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7560 = 12'h433 == _T_6[11:0] ? ram_1075 : _GEN_7559; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7561 = 12'h434 == _T_6[11:0] ? ram_1076 : _GEN_7560; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7562 = 12'h435 == _T_6[11:0] ? ram_1077 : _GEN_7561; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7563 = 12'h436 == _T_6[11:0] ? ram_1078 : _GEN_7562; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7564 = 12'h437 == _T_6[11:0] ? ram_1079 : _GEN_7563; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7565 = 12'h438 == _T_6[11:0] ? ram_1080 : _GEN_7564; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7566 = 12'h439 == _T_6[11:0] ? ram_1081 : _GEN_7565; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7567 = 12'h43a == _T_6[11:0] ? ram_1082 : _GEN_7566; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7568 = 12'h43b == _T_6[11:0] ? ram_1083 : _GEN_7567; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7569 = 12'h43c == _T_6[11:0] ? ram_1084 : _GEN_7568; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7570 = 12'h43d == _T_6[11:0] ? ram_1085 : _GEN_7569; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7571 = 12'h43e == _T_6[11:0] ? ram_1086 : _GEN_7570; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7572 = 12'h43f == _T_6[11:0] ? ram_1087 : _GEN_7571; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7573 = 12'h440 == _T_6[11:0] ? ram_1088 : _GEN_7572; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7574 = 12'h441 == _T_6[11:0] ? ram_1089 : _GEN_7573; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7575 = 12'h442 == _T_6[11:0] ? ram_1090 : _GEN_7574; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7576 = 12'h443 == _T_6[11:0] ? ram_1091 : _GEN_7575; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7577 = 12'h444 == _T_6[11:0] ? ram_1092 : _GEN_7576; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7578 = 12'h445 == _T_6[11:0] ? ram_1093 : _GEN_7577; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7579 = 12'h446 == _T_6[11:0] ? ram_1094 : _GEN_7578; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7580 = 12'h447 == _T_6[11:0] ? ram_1095 : _GEN_7579; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7581 = 12'h448 == _T_6[11:0] ? ram_1096 : _GEN_7580; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7582 = 12'h449 == _T_6[11:0] ? ram_1097 : _GEN_7581; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7583 = 12'h44a == _T_6[11:0] ? ram_1098 : _GEN_7582; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7584 = 12'h44b == _T_6[11:0] ? ram_1099 : _GEN_7583; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7585 = 12'h44c == _T_6[11:0] ? ram_1100 : _GEN_7584; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7586 = 12'h44d == _T_6[11:0] ? ram_1101 : _GEN_7585; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7587 = 12'h44e == _T_6[11:0] ? ram_1102 : _GEN_7586; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7588 = 12'h44f == _T_6[11:0] ? ram_1103 : _GEN_7587; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7589 = 12'h450 == _T_6[11:0] ? ram_1104 : _GEN_7588; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7590 = 12'h451 == _T_6[11:0] ? ram_1105 : _GEN_7589; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7591 = 12'h452 == _T_6[11:0] ? ram_1106 : _GEN_7590; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7592 = 12'h453 == _T_6[11:0] ? ram_1107 : _GEN_7591; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7593 = 12'h454 == _T_6[11:0] ? ram_1108 : _GEN_7592; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7594 = 12'h455 == _T_6[11:0] ? ram_1109 : _GEN_7593; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7595 = 12'h456 == _T_6[11:0] ? ram_1110 : _GEN_7594; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7596 = 12'h457 == _T_6[11:0] ? ram_1111 : _GEN_7595; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7597 = 12'h458 == _T_6[11:0] ? ram_1112 : _GEN_7596; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7598 = 12'h459 == _T_6[11:0] ? ram_1113 : _GEN_7597; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7599 = 12'h45a == _T_6[11:0] ? ram_1114 : _GEN_7598; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7600 = 12'h45b == _T_6[11:0] ? ram_1115 : _GEN_7599; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7601 = 12'h45c == _T_6[11:0] ? ram_1116 : _GEN_7600; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7602 = 12'h45d == _T_6[11:0] ? ram_1117 : _GEN_7601; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7603 = 12'h45e == _T_6[11:0] ? ram_1118 : _GEN_7602; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7604 = 12'h45f == _T_6[11:0] ? ram_1119 : _GEN_7603; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7605 = 12'h460 == _T_6[11:0] ? ram_1120 : _GEN_7604; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7606 = 12'h461 == _T_6[11:0] ? ram_1121 : _GEN_7605; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7607 = 12'h462 == _T_6[11:0] ? ram_1122 : _GEN_7606; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7608 = 12'h463 == _T_6[11:0] ? ram_1123 : _GEN_7607; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7609 = 12'h464 == _T_6[11:0] ? ram_1124 : _GEN_7608; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7610 = 12'h465 == _T_6[11:0] ? ram_1125 : _GEN_7609; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7611 = 12'h466 == _T_6[11:0] ? ram_1126 : _GEN_7610; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7612 = 12'h467 == _T_6[11:0] ? ram_1127 : _GEN_7611; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7613 = 12'h468 == _T_6[11:0] ? ram_1128 : _GEN_7612; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7614 = 12'h469 == _T_6[11:0] ? ram_1129 : _GEN_7613; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7615 = 12'h46a == _T_6[11:0] ? ram_1130 : _GEN_7614; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7616 = 12'h46b == _T_6[11:0] ? ram_1131 : _GEN_7615; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7617 = 12'h46c == _T_6[11:0] ? ram_1132 : _GEN_7616; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7618 = 12'h46d == _T_6[11:0] ? ram_1133 : _GEN_7617; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7619 = 12'h46e == _T_6[11:0] ? ram_1134 : _GEN_7618; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7620 = 12'h46f == _T_6[11:0] ? ram_1135 : _GEN_7619; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7621 = 12'h470 == _T_6[11:0] ? ram_1136 : _GEN_7620; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7622 = 12'h471 == _T_6[11:0] ? ram_1137 : _GEN_7621; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7623 = 12'h472 == _T_6[11:0] ? ram_1138 : _GEN_7622; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7624 = 12'h473 == _T_6[11:0] ? ram_1139 : _GEN_7623; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7625 = 12'h474 == _T_6[11:0] ? ram_1140 : _GEN_7624; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7626 = 12'h475 == _T_6[11:0] ? ram_1141 : _GEN_7625; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7627 = 12'h476 == _T_6[11:0] ? ram_1142 : _GEN_7626; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7628 = 12'h477 == _T_6[11:0] ? ram_1143 : _GEN_7627; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7629 = 12'h478 == _T_6[11:0] ? ram_1144 : _GEN_7628; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7630 = 12'h479 == _T_6[11:0] ? ram_1145 : _GEN_7629; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7631 = 12'h47a == _T_6[11:0] ? ram_1146 : _GEN_7630; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7632 = 12'h47b == _T_6[11:0] ? ram_1147 : _GEN_7631; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7633 = 12'h47c == _T_6[11:0] ? ram_1148 : _GEN_7632; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7634 = 12'h47d == _T_6[11:0] ? ram_1149 : _GEN_7633; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7635 = 12'h47e == _T_6[11:0] ? ram_1150 : _GEN_7634; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7636 = 12'h47f == _T_6[11:0] ? ram_1151 : _GEN_7635; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7637 = 12'h480 == _T_6[11:0] ? ram_1152 : _GEN_7636; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7638 = 12'h481 == _T_6[11:0] ? ram_1153 : _GEN_7637; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7639 = 12'h482 == _T_6[11:0] ? ram_1154 : _GEN_7638; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7640 = 12'h483 == _T_6[11:0] ? ram_1155 : _GEN_7639; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7641 = 12'h484 == _T_6[11:0] ? ram_1156 : _GEN_7640; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7642 = 12'h485 == _T_6[11:0] ? ram_1157 : _GEN_7641; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7643 = 12'h486 == _T_6[11:0] ? ram_1158 : _GEN_7642; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7644 = 12'h487 == _T_6[11:0] ? ram_1159 : _GEN_7643; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7645 = 12'h488 == _T_6[11:0] ? ram_1160 : _GEN_7644; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7646 = 12'h489 == _T_6[11:0] ? ram_1161 : _GEN_7645; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7647 = 12'h48a == _T_6[11:0] ? ram_1162 : _GEN_7646; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7648 = 12'h48b == _T_6[11:0] ? ram_1163 : _GEN_7647; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7649 = 12'h48c == _T_6[11:0] ? ram_1164 : _GEN_7648; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7650 = 12'h48d == _T_6[11:0] ? ram_1165 : _GEN_7649; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7651 = 12'h48e == _T_6[11:0] ? ram_1166 : _GEN_7650; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7652 = 12'h48f == _T_6[11:0] ? ram_1167 : _GEN_7651; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7653 = 12'h490 == _T_6[11:0] ? ram_1168 : _GEN_7652; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7654 = 12'h491 == _T_6[11:0] ? ram_1169 : _GEN_7653; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7655 = 12'h492 == _T_6[11:0] ? ram_1170 : _GEN_7654; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7656 = 12'h493 == _T_6[11:0] ? ram_1171 : _GEN_7655; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7657 = 12'h494 == _T_6[11:0] ? ram_1172 : _GEN_7656; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7658 = 12'h495 == _T_6[11:0] ? ram_1173 : _GEN_7657; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7659 = 12'h496 == _T_6[11:0] ? ram_1174 : _GEN_7658; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7660 = 12'h497 == _T_6[11:0] ? ram_1175 : _GEN_7659; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7661 = 12'h498 == _T_6[11:0] ? ram_1176 : _GEN_7660; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7662 = 12'h499 == _T_6[11:0] ? ram_1177 : _GEN_7661; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7663 = 12'h49a == _T_6[11:0] ? ram_1178 : _GEN_7662; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7664 = 12'h49b == _T_6[11:0] ? ram_1179 : _GEN_7663; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7665 = 12'h49c == _T_6[11:0] ? ram_1180 : _GEN_7664; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7666 = 12'h49d == _T_6[11:0] ? ram_1181 : _GEN_7665; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7667 = 12'h49e == _T_6[11:0] ? ram_1182 : _GEN_7666; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7668 = 12'h49f == _T_6[11:0] ? ram_1183 : _GEN_7667; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7669 = 12'h4a0 == _T_6[11:0] ? ram_1184 : _GEN_7668; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7670 = 12'h4a1 == _T_6[11:0] ? ram_1185 : _GEN_7669; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7671 = 12'h4a2 == _T_6[11:0] ? ram_1186 : _GEN_7670; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7672 = 12'h4a3 == _T_6[11:0] ? ram_1187 : _GEN_7671; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7673 = 12'h4a4 == _T_6[11:0] ? ram_1188 : _GEN_7672; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7674 = 12'h4a5 == _T_6[11:0] ? ram_1189 : _GEN_7673; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7675 = 12'h4a6 == _T_6[11:0] ? ram_1190 : _GEN_7674; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7676 = 12'h4a7 == _T_6[11:0] ? ram_1191 : _GEN_7675; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7677 = 12'h4a8 == _T_6[11:0] ? ram_1192 : _GEN_7676; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7678 = 12'h4a9 == _T_6[11:0] ? ram_1193 : _GEN_7677; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7679 = 12'h4aa == _T_6[11:0] ? ram_1194 : _GEN_7678; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7680 = 12'h4ab == _T_6[11:0] ? ram_1195 : _GEN_7679; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7681 = 12'h4ac == _T_6[11:0] ? ram_1196 : _GEN_7680; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7682 = 12'h4ad == _T_6[11:0] ? ram_1197 : _GEN_7681; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7683 = 12'h4ae == _T_6[11:0] ? ram_1198 : _GEN_7682; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7684 = 12'h4af == _T_6[11:0] ? ram_1199 : _GEN_7683; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7685 = 12'h4b0 == _T_6[11:0] ? ram_1200 : _GEN_7684; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7686 = 12'h4b1 == _T_6[11:0] ? ram_1201 : _GEN_7685; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7687 = 12'h4b2 == _T_6[11:0] ? ram_1202 : _GEN_7686; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7688 = 12'h4b3 == _T_6[11:0] ? ram_1203 : _GEN_7687; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7689 = 12'h4b4 == _T_6[11:0] ? ram_1204 : _GEN_7688; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7690 = 12'h4b5 == _T_6[11:0] ? ram_1205 : _GEN_7689; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7691 = 12'h4b6 == _T_6[11:0] ? ram_1206 : _GEN_7690; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7692 = 12'h4b7 == _T_6[11:0] ? ram_1207 : _GEN_7691; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7693 = 12'h4b8 == _T_6[11:0] ? ram_1208 : _GEN_7692; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7694 = 12'h4b9 == _T_6[11:0] ? ram_1209 : _GEN_7693; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7695 = 12'h4ba == _T_6[11:0] ? ram_1210 : _GEN_7694; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7696 = 12'h4bb == _T_6[11:0] ? ram_1211 : _GEN_7695; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7697 = 12'h4bc == _T_6[11:0] ? ram_1212 : _GEN_7696; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7698 = 12'h4bd == _T_6[11:0] ? ram_1213 : _GEN_7697; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7699 = 12'h4be == _T_6[11:0] ? ram_1214 : _GEN_7698; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7700 = 12'h4bf == _T_6[11:0] ? ram_1215 : _GEN_7699; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7701 = 12'h4c0 == _T_6[11:0] ? ram_1216 : _GEN_7700; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7702 = 12'h4c1 == _T_6[11:0] ? ram_1217 : _GEN_7701; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7703 = 12'h4c2 == _T_6[11:0] ? ram_1218 : _GEN_7702; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7704 = 12'h4c3 == _T_6[11:0] ? ram_1219 : _GEN_7703; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7705 = 12'h4c4 == _T_6[11:0] ? ram_1220 : _GEN_7704; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7706 = 12'h4c5 == _T_6[11:0] ? ram_1221 : _GEN_7705; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7707 = 12'h4c6 == _T_6[11:0] ? ram_1222 : _GEN_7706; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7708 = 12'h4c7 == _T_6[11:0] ? ram_1223 : _GEN_7707; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7709 = 12'h4c8 == _T_6[11:0] ? ram_1224 : _GEN_7708; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7710 = 12'h4c9 == _T_6[11:0] ? ram_1225 : _GEN_7709; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7711 = 12'h4ca == _T_6[11:0] ? ram_1226 : _GEN_7710; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7712 = 12'h4cb == _T_6[11:0] ? ram_1227 : _GEN_7711; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7713 = 12'h4cc == _T_6[11:0] ? ram_1228 : _GEN_7712; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7714 = 12'h4cd == _T_6[11:0] ? ram_1229 : _GEN_7713; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7715 = 12'h4ce == _T_6[11:0] ? ram_1230 : _GEN_7714; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7716 = 12'h4cf == _T_6[11:0] ? ram_1231 : _GEN_7715; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7717 = 12'h4d0 == _T_6[11:0] ? ram_1232 : _GEN_7716; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7718 = 12'h4d1 == _T_6[11:0] ? ram_1233 : _GEN_7717; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7719 = 12'h4d2 == _T_6[11:0] ? ram_1234 : _GEN_7718; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7720 = 12'h4d3 == _T_6[11:0] ? ram_1235 : _GEN_7719; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7721 = 12'h4d4 == _T_6[11:0] ? ram_1236 : _GEN_7720; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7722 = 12'h4d5 == _T_6[11:0] ? ram_1237 : _GEN_7721; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7723 = 12'h4d6 == _T_6[11:0] ? ram_1238 : _GEN_7722; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7724 = 12'h4d7 == _T_6[11:0] ? ram_1239 : _GEN_7723; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7725 = 12'h4d8 == _T_6[11:0] ? ram_1240 : _GEN_7724; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7726 = 12'h4d9 == _T_6[11:0] ? ram_1241 : _GEN_7725; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7727 = 12'h4da == _T_6[11:0] ? ram_1242 : _GEN_7726; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7728 = 12'h4db == _T_6[11:0] ? ram_1243 : _GEN_7727; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7729 = 12'h4dc == _T_6[11:0] ? ram_1244 : _GEN_7728; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7730 = 12'h4dd == _T_6[11:0] ? ram_1245 : _GEN_7729; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7731 = 12'h4de == _T_6[11:0] ? ram_1246 : _GEN_7730; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7732 = 12'h4df == _T_6[11:0] ? ram_1247 : _GEN_7731; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7733 = 12'h4e0 == _T_6[11:0] ? ram_1248 : _GEN_7732; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7734 = 12'h4e1 == _T_6[11:0] ? ram_1249 : _GEN_7733; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7735 = 12'h4e2 == _T_6[11:0] ? ram_1250 : _GEN_7734; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7736 = 12'h4e3 == _T_6[11:0] ? ram_1251 : _GEN_7735; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7737 = 12'h4e4 == _T_6[11:0] ? ram_1252 : _GEN_7736; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7738 = 12'h4e5 == _T_6[11:0] ? ram_1253 : _GEN_7737; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7739 = 12'h4e6 == _T_6[11:0] ? ram_1254 : _GEN_7738; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7740 = 12'h4e7 == _T_6[11:0] ? ram_1255 : _GEN_7739; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7741 = 12'h4e8 == _T_6[11:0] ? ram_1256 : _GEN_7740; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7742 = 12'h4e9 == _T_6[11:0] ? ram_1257 : _GEN_7741; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7743 = 12'h4ea == _T_6[11:0] ? ram_1258 : _GEN_7742; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7744 = 12'h4eb == _T_6[11:0] ? ram_1259 : _GEN_7743; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7745 = 12'h4ec == _T_6[11:0] ? ram_1260 : _GEN_7744; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7746 = 12'h4ed == _T_6[11:0] ? ram_1261 : _GEN_7745; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7747 = 12'h4ee == _T_6[11:0] ? ram_1262 : _GEN_7746; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7748 = 12'h4ef == _T_6[11:0] ? ram_1263 : _GEN_7747; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7749 = 12'h4f0 == _T_6[11:0] ? ram_1264 : _GEN_7748; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7750 = 12'h4f1 == _T_6[11:0] ? ram_1265 : _GEN_7749; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7751 = 12'h4f2 == _T_6[11:0] ? ram_1266 : _GEN_7750; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7752 = 12'h4f3 == _T_6[11:0] ? ram_1267 : _GEN_7751; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7753 = 12'h4f4 == _T_6[11:0] ? ram_1268 : _GEN_7752; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7754 = 12'h4f5 == _T_6[11:0] ? ram_1269 : _GEN_7753; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7755 = 12'h4f6 == _T_6[11:0] ? ram_1270 : _GEN_7754; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7756 = 12'h4f7 == _T_6[11:0] ? ram_1271 : _GEN_7755; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7757 = 12'h4f8 == _T_6[11:0] ? ram_1272 : _GEN_7756; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7758 = 12'h4f9 == _T_6[11:0] ? ram_1273 : _GEN_7757; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7759 = 12'h4fa == _T_6[11:0] ? ram_1274 : _GEN_7758; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7760 = 12'h4fb == _T_6[11:0] ? ram_1275 : _GEN_7759; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7761 = 12'h4fc == _T_6[11:0] ? ram_1276 : _GEN_7760; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7762 = 12'h4fd == _T_6[11:0] ? ram_1277 : _GEN_7761; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7763 = 12'h4fe == _T_6[11:0] ? ram_1278 : _GEN_7762; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7764 = 12'h4ff == _T_6[11:0] ? ram_1279 : _GEN_7763; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7765 = 12'h500 == _T_6[11:0] ? ram_1280 : _GEN_7764; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7766 = 12'h501 == _T_6[11:0] ? ram_1281 : _GEN_7765; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7767 = 12'h502 == _T_6[11:0] ? ram_1282 : _GEN_7766; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7768 = 12'h503 == _T_6[11:0] ? ram_1283 : _GEN_7767; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7769 = 12'h504 == _T_6[11:0] ? ram_1284 : _GEN_7768; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7770 = 12'h505 == _T_6[11:0] ? ram_1285 : _GEN_7769; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7771 = 12'h506 == _T_6[11:0] ? ram_1286 : _GEN_7770; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7772 = 12'h507 == _T_6[11:0] ? ram_1287 : _GEN_7771; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7773 = 12'h508 == _T_6[11:0] ? ram_1288 : _GEN_7772; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7774 = 12'h509 == _T_6[11:0] ? ram_1289 : _GEN_7773; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7775 = 12'h50a == _T_6[11:0] ? ram_1290 : _GEN_7774; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7776 = 12'h50b == _T_6[11:0] ? ram_1291 : _GEN_7775; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7777 = 12'h50c == _T_6[11:0] ? ram_1292 : _GEN_7776; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7778 = 12'h50d == _T_6[11:0] ? ram_1293 : _GEN_7777; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7779 = 12'h50e == _T_6[11:0] ? ram_1294 : _GEN_7778; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7780 = 12'h50f == _T_6[11:0] ? ram_1295 : _GEN_7779; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7781 = 12'h510 == _T_6[11:0] ? ram_1296 : _GEN_7780; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7782 = 12'h511 == _T_6[11:0] ? ram_1297 : _GEN_7781; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7783 = 12'h512 == _T_6[11:0] ? ram_1298 : _GEN_7782; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7784 = 12'h513 == _T_6[11:0] ? ram_1299 : _GEN_7783; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7785 = 12'h514 == _T_6[11:0] ? ram_1300 : _GEN_7784; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7786 = 12'h515 == _T_6[11:0] ? ram_1301 : _GEN_7785; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7787 = 12'h516 == _T_6[11:0] ? ram_1302 : _GEN_7786; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7788 = 12'h517 == _T_6[11:0] ? ram_1303 : _GEN_7787; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7789 = 12'h518 == _T_6[11:0] ? ram_1304 : _GEN_7788; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7790 = 12'h519 == _T_6[11:0] ? ram_1305 : _GEN_7789; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7791 = 12'h51a == _T_6[11:0] ? ram_1306 : _GEN_7790; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7792 = 12'h51b == _T_6[11:0] ? ram_1307 : _GEN_7791; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7793 = 12'h51c == _T_6[11:0] ? ram_1308 : _GEN_7792; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7794 = 12'h51d == _T_6[11:0] ? ram_1309 : _GEN_7793; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7795 = 12'h51e == _T_6[11:0] ? ram_1310 : _GEN_7794; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7796 = 12'h51f == _T_6[11:0] ? ram_1311 : _GEN_7795; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7797 = 12'h520 == _T_6[11:0] ? ram_1312 : _GEN_7796; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7798 = 12'h521 == _T_6[11:0] ? ram_1313 : _GEN_7797; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7799 = 12'h522 == _T_6[11:0] ? ram_1314 : _GEN_7798; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7800 = 12'h523 == _T_6[11:0] ? ram_1315 : _GEN_7799; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7801 = 12'h524 == _T_6[11:0] ? ram_1316 : _GEN_7800; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7802 = 12'h525 == _T_6[11:0] ? ram_1317 : _GEN_7801; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7803 = 12'h526 == _T_6[11:0] ? ram_1318 : _GEN_7802; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7804 = 12'h527 == _T_6[11:0] ? ram_1319 : _GEN_7803; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7805 = 12'h528 == _T_6[11:0] ? ram_1320 : _GEN_7804; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7806 = 12'h529 == _T_6[11:0] ? ram_1321 : _GEN_7805; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7807 = 12'h52a == _T_6[11:0] ? ram_1322 : _GEN_7806; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7808 = 12'h52b == _T_6[11:0] ? ram_1323 : _GEN_7807; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7809 = 12'h52c == _T_6[11:0] ? ram_1324 : _GEN_7808; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7810 = 12'h52d == _T_6[11:0] ? ram_1325 : _GEN_7809; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7811 = 12'h52e == _T_6[11:0] ? ram_1326 : _GEN_7810; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7812 = 12'h52f == _T_6[11:0] ? ram_1327 : _GEN_7811; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7813 = 12'h530 == _T_6[11:0] ? ram_1328 : _GEN_7812; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7814 = 12'h531 == _T_6[11:0] ? ram_1329 : _GEN_7813; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7815 = 12'h532 == _T_6[11:0] ? ram_1330 : _GEN_7814; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7816 = 12'h533 == _T_6[11:0] ? ram_1331 : _GEN_7815; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7817 = 12'h534 == _T_6[11:0] ? ram_1332 : _GEN_7816; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7818 = 12'h535 == _T_6[11:0] ? ram_1333 : _GEN_7817; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7819 = 12'h536 == _T_6[11:0] ? ram_1334 : _GEN_7818; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7820 = 12'h537 == _T_6[11:0] ? ram_1335 : _GEN_7819; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7821 = 12'h538 == _T_6[11:0] ? ram_1336 : _GEN_7820; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7822 = 12'h539 == _T_6[11:0] ? ram_1337 : _GEN_7821; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7823 = 12'h53a == _T_6[11:0] ? ram_1338 : _GEN_7822; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7824 = 12'h53b == _T_6[11:0] ? ram_1339 : _GEN_7823; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7825 = 12'h53c == _T_6[11:0] ? ram_1340 : _GEN_7824; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7826 = 12'h53d == _T_6[11:0] ? ram_1341 : _GEN_7825; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7827 = 12'h53e == _T_6[11:0] ? ram_1342 : _GEN_7826; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7828 = 12'h53f == _T_6[11:0] ? ram_1343 : _GEN_7827; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7829 = 12'h540 == _T_6[11:0] ? ram_1344 : _GEN_7828; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7830 = 12'h541 == _T_6[11:0] ? ram_1345 : _GEN_7829; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7831 = 12'h542 == _T_6[11:0] ? ram_1346 : _GEN_7830; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7832 = 12'h543 == _T_6[11:0] ? ram_1347 : _GEN_7831; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7833 = 12'h544 == _T_6[11:0] ? ram_1348 : _GEN_7832; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7834 = 12'h545 == _T_6[11:0] ? ram_1349 : _GEN_7833; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7835 = 12'h546 == _T_6[11:0] ? ram_1350 : _GEN_7834; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7836 = 12'h547 == _T_6[11:0] ? ram_1351 : _GEN_7835; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7837 = 12'h548 == _T_6[11:0] ? ram_1352 : _GEN_7836; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7838 = 12'h549 == _T_6[11:0] ? ram_1353 : _GEN_7837; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7839 = 12'h54a == _T_6[11:0] ? ram_1354 : _GEN_7838; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7840 = 12'h54b == _T_6[11:0] ? ram_1355 : _GEN_7839; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7841 = 12'h54c == _T_6[11:0] ? ram_1356 : _GEN_7840; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7842 = 12'h54d == _T_6[11:0] ? ram_1357 : _GEN_7841; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7843 = 12'h54e == _T_6[11:0] ? ram_1358 : _GEN_7842; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7844 = 12'h54f == _T_6[11:0] ? ram_1359 : _GEN_7843; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7845 = 12'h550 == _T_6[11:0] ? ram_1360 : _GEN_7844; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7846 = 12'h551 == _T_6[11:0] ? ram_1361 : _GEN_7845; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7847 = 12'h552 == _T_6[11:0] ? ram_1362 : _GEN_7846; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7848 = 12'h553 == _T_6[11:0] ? ram_1363 : _GEN_7847; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7849 = 12'h554 == _T_6[11:0] ? ram_1364 : _GEN_7848; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7850 = 12'h555 == _T_6[11:0] ? ram_1365 : _GEN_7849; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7851 = 12'h556 == _T_6[11:0] ? ram_1366 : _GEN_7850; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7852 = 12'h557 == _T_6[11:0] ? ram_1367 : _GEN_7851; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7853 = 12'h558 == _T_6[11:0] ? ram_1368 : _GEN_7852; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7854 = 12'h559 == _T_6[11:0] ? ram_1369 : _GEN_7853; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7855 = 12'h55a == _T_6[11:0] ? ram_1370 : _GEN_7854; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7856 = 12'h55b == _T_6[11:0] ? ram_1371 : _GEN_7855; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7857 = 12'h55c == _T_6[11:0] ? ram_1372 : _GEN_7856; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7858 = 12'h55d == _T_6[11:0] ? ram_1373 : _GEN_7857; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7859 = 12'h55e == _T_6[11:0] ? ram_1374 : _GEN_7858; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7860 = 12'h55f == _T_6[11:0] ? ram_1375 : _GEN_7859; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7861 = 12'h560 == _T_6[11:0] ? ram_1376 : _GEN_7860; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7862 = 12'h561 == _T_6[11:0] ? ram_1377 : _GEN_7861; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7863 = 12'h562 == _T_6[11:0] ? ram_1378 : _GEN_7862; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7864 = 12'h563 == _T_6[11:0] ? ram_1379 : _GEN_7863; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7865 = 12'h564 == _T_6[11:0] ? ram_1380 : _GEN_7864; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7866 = 12'h565 == _T_6[11:0] ? ram_1381 : _GEN_7865; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7867 = 12'h566 == _T_6[11:0] ? ram_1382 : _GEN_7866; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7868 = 12'h567 == _T_6[11:0] ? ram_1383 : _GEN_7867; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7869 = 12'h568 == _T_6[11:0] ? ram_1384 : _GEN_7868; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7870 = 12'h569 == _T_6[11:0] ? ram_1385 : _GEN_7869; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7871 = 12'h56a == _T_6[11:0] ? ram_1386 : _GEN_7870; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7872 = 12'h56b == _T_6[11:0] ? ram_1387 : _GEN_7871; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7873 = 12'h56c == _T_6[11:0] ? ram_1388 : _GEN_7872; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7874 = 12'h56d == _T_6[11:0] ? ram_1389 : _GEN_7873; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7875 = 12'h56e == _T_6[11:0] ? ram_1390 : _GEN_7874; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7876 = 12'h56f == _T_6[11:0] ? ram_1391 : _GEN_7875; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7877 = 12'h570 == _T_6[11:0] ? ram_1392 : _GEN_7876; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7878 = 12'h571 == _T_6[11:0] ? ram_1393 : _GEN_7877; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7879 = 12'h572 == _T_6[11:0] ? ram_1394 : _GEN_7878; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7880 = 12'h573 == _T_6[11:0] ? ram_1395 : _GEN_7879; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7881 = 12'h574 == _T_6[11:0] ? ram_1396 : _GEN_7880; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7882 = 12'h575 == _T_6[11:0] ? ram_1397 : _GEN_7881; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7883 = 12'h576 == _T_6[11:0] ? ram_1398 : _GEN_7882; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7884 = 12'h577 == _T_6[11:0] ? ram_1399 : _GEN_7883; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7885 = 12'h578 == _T_6[11:0] ? ram_1400 : _GEN_7884; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7886 = 12'h579 == _T_6[11:0] ? ram_1401 : _GEN_7885; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7887 = 12'h57a == _T_6[11:0] ? ram_1402 : _GEN_7886; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7888 = 12'h57b == _T_6[11:0] ? ram_1403 : _GEN_7887; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7889 = 12'h57c == _T_6[11:0] ? ram_1404 : _GEN_7888; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7890 = 12'h57d == _T_6[11:0] ? ram_1405 : _GEN_7889; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7891 = 12'h57e == _T_6[11:0] ? ram_1406 : _GEN_7890; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7892 = 12'h57f == _T_6[11:0] ? ram_1407 : _GEN_7891; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7893 = 12'h580 == _T_6[11:0] ? ram_1408 : _GEN_7892; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7894 = 12'h581 == _T_6[11:0] ? ram_1409 : _GEN_7893; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7895 = 12'h582 == _T_6[11:0] ? ram_1410 : _GEN_7894; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7896 = 12'h583 == _T_6[11:0] ? ram_1411 : _GEN_7895; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7897 = 12'h584 == _T_6[11:0] ? ram_1412 : _GEN_7896; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7898 = 12'h585 == _T_6[11:0] ? ram_1413 : _GEN_7897; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7899 = 12'h586 == _T_6[11:0] ? ram_1414 : _GEN_7898; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7900 = 12'h587 == _T_6[11:0] ? ram_1415 : _GEN_7899; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7901 = 12'h588 == _T_6[11:0] ? ram_1416 : _GEN_7900; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7902 = 12'h589 == _T_6[11:0] ? ram_1417 : _GEN_7901; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7903 = 12'h58a == _T_6[11:0] ? ram_1418 : _GEN_7902; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7904 = 12'h58b == _T_6[11:0] ? ram_1419 : _GEN_7903; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7905 = 12'h58c == _T_6[11:0] ? ram_1420 : _GEN_7904; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7906 = 12'h58d == _T_6[11:0] ? ram_1421 : _GEN_7905; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7907 = 12'h58e == _T_6[11:0] ? ram_1422 : _GEN_7906; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7908 = 12'h58f == _T_6[11:0] ? ram_1423 : _GEN_7907; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7909 = 12'h590 == _T_6[11:0] ? ram_1424 : _GEN_7908; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7910 = 12'h591 == _T_6[11:0] ? ram_1425 : _GEN_7909; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7911 = 12'h592 == _T_6[11:0] ? ram_1426 : _GEN_7910; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7912 = 12'h593 == _T_6[11:0] ? ram_1427 : _GEN_7911; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7913 = 12'h594 == _T_6[11:0] ? ram_1428 : _GEN_7912; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7914 = 12'h595 == _T_6[11:0] ? ram_1429 : _GEN_7913; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7915 = 12'h596 == _T_6[11:0] ? ram_1430 : _GEN_7914; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7916 = 12'h597 == _T_6[11:0] ? ram_1431 : _GEN_7915; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7917 = 12'h598 == _T_6[11:0] ? ram_1432 : _GEN_7916; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7918 = 12'h599 == _T_6[11:0] ? ram_1433 : _GEN_7917; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7919 = 12'h59a == _T_6[11:0] ? ram_1434 : _GEN_7918; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7920 = 12'h59b == _T_6[11:0] ? ram_1435 : _GEN_7919; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7921 = 12'h59c == _T_6[11:0] ? ram_1436 : _GEN_7920; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7922 = 12'h59d == _T_6[11:0] ? ram_1437 : _GEN_7921; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7923 = 12'h59e == _T_6[11:0] ? ram_1438 : _GEN_7922; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7924 = 12'h59f == _T_6[11:0] ? ram_1439 : _GEN_7923; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7925 = 12'h5a0 == _T_6[11:0] ? ram_1440 : _GEN_7924; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7926 = 12'h5a1 == _T_6[11:0] ? ram_1441 : _GEN_7925; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7927 = 12'h5a2 == _T_6[11:0] ? ram_1442 : _GEN_7926; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7928 = 12'h5a3 == _T_6[11:0] ? ram_1443 : _GEN_7927; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7929 = 12'h5a4 == _T_6[11:0] ? ram_1444 : _GEN_7928; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7930 = 12'h5a5 == _T_6[11:0] ? ram_1445 : _GEN_7929; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7931 = 12'h5a6 == _T_6[11:0] ? ram_1446 : _GEN_7930; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7932 = 12'h5a7 == _T_6[11:0] ? ram_1447 : _GEN_7931; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7933 = 12'h5a8 == _T_6[11:0] ? ram_1448 : _GEN_7932; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7934 = 12'h5a9 == _T_6[11:0] ? ram_1449 : _GEN_7933; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7935 = 12'h5aa == _T_6[11:0] ? ram_1450 : _GEN_7934; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7936 = 12'h5ab == _T_6[11:0] ? ram_1451 : _GEN_7935; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7937 = 12'h5ac == _T_6[11:0] ? ram_1452 : _GEN_7936; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7938 = 12'h5ad == _T_6[11:0] ? ram_1453 : _GEN_7937; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7939 = 12'h5ae == _T_6[11:0] ? ram_1454 : _GEN_7938; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7940 = 12'h5af == _T_6[11:0] ? ram_1455 : _GEN_7939; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7941 = 12'h5b0 == _T_6[11:0] ? ram_1456 : _GEN_7940; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7942 = 12'h5b1 == _T_6[11:0] ? ram_1457 : _GEN_7941; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7943 = 12'h5b2 == _T_6[11:0] ? ram_1458 : _GEN_7942; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7944 = 12'h5b3 == _T_6[11:0] ? ram_1459 : _GEN_7943; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7945 = 12'h5b4 == _T_6[11:0] ? ram_1460 : _GEN_7944; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7946 = 12'h5b5 == _T_6[11:0] ? ram_1461 : _GEN_7945; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7947 = 12'h5b6 == _T_6[11:0] ? ram_1462 : _GEN_7946; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7948 = 12'h5b7 == _T_6[11:0] ? ram_1463 : _GEN_7947; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7949 = 12'h5b8 == _T_6[11:0] ? ram_1464 : _GEN_7948; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7950 = 12'h5b9 == _T_6[11:0] ? ram_1465 : _GEN_7949; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7951 = 12'h5ba == _T_6[11:0] ? ram_1466 : _GEN_7950; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7952 = 12'h5bb == _T_6[11:0] ? ram_1467 : _GEN_7951; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7953 = 12'h5bc == _T_6[11:0] ? ram_1468 : _GEN_7952; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7954 = 12'h5bd == _T_6[11:0] ? ram_1469 : _GEN_7953; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7955 = 12'h5be == _T_6[11:0] ? ram_1470 : _GEN_7954; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7956 = 12'h5bf == _T_6[11:0] ? ram_1471 : _GEN_7955; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7957 = 12'h5c0 == _T_6[11:0] ? ram_1472 : _GEN_7956; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7958 = 12'h5c1 == _T_6[11:0] ? ram_1473 : _GEN_7957; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7959 = 12'h5c2 == _T_6[11:0] ? ram_1474 : _GEN_7958; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7960 = 12'h5c3 == _T_6[11:0] ? ram_1475 : _GEN_7959; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7961 = 12'h5c4 == _T_6[11:0] ? ram_1476 : _GEN_7960; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7962 = 12'h5c5 == _T_6[11:0] ? ram_1477 : _GEN_7961; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7963 = 12'h5c6 == _T_6[11:0] ? ram_1478 : _GEN_7962; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7964 = 12'h5c7 == _T_6[11:0] ? ram_1479 : _GEN_7963; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7965 = 12'h5c8 == _T_6[11:0] ? ram_1480 : _GEN_7964; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7966 = 12'h5c9 == _T_6[11:0] ? ram_1481 : _GEN_7965; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7967 = 12'h5ca == _T_6[11:0] ? ram_1482 : _GEN_7966; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7968 = 12'h5cb == _T_6[11:0] ? ram_1483 : _GEN_7967; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7969 = 12'h5cc == _T_6[11:0] ? ram_1484 : _GEN_7968; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7970 = 12'h5cd == _T_6[11:0] ? ram_1485 : _GEN_7969; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7971 = 12'h5ce == _T_6[11:0] ? ram_1486 : _GEN_7970; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7972 = 12'h5cf == _T_6[11:0] ? ram_1487 : _GEN_7971; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7973 = 12'h5d0 == _T_6[11:0] ? ram_1488 : _GEN_7972; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7974 = 12'h5d1 == _T_6[11:0] ? ram_1489 : _GEN_7973; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7975 = 12'h5d2 == _T_6[11:0] ? ram_1490 : _GEN_7974; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7976 = 12'h5d3 == _T_6[11:0] ? ram_1491 : _GEN_7975; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7977 = 12'h5d4 == _T_6[11:0] ? ram_1492 : _GEN_7976; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7978 = 12'h5d5 == _T_6[11:0] ? ram_1493 : _GEN_7977; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7979 = 12'h5d6 == _T_6[11:0] ? ram_1494 : _GEN_7978; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7980 = 12'h5d7 == _T_6[11:0] ? ram_1495 : _GEN_7979; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7981 = 12'h5d8 == _T_6[11:0] ? ram_1496 : _GEN_7980; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7982 = 12'h5d9 == _T_6[11:0] ? ram_1497 : _GEN_7981; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7983 = 12'h5da == _T_6[11:0] ? ram_1498 : _GEN_7982; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7984 = 12'h5db == _T_6[11:0] ? ram_1499 : _GEN_7983; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7985 = 12'h5dc == _T_6[11:0] ? ram_1500 : _GEN_7984; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7986 = 12'h5dd == _T_6[11:0] ? ram_1501 : _GEN_7985; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7987 = 12'h5de == _T_6[11:0] ? ram_1502 : _GEN_7986; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7988 = 12'h5df == _T_6[11:0] ? ram_1503 : _GEN_7987; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7989 = 12'h5e0 == _T_6[11:0] ? ram_1504 : _GEN_7988; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7990 = 12'h5e1 == _T_6[11:0] ? ram_1505 : _GEN_7989; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7991 = 12'h5e2 == _T_6[11:0] ? ram_1506 : _GEN_7990; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7992 = 12'h5e3 == _T_6[11:0] ? ram_1507 : _GEN_7991; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7993 = 12'h5e4 == _T_6[11:0] ? ram_1508 : _GEN_7992; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7994 = 12'h5e5 == _T_6[11:0] ? ram_1509 : _GEN_7993; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7995 = 12'h5e6 == _T_6[11:0] ? ram_1510 : _GEN_7994; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7996 = 12'h5e7 == _T_6[11:0] ? ram_1511 : _GEN_7995; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7997 = 12'h5e8 == _T_6[11:0] ? ram_1512 : _GEN_7996; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7998 = 12'h5e9 == _T_6[11:0] ? ram_1513 : _GEN_7997; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_7999 = 12'h5ea == _T_6[11:0] ? ram_1514 : _GEN_7998; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8000 = 12'h5eb == _T_6[11:0] ? ram_1515 : _GEN_7999; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8001 = 12'h5ec == _T_6[11:0] ? ram_1516 : _GEN_8000; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8002 = 12'h5ed == _T_6[11:0] ? ram_1517 : _GEN_8001; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8003 = 12'h5ee == _T_6[11:0] ? ram_1518 : _GEN_8002; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8004 = 12'h5ef == _T_6[11:0] ? ram_1519 : _GEN_8003; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8005 = 12'h5f0 == _T_6[11:0] ? ram_1520 : _GEN_8004; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8006 = 12'h5f1 == _T_6[11:0] ? ram_1521 : _GEN_8005; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8007 = 12'h5f2 == _T_6[11:0] ? ram_1522 : _GEN_8006; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8008 = 12'h5f3 == _T_6[11:0] ? ram_1523 : _GEN_8007; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8009 = 12'h5f4 == _T_6[11:0] ? ram_1524 : _GEN_8008; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8010 = 12'h5f5 == _T_6[11:0] ? ram_1525 : _GEN_8009; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8011 = 12'h5f6 == _T_6[11:0] ? ram_1526 : _GEN_8010; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8012 = 12'h5f7 == _T_6[11:0] ? ram_1527 : _GEN_8011; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8013 = 12'h5f8 == _T_6[11:0] ? ram_1528 : _GEN_8012; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8014 = 12'h5f9 == _T_6[11:0] ? ram_1529 : _GEN_8013; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8015 = 12'h5fa == _T_6[11:0] ? ram_1530 : _GEN_8014; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8016 = 12'h5fb == _T_6[11:0] ? ram_1531 : _GEN_8015; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8017 = 12'h5fc == _T_6[11:0] ? ram_1532 : _GEN_8016; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8018 = 12'h5fd == _T_6[11:0] ? ram_1533 : _GEN_8017; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8019 = 12'h5fe == _T_6[11:0] ? ram_1534 : _GEN_8018; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8020 = 12'h5ff == _T_6[11:0] ? ram_1535 : _GEN_8019; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8021 = 12'h600 == _T_6[11:0] ? ram_1536 : _GEN_8020; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8022 = 12'h601 == _T_6[11:0] ? ram_1537 : _GEN_8021; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8023 = 12'h602 == _T_6[11:0] ? ram_1538 : _GEN_8022; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8024 = 12'h603 == _T_6[11:0] ? ram_1539 : _GEN_8023; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8025 = 12'h604 == _T_6[11:0] ? ram_1540 : _GEN_8024; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8026 = 12'h605 == _T_6[11:0] ? ram_1541 : _GEN_8025; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8027 = 12'h606 == _T_6[11:0] ? ram_1542 : _GEN_8026; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8028 = 12'h607 == _T_6[11:0] ? ram_1543 : _GEN_8027; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8029 = 12'h608 == _T_6[11:0] ? ram_1544 : _GEN_8028; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8030 = 12'h609 == _T_6[11:0] ? ram_1545 : _GEN_8029; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8031 = 12'h60a == _T_6[11:0] ? ram_1546 : _GEN_8030; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8032 = 12'h60b == _T_6[11:0] ? ram_1547 : _GEN_8031; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8033 = 12'h60c == _T_6[11:0] ? ram_1548 : _GEN_8032; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8034 = 12'h60d == _T_6[11:0] ? ram_1549 : _GEN_8033; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8035 = 12'h60e == _T_6[11:0] ? ram_1550 : _GEN_8034; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8036 = 12'h60f == _T_6[11:0] ? ram_1551 : _GEN_8035; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8037 = 12'h610 == _T_6[11:0] ? ram_1552 : _GEN_8036; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8038 = 12'h611 == _T_6[11:0] ? ram_1553 : _GEN_8037; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8039 = 12'h612 == _T_6[11:0] ? ram_1554 : _GEN_8038; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8040 = 12'h613 == _T_6[11:0] ? ram_1555 : _GEN_8039; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8041 = 12'h614 == _T_6[11:0] ? ram_1556 : _GEN_8040; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8042 = 12'h615 == _T_6[11:0] ? ram_1557 : _GEN_8041; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8043 = 12'h616 == _T_6[11:0] ? ram_1558 : _GEN_8042; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8044 = 12'h617 == _T_6[11:0] ? ram_1559 : _GEN_8043; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8045 = 12'h618 == _T_6[11:0] ? ram_1560 : _GEN_8044; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8046 = 12'h619 == _T_6[11:0] ? ram_1561 : _GEN_8045; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8047 = 12'h61a == _T_6[11:0] ? ram_1562 : _GEN_8046; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8048 = 12'h61b == _T_6[11:0] ? ram_1563 : _GEN_8047; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8049 = 12'h61c == _T_6[11:0] ? ram_1564 : _GEN_8048; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8050 = 12'h61d == _T_6[11:0] ? ram_1565 : _GEN_8049; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8051 = 12'h61e == _T_6[11:0] ? ram_1566 : _GEN_8050; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8052 = 12'h61f == _T_6[11:0] ? ram_1567 : _GEN_8051; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8053 = 12'h620 == _T_6[11:0] ? ram_1568 : _GEN_8052; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8054 = 12'h621 == _T_6[11:0] ? ram_1569 : _GEN_8053; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8055 = 12'h622 == _T_6[11:0] ? ram_1570 : _GEN_8054; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8056 = 12'h623 == _T_6[11:0] ? ram_1571 : _GEN_8055; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8057 = 12'h624 == _T_6[11:0] ? ram_1572 : _GEN_8056; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8058 = 12'h625 == _T_6[11:0] ? ram_1573 : _GEN_8057; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8059 = 12'h626 == _T_6[11:0] ? ram_1574 : _GEN_8058; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8060 = 12'h627 == _T_6[11:0] ? ram_1575 : _GEN_8059; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8061 = 12'h628 == _T_6[11:0] ? ram_1576 : _GEN_8060; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8062 = 12'h629 == _T_6[11:0] ? ram_1577 : _GEN_8061; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8063 = 12'h62a == _T_6[11:0] ? ram_1578 : _GEN_8062; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8064 = 12'h62b == _T_6[11:0] ? ram_1579 : _GEN_8063; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8065 = 12'h62c == _T_6[11:0] ? ram_1580 : _GEN_8064; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8066 = 12'h62d == _T_6[11:0] ? ram_1581 : _GEN_8065; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8067 = 12'h62e == _T_6[11:0] ? ram_1582 : _GEN_8066; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8068 = 12'h62f == _T_6[11:0] ? ram_1583 : _GEN_8067; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8069 = 12'h630 == _T_6[11:0] ? ram_1584 : _GEN_8068; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8070 = 12'h631 == _T_6[11:0] ? ram_1585 : _GEN_8069; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8071 = 12'h632 == _T_6[11:0] ? ram_1586 : _GEN_8070; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8072 = 12'h633 == _T_6[11:0] ? ram_1587 : _GEN_8071; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8073 = 12'h634 == _T_6[11:0] ? ram_1588 : _GEN_8072; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8074 = 12'h635 == _T_6[11:0] ? ram_1589 : _GEN_8073; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8075 = 12'h636 == _T_6[11:0] ? ram_1590 : _GEN_8074; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8076 = 12'h637 == _T_6[11:0] ? ram_1591 : _GEN_8075; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8077 = 12'h638 == _T_6[11:0] ? ram_1592 : _GEN_8076; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8078 = 12'h639 == _T_6[11:0] ? ram_1593 : _GEN_8077; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8079 = 12'h63a == _T_6[11:0] ? ram_1594 : _GEN_8078; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8080 = 12'h63b == _T_6[11:0] ? ram_1595 : _GEN_8079; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8081 = 12'h63c == _T_6[11:0] ? ram_1596 : _GEN_8080; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8082 = 12'h63d == _T_6[11:0] ? ram_1597 : _GEN_8081; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8083 = 12'h63e == _T_6[11:0] ? ram_1598 : _GEN_8082; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8084 = 12'h63f == _T_6[11:0] ? ram_1599 : _GEN_8083; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8085 = 12'h640 == _T_6[11:0] ? ram_1600 : _GEN_8084; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8086 = 12'h641 == _T_6[11:0] ? ram_1601 : _GEN_8085; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8087 = 12'h642 == _T_6[11:0] ? ram_1602 : _GEN_8086; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8088 = 12'h643 == _T_6[11:0] ? ram_1603 : _GEN_8087; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8089 = 12'h644 == _T_6[11:0] ? ram_1604 : _GEN_8088; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8090 = 12'h645 == _T_6[11:0] ? ram_1605 : _GEN_8089; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8091 = 12'h646 == _T_6[11:0] ? ram_1606 : _GEN_8090; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8092 = 12'h647 == _T_6[11:0] ? ram_1607 : _GEN_8091; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8093 = 12'h648 == _T_6[11:0] ? ram_1608 : _GEN_8092; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8094 = 12'h649 == _T_6[11:0] ? ram_1609 : _GEN_8093; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8095 = 12'h64a == _T_6[11:0] ? ram_1610 : _GEN_8094; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8096 = 12'h64b == _T_6[11:0] ? ram_1611 : _GEN_8095; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8097 = 12'h64c == _T_6[11:0] ? ram_1612 : _GEN_8096; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8098 = 12'h64d == _T_6[11:0] ? ram_1613 : _GEN_8097; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8099 = 12'h64e == _T_6[11:0] ? ram_1614 : _GEN_8098; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8100 = 12'h64f == _T_6[11:0] ? ram_1615 : _GEN_8099; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8101 = 12'h650 == _T_6[11:0] ? ram_1616 : _GEN_8100; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8102 = 12'h651 == _T_6[11:0] ? ram_1617 : _GEN_8101; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8103 = 12'h652 == _T_6[11:0] ? ram_1618 : _GEN_8102; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8104 = 12'h653 == _T_6[11:0] ? ram_1619 : _GEN_8103; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8105 = 12'h654 == _T_6[11:0] ? ram_1620 : _GEN_8104; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8106 = 12'h655 == _T_6[11:0] ? ram_1621 : _GEN_8105; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8107 = 12'h656 == _T_6[11:0] ? ram_1622 : _GEN_8106; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8108 = 12'h657 == _T_6[11:0] ? ram_1623 : _GEN_8107; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8109 = 12'h658 == _T_6[11:0] ? ram_1624 : _GEN_8108; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8110 = 12'h659 == _T_6[11:0] ? ram_1625 : _GEN_8109; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8111 = 12'h65a == _T_6[11:0] ? ram_1626 : _GEN_8110; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8112 = 12'h65b == _T_6[11:0] ? ram_1627 : _GEN_8111; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8113 = 12'h65c == _T_6[11:0] ? ram_1628 : _GEN_8112; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8114 = 12'h65d == _T_6[11:0] ? ram_1629 : _GEN_8113; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8115 = 12'h65e == _T_6[11:0] ? ram_1630 : _GEN_8114; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8116 = 12'h65f == _T_6[11:0] ? ram_1631 : _GEN_8115; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8117 = 12'h660 == _T_6[11:0] ? ram_1632 : _GEN_8116; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8118 = 12'h661 == _T_6[11:0] ? ram_1633 : _GEN_8117; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8119 = 12'h662 == _T_6[11:0] ? ram_1634 : _GEN_8118; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8120 = 12'h663 == _T_6[11:0] ? ram_1635 : _GEN_8119; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8121 = 12'h664 == _T_6[11:0] ? ram_1636 : _GEN_8120; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8122 = 12'h665 == _T_6[11:0] ? ram_1637 : _GEN_8121; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8123 = 12'h666 == _T_6[11:0] ? ram_1638 : _GEN_8122; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8124 = 12'h667 == _T_6[11:0] ? ram_1639 : _GEN_8123; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8125 = 12'h668 == _T_6[11:0] ? ram_1640 : _GEN_8124; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8126 = 12'h669 == _T_6[11:0] ? ram_1641 : _GEN_8125; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8127 = 12'h66a == _T_6[11:0] ? ram_1642 : _GEN_8126; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8128 = 12'h66b == _T_6[11:0] ? ram_1643 : _GEN_8127; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8129 = 12'h66c == _T_6[11:0] ? ram_1644 : _GEN_8128; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8130 = 12'h66d == _T_6[11:0] ? ram_1645 : _GEN_8129; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8131 = 12'h66e == _T_6[11:0] ? ram_1646 : _GEN_8130; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8132 = 12'h66f == _T_6[11:0] ? ram_1647 : _GEN_8131; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8133 = 12'h670 == _T_6[11:0] ? ram_1648 : _GEN_8132; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8134 = 12'h671 == _T_6[11:0] ? ram_1649 : _GEN_8133; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8135 = 12'h672 == _T_6[11:0] ? ram_1650 : _GEN_8134; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8136 = 12'h673 == _T_6[11:0] ? ram_1651 : _GEN_8135; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8137 = 12'h674 == _T_6[11:0] ? ram_1652 : _GEN_8136; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8138 = 12'h675 == _T_6[11:0] ? ram_1653 : _GEN_8137; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8139 = 12'h676 == _T_6[11:0] ? ram_1654 : _GEN_8138; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8140 = 12'h677 == _T_6[11:0] ? ram_1655 : _GEN_8139; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8141 = 12'h678 == _T_6[11:0] ? ram_1656 : _GEN_8140; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8142 = 12'h679 == _T_6[11:0] ? ram_1657 : _GEN_8141; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8143 = 12'h67a == _T_6[11:0] ? ram_1658 : _GEN_8142; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8144 = 12'h67b == _T_6[11:0] ? ram_1659 : _GEN_8143; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8145 = 12'h67c == _T_6[11:0] ? ram_1660 : _GEN_8144; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8146 = 12'h67d == _T_6[11:0] ? ram_1661 : _GEN_8145; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8147 = 12'h67e == _T_6[11:0] ? ram_1662 : _GEN_8146; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8148 = 12'h67f == _T_6[11:0] ? ram_1663 : _GEN_8147; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8149 = 12'h680 == _T_6[11:0] ? ram_1664 : _GEN_8148; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8150 = 12'h681 == _T_6[11:0] ? ram_1665 : _GEN_8149; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8151 = 12'h682 == _T_6[11:0] ? ram_1666 : _GEN_8150; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8152 = 12'h683 == _T_6[11:0] ? ram_1667 : _GEN_8151; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8153 = 12'h684 == _T_6[11:0] ? ram_1668 : _GEN_8152; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8154 = 12'h685 == _T_6[11:0] ? ram_1669 : _GEN_8153; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8155 = 12'h686 == _T_6[11:0] ? ram_1670 : _GEN_8154; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8156 = 12'h687 == _T_6[11:0] ? ram_1671 : _GEN_8155; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8157 = 12'h688 == _T_6[11:0] ? ram_1672 : _GEN_8156; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8158 = 12'h689 == _T_6[11:0] ? ram_1673 : _GEN_8157; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8159 = 12'h68a == _T_6[11:0] ? ram_1674 : _GEN_8158; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8160 = 12'h68b == _T_6[11:0] ? ram_1675 : _GEN_8159; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8161 = 12'h68c == _T_6[11:0] ? ram_1676 : _GEN_8160; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8162 = 12'h68d == _T_6[11:0] ? ram_1677 : _GEN_8161; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8163 = 12'h68e == _T_6[11:0] ? ram_1678 : _GEN_8162; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8164 = 12'h68f == _T_6[11:0] ? ram_1679 : _GEN_8163; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8165 = 12'h690 == _T_6[11:0] ? ram_1680 : _GEN_8164; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8166 = 12'h691 == _T_6[11:0] ? ram_1681 : _GEN_8165; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8167 = 12'h692 == _T_6[11:0] ? ram_1682 : _GEN_8166; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8168 = 12'h693 == _T_6[11:0] ? ram_1683 : _GEN_8167; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8169 = 12'h694 == _T_6[11:0] ? ram_1684 : _GEN_8168; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8170 = 12'h695 == _T_6[11:0] ? ram_1685 : _GEN_8169; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8171 = 12'h696 == _T_6[11:0] ? ram_1686 : _GEN_8170; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8172 = 12'h697 == _T_6[11:0] ? ram_1687 : _GEN_8171; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8173 = 12'h698 == _T_6[11:0] ? ram_1688 : _GEN_8172; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8174 = 12'h699 == _T_6[11:0] ? ram_1689 : _GEN_8173; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8175 = 12'h69a == _T_6[11:0] ? ram_1690 : _GEN_8174; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8176 = 12'h69b == _T_6[11:0] ? ram_1691 : _GEN_8175; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8177 = 12'h69c == _T_6[11:0] ? ram_1692 : _GEN_8176; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8178 = 12'h69d == _T_6[11:0] ? ram_1693 : _GEN_8177; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8179 = 12'h69e == _T_6[11:0] ? ram_1694 : _GEN_8178; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8180 = 12'h69f == _T_6[11:0] ? ram_1695 : _GEN_8179; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8181 = 12'h6a0 == _T_6[11:0] ? ram_1696 : _GEN_8180; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8182 = 12'h6a1 == _T_6[11:0] ? ram_1697 : _GEN_8181; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8183 = 12'h6a2 == _T_6[11:0] ? ram_1698 : _GEN_8182; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8184 = 12'h6a3 == _T_6[11:0] ? ram_1699 : _GEN_8183; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8185 = 12'h6a4 == _T_6[11:0] ? ram_1700 : _GEN_8184; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8186 = 12'h6a5 == _T_6[11:0] ? ram_1701 : _GEN_8185; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8187 = 12'h6a6 == _T_6[11:0] ? ram_1702 : _GEN_8186; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8188 = 12'h6a7 == _T_6[11:0] ? ram_1703 : _GEN_8187; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8189 = 12'h6a8 == _T_6[11:0] ? ram_1704 : _GEN_8188; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8190 = 12'h6a9 == _T_6[11:0] ? ram_1705 : _GEN_8189; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8191 = 12'h6aa == _T_6[11:0] ? ram_1706 : _GEN_8190; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8192 = 12'h6ab == _T_6[11:0] ? ram_1707 : _GEN_8191; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8193 = 12'h6ac == _T_6[11:0] ? ram_1708 : _GEN_8192; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8194 = 12'h6ad == _T_6[11:0] ? ram_1709 : _GEN_8193; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8195 = 12'h6ae == _T_6[11:0] ? ram_1710 : _GEN_8194; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8196 = 12'h6af == _T_6[11:0] ? ram_1711 : _GEN_8195; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8197 = 12'h6b0 == _T_6[11:0] ? ram_1712 : _GEN_8196; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8198 = 12'h6b1 == _T_6[11:0] ? ram_1713 : _GEN_8197; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8199 = 12'h6b2 == _T_6[11:0] ? ram_1714 : _GEN_8198; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8200 = 12'h6b3 == _T_6[11:0] ? ram_1715 : _GEN_8199; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8201 = 12'h6b4 == _T_6[11:0] ? ram_1716 : _GEN_8200; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8202 = 12'h6b5 == _T_6[11:0] ? ram_1717 : _GEN_8201; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8203 = 12'h6b6 == _T_6[11:0] ? ram_1718 : _GEN_8202; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8204 = 12'h6b7 == _T_6[11:0] ? ram_1719 : _GEN_8203; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8205 = 12'h6b8 == _T_6[11:0] ? ram_1720 : _GEN_8204; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8206 = 12'h6b9 == _T_6[11:0] ? ram_1721 : _GEN_8205; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8207 = 12'h6ba == _T_6[11:0] ? ram_1722 : _GEN_8206; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8208 = 12'h6bb == _T_6[11:0] ? ram_1723 : _GEN_8207; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8209 = 12'h6bc == _T_6[11:0] ? ram_1724 : _GEN_8208; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8210 = 12'h6bd == _T_6[11:0] ? ram_1725 : _GEN_8209; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8211 = 12'h6be == _T_6[11:0] ? ram_1726 : _GEN_8210; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8212 = 12'h6bf == _T_6[11:0] ? ram_1727 : _GEN_8211; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8213 = 12'h6c0 == _T_6[11:0] ? ram_1728 : _GEN_8212; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8214 = 12'h6c1 == _T_6[11:0] ? ram_1729 : _GEN_8213; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8215 = 12'h6c2 == _T_6[11:0] ? ram_1730 : _GEN_8214; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8216 = 12'h6c3 == _T_6[11:0] ? ram_1731 : _GEN_8215; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8217 = 12'h6c4 == _T_6[11:0] ? ram_1732 : _GEN_8216; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8218 = 12'h6c5 == _T_6[11:0] ? ram_1733 : _GEN_8217; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8219 = 12'h6c6 == _T_6[11:0] ? ram_1734 : _GEN_8218; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8220 = 12'h6c7 == _T_6[11:0] ? ram_1735 : _GEN_8219; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8221 = 12'h6c8 == _T_6[11:0] ? ram_1736 : _GEN_8220; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8222 = 12'h6c9 == _T_6[11:0] ? ram_1737 : _GEN_8221; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8223 = 12'h6ca == _T_6[11:0] ? ram_1738 : _GEN_8222; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8224 = 12'h6cb == _T_6[11:0] ? ram_1739 : _GEN_8223; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8225 = 12'h6cc == _T_6[11:0] ? ram_1740 : _GEN_8224; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8226 = 12'h6cd == _T_6[11:0] ? ram_1741 : _GEN_8225; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8227 = 12'h6ce == _T_6[11:0] ? ram_1742 : _GEN_8226; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8228 = 12'h6cf == _T_6[11:0] ? ram_1743 : _GEN_8227; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8229 = 12'h6d0 == _T_6[11:0] ? ram_1744 : _GEN_8228; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8230 = 12'h6d1 == _T_6[11:0] ? ram_1745 : _GEN_8229; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8231 = 12'h6d2 == _T_6[11:0] ? ram_1746 : _GEN_8230; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8232 = 12'h6d3 == _T_6[11:0] ? ram_1747 : _GEN_8231; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8233 = 12'h6d4 == _T_6[11:0] ? ram_1748 : _GEN_8232; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8234 = 12'h6d5 == _T_6[11:0] ? ram_1749 : _GEN_8233; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8235 = 12'h6d6 == _T_6[11:0] ? ram_1750 : _GEN_8234; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8236 = 12'h6d7 == _T_6[11:0] ? ram_1751 : _GEN_8235; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8237 = 12'h6d8 == _T_6[11:0] ? ram_1752 : _GEN_8236; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8238 = 12'h6d9 == _T_6[11:0] ? ram_1753 : _GEN_8237; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8239 = 12'h6da == _T_6[11:0] ? ram_1754 : _GEN_8238; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8240 = 12'h6db == _T_6[11:0] ? ram_1755 : _GEN_8239; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8241 = 12'h6dc == _T_6[11:0] ? ram_1756 : _GEN_8240; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8242 = 12'h6dd == _T_6[11:0] ? ram_1757 : _GEN_8241; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8243 = 12'h6de == _T_6[11:0] ? ram_1758 : _GEN_8242; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8244 = 12'h6df == _T_6[11:0] ? ram_1759 : _GEN_8243; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8245 = 12'h6e0 == _T_6[11:0] ? ram_1760 : _GEN_8244; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8246 = 12'h6e1 == _T_6[11:0] ? ram_1761 : _GEN_8245; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8247 = 12'h6e2 == _T_6[11:0] ? ram_1762 : _GEN_8246; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8248 = 12'h6e3 == _T_6[11:0] ? ram_1763 : _GEN_8247; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8249 = 12'h6e4 == _T_6[11:0] ? ram_1764 : _GEN_8248; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8250 = 12'h6e5 == _T_6[11:0] ? ram_1765 : _GEN_8249; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8251 = 12'h6e6 == _T_6[11:0] ? ram_1766 : _GEN_8250; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8252 = 12'h6e7 == _T_6[11:0] ? ram_1767 : _GEN_8251; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8253 = 12'h6e8 == _T_6[11:0] ? ram_1768 : _GEN_8252; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8254 = 12'h6e9 == _T_6[11:0] ? ram_1769 : _GEN_8253; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8255 = 12'h6ea == _T_6[11:0] ? ram_1770 : _GEN_8254; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8256 = 12'h6eb == _T_6[11:0] ? ram_1771 : _GEN_8255; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8257 = 12'h6ec == _T_6[11:0] ? ram_1772 : _GEN_8256; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8258 = 12'h6ed == _T_6[11:0] ? ram_1773 : _GEN_8257; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8259 = 12'h6ee == _T_6[11:0] ? ram_1774 : _GEN_8258; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8260 = 12'h6ef == _T_6[11:0] ? ram_1775 : _GEN_8259; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8261 = 12'h6f0 == _T_6[11:0] ? ram_1776 : _GEN_8260; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8262 = 12'h6f1 == _T_6[11:0] ? ram_1777 : _GEN_8261; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8263 = 12'h6f2 == _T_6[11:0] ? ram_1778 : _GEN_8262; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8264 = 12'h6f3 == _T_6[11:0] ? ram_1779 : _GEN_8263; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8265 = 12'h6f4 == _T_6[11:0] ? ram_1780 : _GEN_8264; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8266 = 12'h6f5 == _T_6[11:0] ? ram_1781 : _GEN_8265; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8267 = 12'h6f6 == _T_6[11:0] ? ram_1782 : _GEN_8266; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8268 = 12'h6f7 == _T_6[11:0] ? ram_1783 : _GEN_8267; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8269 = 12'h6f8 == _T_6[11:0] ? ram_1784 : _GEN_8268; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8270 = 12'h6f9 == _T_6[11:0] ? ram_1785 : _GEN_8269; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8271 = 12'h6fa == _T_6[11:0] ? ram_1786 : _GEN_8270; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8272 = 12'h6fb == _T_6[11:0] ? ram_1787 : _GEN_8271; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8273 = 12'h6fc == _T_6[11:0] ? ram_1788 : _GEN_8272; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8274 = 12'h6fd == _T_6[11:0] ? ram_1789 : _GEN_8273; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8275 = 12'h6fe == _T_6[11:0] ? ram_1790 : _GEN_8274; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8276 = 12'h6ff == _T_6[11:0] ? ram_1791 : _GEN_8275; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8277 = 12'h700 == _T_6[11:0] ? ram_1792 : _GEN_8276; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8278 = 12'h701 == _T_6[11:0] ? ram_1793 : _GEN_8277; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8279 = 12'h702 == _T_6[11:0] ? ram_1794 : _GEN_8278; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8280 = 12'h703 == _T_6[11:0] ? ram_1795 : _GEN_8279; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8281 = 12'h704 == _T_6[11:0] ? ram_1796 : _GEN_8280; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8282 = 12'h705 == _T_6[11:0] ? ram_1797 : _GEN_8281; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8283 = 12'h706 == _T_6[11:0] ? ram_1798 : _GEN_8282; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8284 = 12'h707 == _T_6[11:0] ? ram_1799 : _GEN_8283; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8285 = 12'h708 == _T_6[11:0] ? ram_1800 : _GEN_8284; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8286 = 12'h709 == _T_6[11:0] ? ram_1801 : _GEN_8285; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8287 = 12'h70a == _T_6[11:0] ? ram_1802 : _GEN_8286; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8288 = 12'h70b == _T_6[11:0] ? ram_1803 : _GEN_8287; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8289 = 12'h70c == _T_6[11:0] ? ram_1804 : _GEN_8288; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8290 = 12'h70d == _T_6[11:0] ? ram_1805 : _GEN_8289; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8291 = 12'h70e == _T_6[11:0] ? ram_1806 : _GEN_8290; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8292 = 12'h70f == _T_6[11:0] ? ram_1807 : _GEN_8291; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8293 = 12'h710 == _T_6[11:0] ? ram_1808 : _GEN_8292; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8294 = 12'h711 == _T_6[11:0] ? ram_1809 : _GEN_8293; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8295 = 12'h712 == _T_6[11:0] ? ram_1810 : _GEN_8294; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8296 = 12'h713 == _T_6[11:0] ? ram_1811 : _GEN_8295; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8297 = 12'h714 == _T_6[11:0] ? ram_1812 : _GEN_8296; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8298 = 12'h715 == _T_6[11:0] ? ram_1813 : _GEN_8297; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8299 = 12'h716 == _T_6[11:0] ? ram_1814 : _GEN_8298; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8300 = 12'h717 == _T_6[11:0] ? ram_1815 : _GEN_8299; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8301 = 12'h718 == _T_6[11:0] ? ram_1816 : _GEN_8300; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8302 = 12'h719 == _T_6[11:0] ? ram_1817 : _GEN_8301; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8303 = 12'h71a == _T_6[11:0] ? ram_1818 : _GEN_8302; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8304 = 12'h71b == _T_6[11:0] ? ram_1819 : _GEN_8303; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8305 = 12'h71c == _T_6[11:0] ? ram_1820 : _GEN_8304; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8306 = 12'h71d == _T_6[11:0] ? ram_1821 : _GEN_8305; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8307 = 12'h71e == _T_6[11:0] ? ram_1822 : _GEN_8306; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8308 = 12'h71f == _T_6[11:0] ? ram_1823 : _GEN_8307; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8309 = 12'h720 == _T_6[11:0] ? ram_1824 : _GEN_8308; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8310 = 12'h721 == _T_6[11:0] ? ram_1825 : _GEN_8309; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8311 = 12'h722 == _T_6[11:0] ? ram_1826 : _GEN_8310; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8312 = 12'h723 == _T_6[11:0] ? ram_1827 : _GEN_8311; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8313 = 12'h724 == _T_6[11:0] ? ram_1828 : _GEN_8312; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8314 = 12'h725 == _T_6[11:0] ? ram_1829 : _GEN_8313; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8315 = 12'h726 == _T_6[11:0] ? ram_1830 : _GEN_8314; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8316 = 12'h727 == _T_6[11:0] ? ram_1831 : _GEN_8315; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8317 = 12'h728 == _T_6[11:0] ? ram_1832 : _GEN_8316; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8318 = 12'h729 == _T_6[11:0] ? ram_1833 : _GEN_8317; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8319 = 12'h72a == _T_6[11:0] ? ram_1834 : _GEN_8318; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8320 = 12'h72b == _T_6[11:0] ? ram_1835 : _GEN_8319; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8321 = 12'h72c == _T_6[11:0] ? ram_1836 : _GEN_8320; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8322 = 12'h72d == _T_6[11:0] ? ram_1837 : _GEN_8321; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8323 = 12'h72e == _T_6[11:0] ? ram_1838 : _GEN_8322; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8324 = 12'h72f == _T_6[11:0] ? ram_1839 : _GEN_8323; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8325 = 12'h730 == _T_6[11:0] ? ram_1840 : _GEN_8324; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8326 = 12'h731 == _T_6[11:0] ? ram_1841 : _GEN_8325; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8327 = 12'h732 == _T_6[11:0] ? ram_1842 : _GEN_8326; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8328 = 12'h733 == _T_6[11:0] ? ram_1843 : _GEN_8327; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8329 = 12'h734 == _T_6[11:0] ? ram_1844 : _GEN_8328; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8330 = 12'h735 == _T_6[11:0] ? ram_1845 : _GEN_8329; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8331 = 12'h736 == _T_6[11:0] ? ram_1846 : _GEN_8330; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8332 = 12'h737 == _T_6[11:0] ? ram_1847 : _GEN_8331; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8333 = 12'h738 == _T_6[11:0] ? ram_1848 : _GEN_8332; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8334 = 12'h739 == _T_6[11:0] ? ram_1849 : _GEN_8333; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8335 = 12'h73a == _T_6[11:0] ? ram_1850 : _GEN_8334; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8336 = 12'h73b == _T_6[11:0] ? ram_1851 : _GEN_8335; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8337 = 12'h73c == _T_6[11:0] ? ram_1852 : _GEN_8336; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8338 = 12'h73d == _T_6[11:0] ? ram_1853 : _GEN_8337; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8339 = 12'h73e == _T_6[11:0] ? ram_1854 : _GEN_8338; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8340 = 12'h73f == _T_6[11:0] ? ram_1855 : _GEN_8339; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8341 = 12'h740 == _T_6[11:0] ? ram_1856 : _GEN_8340; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8342 = 12'h741 == _T_6[11:0] ? ram_1857 : _GEN_8341; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8343 = 12'h742 == _T_6[11:0] ? ram_1858 : _GEN_8342; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8344 = 12'h743 == _T_6[11:0] ? ram_1859 : _GEN_8343; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8345 = 12'h744 == _T_6[11:0] ? ram_1860 : _GEN_8344; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8346 = 12'h745 == _T_6[11:0] ? ram_1861 : _GEN_8345; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8347 = 12'h746 == _T_6[11:0] ? ram_1862 : _GEN_8346; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8348 = 12'h747 == _T_6[11:0] ? ram_1863 : _GEN_8347; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8349 = 12'h748 == _T_6[11:0] ? ram_1864 : _GEN_8348; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8350 = 12'h749 == _T_6[11:0] ? ram_1865 : _GEN_8349; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8351 = 12'h74a == _T_6[11:0] ? ram_1866 : _GEN_8350; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8352 = 12'h74b == _T_6[11:0] ? ram_1867 : _GEN_8351; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8353 = 12'h74c == _T_6[11:0] ? ram_1868 : _GEN_8352; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8354 = 12'h74d == _T_6[11:0] ? ram_1869 : _GEN_8353; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8355 = 12'h74e == _T_6[11:0] ? ram_1870 : _GEN_8354; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8356 = 12'h74f == _T_6[11:0] ? ram_1871 : _GEN_8355; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8357 = 12'h750 == _T_6[11:0] ? ram_1872 : _GEN_8356; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8358 = 12'h751 == _T_6[11:0] ? ram_1873 : _GEN_8357; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8359 = 12'h752 == _T_6[11:0] ? ram_1874 : _GEN_8358; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8360 = 12'h753 == _T_6[11:0] ? ram_1875 : _GEN_8359; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8361 = 12'h754 == _T_6[11:0] ? ram_1876 : _GEN_8360; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8362 = 12'h755 == _T_6[11:0] ? ram_1877 : _GEN_8361; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8363 = 12'h756 == _T_6[11:0] ? ram_1878 : _GEN_8362; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8364 = 12'h757 == _T_6[11:0] ? ram_1879 : _GEN_8363; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8365 = 12'h758 == _T_6[11:0] ? ram_1880 : _GEN_8364; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8366 = 12'h759 == _T_6[11:0] ? ram_1881 : _GEN_8365; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8367 = 12'h75a == _T_6[11:0] ? ram_1882 : _GEN_8366; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8368 = 12'h75b == _T_6[11:0] ? ram_1883 : _GEN_8367; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8369 = 12'h75c == _T_6[11:0] ? ram_1884 : _GEN_8368; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8370 = 12'h75d == _T_6[11:0] ? ram_1885 : _GEN_8369; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8371 = 12'h75e == _T_6[11:0] ? ram_1886 : _GEN_8370; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8372 = 12'h75f == _T_6[11:0] ? ram_1887 : _GEN_8371; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8373 = 12'h760 == _T_6[11:0] ? ram_1888 : _GEN_8372; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8374 = 12'h761 == _T_6[11:0] ? ram_1889 : _GEN_8373; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8375 = 12'h762 == _T_6[11:0] ? ram_1890 : _GEN_8374; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8376 = 12'h763 == _T_6[11:0] ? ram_1891 : _GEN_8375; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8377 = 12'h764 == _T_6[11:0] ? ram_1892 : _GEN_8376; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8378 = 12'h765 == _T_6[11:0] ? ram_1893 : _GEN_8377; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8379 = 12'h766 == _T_6[11:0] ? ram_1894 : _GEN_8378; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8380 = 12'h767 == _T_6[11:0] ? ram_1895 : _GEN_8379; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8381 = 12'h768 == _T_6[11:0] ? ram_1896 : _GEN_8380; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8382 = 12'h769 == _T_6[11:0] ? ram_1897 : _GEN_8381; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8383 = 12'h76a == _T_6[11:0] ? ram_1898 : _GEN_8382; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8384 = 12'h76b == _T_6[11:0] ? ram_1899 : _GEN_8383; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8385 = 12'h76c == _T_6[11:0] ? ram_1900 : _GEN_8384; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8386 = 12'h76d == _T_6[11:0] ? ram_1901 : _GEN_8385; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8387 = 12'h76e == _T_6[11:0] ? ram_1902 : _GEN_8386; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8388 = 12'h76f == _T_6[11:0] ? ram_1903 : _GEN_8387; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8389 = 12'h770 == _T_6[11:0] ? ram_1904 : _GEN_8388; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8390 = 12'h771 == _T_6[11:0] ? ram_1905 : _GEN_8389; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8391 = 12'h772 == _T_6[11:0] ? ram_1906 : _GEN_8390; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8392 = 12'h773 == _T_6[11:0] ? ram_1907 : _GEN_8391; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8393 = 12'h774 == _T_6[11:0] ? ram_1908 : _GEN_8392; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8394 = 12'h775 == _T_6[11:0] ? ram_1909 : _GEN_8393; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8395 = 12'h776 == _T_6[11:0] ? ram_1910 : _GEN_8394; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8396 = 12'h777 == _T_6[11:0] ? ram_1911 : _GEN_8395; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8397 = 12'h778 == _T_6[11:0] ? ram_1912 : _GEN_8396; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8398 = 12'h779 == _T_6[11:0] ? ram_1913 : _GEN_8397; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8399 = 12'h77a == _T_6[11:0] ? ram_1914 : _GEN_8398; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8400 = 12'h77b == _T_6[11:0] ? ram_1915 : _GEN_8399; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8401 = 12'h77c == _T_6[11:0] ? ram_1916 : _GEN_8400; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8402 = 12'h77d == _T_6[11:0] ? ram_1917 : _GEN_8401; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8403 = 12'h77e == _T_6[11:0] ? ram_1918 : _GEN_8402; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8404 = 12'h77f == _T_6[11:0] ? ram_1919 : _GEN_8403; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8405 = 12'h780 == _T_6[11:0] ? ram_1920 : _GEN_8404; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8406 = 12'h781 == _T_6[11:0] ? ram_1921 : _GEN_8405; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8407 = 12'h782 == _T_6[11:0] ? ram_1922 : _GEN_8406; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8408 = 12'h783 == _T_6[11:0] ? ram_1923 : _GEN_8407; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8409 = 12'h784 == _T_6[11:0] ? ram_1924 : _GEN_8408; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8410 = 12'h785 == _T_6[11:0] ? ram_1925 : _GEN_8409; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8411 = 12'h786 == _T_6[11:0] ? ram_1926 : _GEN_8410; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8412 = 12'h787 == _T_6[11:0] ? ram_1927 : _GEN_8411; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8413 = 12'h788 == _T_6[11:0] ? ram_1928 : _GEN_8412; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8414 = 12'h789 == _T_6[11:0] ? ram_1929 : _GEN_8413; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8415 = 12'h78a == _T_6[11:0] ? ram_1930 : _GEN_8414; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8416 = 12'h78b == _T_6[11:0] ? ram_1931 : _GEN_8415; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8417 = 12'h78c == _T_6[11:0] ? ram_1932 : _GEN_8416; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8418 = 12'h78d == _T_6[11:0] ? ram_1933 : _GEN_8417; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8419 = 12'h78e == _T_6[11:0] ? ram_1934 : _GEN_8418; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8420 = 12'h78f == _T_6[11:0] ? ram_1935 : _GEN_8419; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8421 = 12'h790 == _T_6[11:0] ? ram_1936 : _GEN_8420; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8422 = 12'h791 == _T_6[11:0] ? ram_1937 : _GEN_8421; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8423 = 12'h792 == _T_6[11:0] ? ram_1938 : _GEN_8422; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8424 = 12'h793 == _T_6[11:0] ? ram_1939 : _GEN_8423; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8425 = 12'h794 == _T_6[11:0] ? ram_1940 : _GEN_8424; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8426 = 12'h795 == _T_6[11:0] ? ram_1941 : _GEN_8425; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8427 = 12'h796 == _T_6[11:0] ? ram_1942 : _GEN_8426; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8428 = 12'h797 == _T_6[11:0] ? ram_1943 : _GEN_8427; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8429 = 12'h798 == _T_6[11:0] ? ram_1944 : _GEN_8428; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8430 = 12'h799 == _T_6[11:0] ? ram_1945 : _GEN_8429; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8431 = 12'h79a == _T_6[11:0] ? ram_1946 : _GEN_8430; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8432 = 12'h79b == _T_6[11:0] ? ram_1947 : _GEN_8431; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8433 = 12'h79c == _T_6[11:0] ? ram_1948 : _GEN_8432; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8434 = 12'h79d == _T_6[11:0] ? ram_1949 : _GEN_8433; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8435 = 12'h79e == _T_6[11:0] ? ram_1950 : _GEN_8434; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8436 = 12'h79f == _T_6[11:0] ? ram_1951 : _GEN_8435; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8437 = 12'h7a0 == _T_6[11:0] ? ram_1952 : _GEN_8436; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8438 = 12'h7a1 == _T_6[11:0] ? ram_1953 : _GEN_8437; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8439 = 12'h7a2 == _T_6[11:0] ? ram_1954 : _GEN_8438; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8440 = 12'h7a3 == _T_6[11:0] ? ram_1955 : _GEN_8439; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8441 = 12'h7a4 == _T_6[11:0] ? ram_1956 : _GEN_8440; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8442 = 12'h7a5 == _T_6[11:0] ? ram_1957 : _GEN_8441; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8443 = 12'h7a6 == _T_6[11:0] ? ram_1958 : _GEN_8442; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8444 = 12'h7a7 == _T_6[11:0] ? ram_1959 : _GEN_8443; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8445 = 12'h7a8 == _T_6[11:0] ? ram_1960 : _GEN_8444; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8446 = 12'h7a9 == _T_6[11:0] ? ram_1961 : _GEN_8445; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8447 = 12'h7aa == _T_6[11:0] ? ram_1962 : _GEN_8446; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8448 = 12'h7ab == _T_6[11:0] ? ram_1963 : _GEN_8447; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8449 = 12'h7ac == _T_6[11:0] ? ram_1964 : _GEN_8448; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8450 = 12'h7ad == _T_6[11:0] ? ram_1965 : _GEN_8449; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8451 = 12'h7ae == _T_6[11:0] ? ram_1966 : _GEN_8450; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8452 = 12'h7af == _T_6[11:0] ? ram_1967 : _GEN_8451; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8453 = 12'h7b0 == _T_6[11:0] ? ram_1968 : _GEN_8452; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8454 = 12'h7b1 == _T_6[11:0] ? ram_1969 : _GEN_8453; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8455 = 12'h7b2 == _T_6[11:0] ? ram_1970 : _GEN_8454; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8456 = 12'h7b3 == _T_6[11:0] ? ram_1971 : _GEN_8455; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8457 = 12'h7b4 == _T_6[11:0] ? ram_1972 : _GEN_8456; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8458 = 12'h7b5 == _T_6[11:0] ? ram_1973 : _GEN_8457; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8459 = 12'h7b6 == _T_6[11:0] ? ram_1974 : _GEN_8458; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8460 = 12'h7b7 == _T_6[11:0] ? ram_1975 : _GEN_8459; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8461 = 12'h7b8 == _T_6[11:0] ? ram_1976 : _GEN_8460; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8462 = 12'h7b9 == _T_6[11:0] ? ram_1977 : _GEN_8461; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8463 = 12'h7ba == _T_6[11:0] ? ram_1978 : _GEN_8462; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8464 = 12'h7bb == _T_6[11:0] ? ram_1979 : _GEN_8463; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8465 = 12'h7bc == _T_6[11:0] ? ram_1980 : _GEN_8464; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8466 = 12'h7bd == _T_6[11:0] ? ram_1981 : _GEN_8465; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8467 = 12'h7be == _T_6[11:0] ? ram_1982 : _GEN_8466; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8468 = 12'h7bf == _T_6[11:0] ? ram_1983 : _GEN_8467; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8469 = 12'h7c0 == _T_6[11:0] ? ram_1984 : _GEN_8468; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8470 = 12'h7c1 == _T_6[11:0] ? ram_1985 : _GEN_8469; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8471 = 12'h7c2 == _T_6[11:0] ? ram_1986 : _GEN_8470; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8472 = 12'h7c3 == _T_6[11:0] ? ram_1987 : _GEN_8471; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8473 = 12'h7c4 == _T_6[11:0] ? ram_1988 : _GEN_8472; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8474 = 12'h7c5 == _T_6[11:0] ? ram_1989 : _GEN_8473; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8475 = 12'h7c6 == _T_6[11:0] ? ram_1990 : _GEN_8474; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8476 = 12'h7c7 == _T_6[11:0] ? ram_1991 : _GEN_8475; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8477 = 12'h7c8 == _T_6[11:0] ? ram_1992 : _GEN_8476; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8478 = 12'h7c9 == _T_6[11:0] ? ram_1993 : _GEN_8477; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8479 = 12'h7ca == _T_6[11:0] ? ram_1994 : _GEN_8478; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8480 = 12'h7cb == _T_6[11:0] ? ram_1995 : _GEN_8479; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8481 = 12'h7cc == _T_6[11:0] ? ram_1996 : _GEN_8480; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8482 = 12'h7cd == _T_6[11:0] ? ram_1997 : _GEN_8481; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8483 = 12'h7ce == _T_6[11:0] ? ram_1998 : _GEN_8482; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8484 = 12'h7cf == _T_6[11:0] ? ram_1999 : _GEN_8483; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8485 = 12'h7d0 == _T_6[11:0] ? ram_2000 : _GEN_8484; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8486 = 12'h7d1 == _T_6[11:0] ? ram_2001 : _GEN_8485; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8487 = 12'h7d2 == _T_6[11:0] ? ram_2002 : _GEN_8486; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8488 = 12'h7d3 == _T_6[11:0] ? ram_2003 : _GEN_8487; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8489 = 12'h7d4 == _T_6[11:0] ? ram_2004 : _GEN_8488; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8490 = 12'h7d5 == _T_6[11:0] ? ram_2005 : _GEN_8489; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8491 = 12'h7d6 == _T_6[11:0] ? ram_2006 : _GEN_8490; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8492 = 12'h7d7 == _T_6[11:0] ? ram_2007 : _GEN_8491; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8493 = 12'h7d8 == _T_6[11:0] ? ram_2008 : _GEN_8492; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8494 = 12'h7d9 == _T_6[11:0] ? ram_2009 : _GEN_8493; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8495 = 12'h7da == _T_6[11:0] ? ram_2010 : _GEN_8494; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8496 = 12'h7db == _T_6[11:0] ? ram_2011 : _GEN_8495; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8497 = 12'h7dc == _T_6[11:0] ? ram_2012 : _GEN_8496; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8498 = 12'h7dd == _T_6[11:0] ? ram_2013 : _GEN_8497; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8499 = 12'h7de == _T_6[11:0] ? ram_2014 : _GEN_8498; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8500 = 12'h7df == _T_6[11:0] ? ram_2015 : _GEN_8499; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8501 = 12'h7e0 == _T_6[11:0] ? ram_2016 : _GEN_8500; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8502 = 12'h7e1 == _T_6[11:0] ? ram_2017 : _GEN_8501; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8503 = 12'h7e2 == _T_6[11:0] ? ram_2018 : _GEN_8502; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8504 = 12'h7e3 == _T_6[11:0] ? ram_2019 : _GEN_8503; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8505 = 12'h7e4 == _T_6[11:0] ? ram_2020 : _GEN_8504; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8506 = 12'h7e5 == _T_6[11:0] ? ram_2021 : _GEN_8505; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8507 = 12'h7e6 == _T_6[11:0] ? ram_2022 : _GEN_8506; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8508 = 12'h7e7 == _T_6[11:0] ? ram_2023 : _GEN_8507; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8509 = 12'h7e8 == _T_6[11:0] ? ram_2024 : _GEN_8508; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8510 = 12'h7e9 == _T_6[11:0] ? ram_2025 : _GEN_8509; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8511 = 12'h7ea == _T_6[11:0] ? ram_2026 : _GEN_8510; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8512 = 12'h7eb == _T_6[11:0] ? ram_2027 : _GEN_8511; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8513 = 12'h7ec == _T_6[11:0] ? ram_2028 : _GEN_8512; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8514 = 12'h7ed == _T_6[11:0] ? ram_2029 : _GEN_8513; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8515 = 12'h7ee == _T_6[11:0] ? ram_2030 : _GEN_8514; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8516 = 12'h7ef == _T_6[11:0] ? ram_2031 : _GEN_8515; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8517 = 12'h7f0 == _T_6[11:0] ? ram_2032 : _GEN_8516; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8518 = 12'h7f1 == _T_6[11:0] ? ram_2033 : _GEN_8517; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8519 = 12'h7f2 == _T_6[11:0] ? ram_2034 : _GEN_8518; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8520 = 12'h7f3 == _T_6[11:0] ? ram_2035 : _GEN_8519; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8521 = 12'h7f4 == _T_6[11:0] ? ram_2036 : _GEN_8520; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8522 = 12'h7f5 == _T_6[11:0] ? ram_2037 : _GEN_8521; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8523 = 12'h7f6 == _T_6[11:0] ? ram_2038 : _GEN_8522; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8524 = 12'h7f7 == _T_6[11:0] ? ram_2039 : _GEN_8523; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8525 = 12'h7f8 == _T_6[11:0] ? ram_2040 : _GEN_8524; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8526 = 12'h7f9 == _T_6[11:0] ? ram_2041 : _GEN_8525; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8527 = 12'h7fa == _T_6[11:0] ? ram_2042 : _GEN_8526; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8528 = 12'h7fb == _T_6[11:0] ? ram_2043 : _GEN_8527; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8529 = 12'h7fc == _T_6[11:0] ? ram_2044 : _GEN_8528; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8530 = 12'h7fd == _T_6[11:0] ? ram_2045 : _GEN_8529; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8531 = 12'h7fe == _T_6[11:0] ? ram_2046 : _GEN_8530; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8532 = 12'h7ff == _T_6[11:0] ? ram_2047 : _GEN_8531; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8533 = 12'h800 == _T_6[11:0] ? ram_2048 : _GEN_8532; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8534 = 12'h801 == _T_6[11:0] ? ram_2049 : _GEN_8533; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8535 = 12'h802 == _T_6[11:0] ? ram_2050 : _GEN_8534; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8536 = 12'h803 == _T_6[11:0] ? ram_2051 : _GEN_8535; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8537 = 12'h804 == _T_6[11:0] ? ram_2052 : _GEN_8536; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8538 = 12'h805 == _T_6[11:0] ? ram_2053 : _GEN_8537; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8539 = 12'h806 == _T_6[11:0] ? ram_2054 : _GEN_8538; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8540 = 12'h807 == _T_6[11:0] ? ram_2055 : _GEN_8539; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8541 = 12'h808 == _T_6[11:0] ? ram_2056 : _GEN_8540; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8542 = 12'h809 == _T_6[11:0] ? ram_2057 : _GEN_8541; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8543 = 12'h80a == _T_6[11:0] ? ram_2058 : _GEN_8542; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8544 = 12'h80b == _T_6[11:0] ? ram_2059 : _GEN_8543; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8545 = 12'h80c == _T_6[11:0] ? ram_2060 : _GEN_8544; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8546 = 12'h80d == _T_6[11:0] ? ram_2061 : _GEN_8545; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8547 = 12'h80e == _T_6[11:0] ? ram_2062 : _GEN_8546; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8548 = 12'h80f == _T_6[11:0] ? ram_2063 : _GEN_8547; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8549 = 12'h810 == _T_6[11:0] ? ram_2064 : _GEN_8548; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8550 = 12'h811 == _T_6[11:0] ? ram_2065 : _GEN_8549; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8551 = 12'h812 == _T_6[11:0] ? ram_2066 : _GEN_8550; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8552 = 12'h813 == _T_6[11:0] ? ram_2067 : _GEN_8551; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8553 = 12'h814 == _T_6[11:0] ? ram_2068 : _GEN_8552; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8554 = 12'h815 == _T_6[11:0] ? ram_2069 : _GEN_8553; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8555 = 12'h816 == _T_6[11:0] ? ram_2070 : _GEN_8554; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8556 = 12'h817 == _T_6[11:0] ? ram_2071 : _GEN_8555; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8557 = 12'h818 == _T_6[11:0] ? ram_2072 : _GEN_8556; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8558 = 12'h819 == _T_6[11:0] ? ram_2073 : _GEN_8557; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8559 = 12'h81a == _T_6[11:0] ? ram_2074 : _GEN_8558; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8560 = 12'h81b == _T_6[11:0] ? ram_2075 : _GEN_8559; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8561 = 12'h81c == _T_6[11:0] ? ram_2076 : _GEN_8560; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8562 = 12'h81d == _T_6[11:0] ? ram_2077 : _GEN_8561; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8563 = 12'h81e == _T_6[11:0] ? ram_2078 : _GEN_8562; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8564 = 12'h81f == _T_6[11:0] ? ram_2079 : _GEN_8563; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8565 = 12'h820 == _T_6[11:0] ? ram_2080 : _GEN_8564; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8566 = 12'h821 == _T_6[11:0] ? ram_2081 : _GEN_8565; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8567 = 12'h822 == _T_6[11:0] ? ram_2082 : _GEN_8566; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8568 = 12'h823 == _T_6[11:0] ? ram_2083 : _GEN_8567; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8569 = 12'h824 == _T_6[11:0] ? ram_2084 : _GEN_8568; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8570 = 12'h825 == _T_6[11:0] ? ram_2085 : _GEN_8569; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8571 = 12'h826 == _T_6[11:0] ? ram_2086 : _GEN_8570; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8572 = 12'h827 == _T_6[11:0] ? ram_2087 : _GEN_8571; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8573 = 12'h828 == _T_6[11:0] ? ram_2088 : _GEN_8572; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8574 = 12'h829 == _T_6[11:0] ? ram_2089 : _GEN_8573; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8575 = 12'h82a == _T_6[11:0] ? ram_2090 : _GEN_8574; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8576 = 12'h82b == _T_6[11:0] ? ram_2091 : _GEN_8575; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8577 = 12'h82c == _T_6[11:0] ? ram_2092 : _GEN_8576; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8578 = 12'h82d == _T_6[11:0] ? ram_2093 : _GEN_8577; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8579 = 12'h82e == _T_6[11:0] ? ram_2094 : _GEN_8578; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8580 = 12'h82f == _T_6[11:0] ? ram_2095 : _GEN_8579; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8581 = 12'h830 == _T_6[11:0] ? ram_2096 : _GEN_8580; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8582 = 12'h831 == _T_6[11:0] ? ram_2097 : _GEN_8581; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8583 = 12'h832 == _T_6[11:0] ? ram_2098 : _GEN_8582; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8584 = 12'h833 == _T_6[11:0] ? ram_2099 : _GEN_8583; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8585 = 12'h834 == _T_6[11:0] ? ram_2100 : _GEN_8584; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8586 = 12'h835 == _T_6[11:0] ? ram_2101 : _GEN_8585; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8587 = 12'h836 == _T_6[11:0] ? ram_2102 : _GEN_8586; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8588 = 12'h837 == _T_6[11:0] ? ram_2103 : _GEN_8587; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8589 = 12'h838 == _T_6[11:0] ? ram_2104 : _GEN_8588; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8590 = 12'h839 == _T_6[11:0] ? ram_2105 : _GEN_8589; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8591 = 12'h83a == _T_6[11:0] ? ram_2106 : _GEN_8590; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8592 = 12'h83b == _T_6[11:0] ? ram_2107 : _GEN_8591; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8593 = 12'h83c == _T_6[11:0] ? ram_2108 : _GEN_8592; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8594 = 12'h83d == _T_6[11:0] ? ram_2109 : _GEN_8593; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8595 = 12'h83e == _T_6[11:0] ? ram_2110 : _GEN_8594; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8596 = 12'h83f == _T_6[11:0] ? ram_2111 : _GEN_8595; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8597 = 12'h840 == _T_6[11:0] ? ram_2112 : _GEN_8596; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8598 = 12'h841 == _T_6[11:0] ? ram_2113 : _GEN_8597; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8599 = 12'h842 == _T_6[11:0] ? ram_2114 : _GEN_8598; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8600 = 12'h843 == _T_6[11:0] ? ram_2115 : _GEN_8599; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8601 = 12'h844 == _T_6[11:0] ? ram_2116 : _GEN_8600; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8602 = 12'h845 == _T_6[11:0] ? ram_2117 : _GEN_8601; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8603 = 12'h846 == _T_6[11:0] ? ram_2118 : _GEN_8602; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8604 = 12'h847 == _T_6[11:0] ? ram_2119 : _GEN_8603; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8605 = 12'h848 == _T_6[11:0] ? ram_2120 : _GEN_8604; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8606 = 12'h849 == _T_6[11:0] ? ram_2121 : _GEN_8605; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8607 = 12'h84a == _T_6[11:0] ? ram_2122 : _GEN_8606; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8608 = 12'h84b == _T_6[11:0] ? ram_2123 : _GEN_8607; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8609 = 12'h84c == _T_6[11:0] ? ram_2124 : _GEN_8608; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8610 = 12'h84d == _T_6[11:0] ? ram_2125 : _GEN_8609; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8611 = 12'h84e == _T_6[11:0] ? ram_2126 : _GEN_8610; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8612 = 12'h84f == _T_6[11:0] ? ram_2127 : _GEN_8611; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8613 = 12'h850 == _T_6[11:0] ? ram_2128 : _GEN_8612; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8614 = 12'h851 == _T_6[11:0] ? ram_2129 : _GEN_8613; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8615 = 12'h852 == _T_6[11:0] ? ram_2130 : _GEN_8614; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8616 = 12'h853 == _T_6[11:0] ? ram_2131 : _GEN_8615; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8617 = 12'h854 == _T_6[11:0] ? ram_2132 : _GEN_8616; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8618 = 12'h855 == _T_6[11:0] ? ram_2133 : _GEN_8617; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8619 = 12'h856 == _T_6[11:0] ? ram_2134 : _GEN_8618; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8620 = 12'h857 == _T_6[11:0] ? ram_2135 : _GEN_8619; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8621 = 12'h858 == _T_6[11:0] ? ram_2136 : _GEN_8620; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8622 = 12'h859 == _T_6[11:0] ? ram_2137 : _GEN_8621; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8623 = 12'h85a == _T_6[11:0] ? ram_2138 : _GEN_8622; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8624 = 12'h85b == _T_6[11:0] ? ram_2139 : _GEN_8623; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8625 = 12'h85c == _T_6[11:0] ? ram_2140 : _GEN_8624; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8626 = 12'h85d == _T_6[11:0] ? ram_2141 : _GEN_8625; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8627 = 12'h85e == _T_6[11:0] ? ram_2142 : _GEN_8626; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8628 = 12'h85f == _T_6[11:0] ? ram_2143 : _GEN_8627; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8629 = 12'h860 == _T_6[11:0] ? ram_2144 : _GEN_8628; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8630 = 12'h861 == _T_6[11:0] ? ram_2145 : _GEN_8629; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8631 = 12'h862 == _T_6[11:0] ? ram_2146 : _GEN_8630; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8632 = 12'h863 == _T_6[11:0] ? ram_2147 : _GEN_8631; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8633 = 12'h864 == _T_6[11:0] ? ram_2148 : _GEN_8632; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8634 = 12'h865 == _T_6[11:0] ? ram_2149 : _GEN_8633; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8635 = 12'h866 == _T_6[11:0] ? ram_2150 : _GEN_8634; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8636 = 12'h867 == _T_6[11:0] ? ram_2151 : _GEN_8635; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8637 = 12'h868 == _T_6[11:0] ? ram_2152 : _GEN_8636; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8638 = 12'h869 == _T_6[11:0] ? ram_2153 : _GEN_8637; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8639 = 12'h86a == _T_6[11:0] ? ram_2154 : _GEN_8638; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8640 = 12'h86b == _T_6[11:0] ? ram_2155 : _GEN_8639; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8641 = 12'h86c == _T_6[11:0] ? ram_2156 : _GEN_8640; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8642 = 12'h86d == _T_6[11:0] ? ram_2157 : _GEN_8641; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8643 = 12'h86e == _T_6[11:0] ? ram_2158 : _GEN_8642; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8644 = 12'h86f == _T_6[11:0] ? ram_2159 : _GEN_8643; // @[vga.scala 29:65 vga.scala 29:65]
  wire [7:0] _GEN_8645 = 12'h870 == _T_6[11:0] ? ram_2160 : _GEN_8644; // @[vga.scala 29:65 vga.scala 29:65]
  wire [11:0] _T_8 = {_GEN_8645, 4'h0}; // @[vga.scala 29:65]
  wire [8:0] _GEN_1 = io_v_addr % 9'h10; // @[vga.scala 29:79]
  wire [4:0] _T_9 = _GEN_1[4:0]; // @[vga.scala 29:79]
  wire [11:0] _GEN_10555 = {{7'd0}, _T_9}; // @[vga.scala 29:69]
  wire [9:0] _GEN_2 = io_h_addr % 10'h9; // @[vga.scala 29:95]
  wire [3:0] _T_12 = _GEN_2[3:0]; // @[vga.scala 29:95]
  wire [11:0] _T_13 = vga_mem_MPORT_data >> _T_12; // @[vga.scala 29:85]
  assign vga_mem_MPORT_addr = vga_mem_MPORT_addr_pipe_0;
  assign vga_mem_MPORT_data = vga_mem[vga_mem_MPORT_addr]; // @[vga.scala 16:30]
  assign io_vga_data = rdwrPort; // @[vga.scala 35:16]
  always @(posedge clock) begin
    vga_mem_MPORT_addr_pipe_0 <= _T_8 + _GEN_10555;
    if (reset) begin // @[vga.scala 13:27]
      rdwrPort <= 24'h0; // @[vga.scala 13:27]
    end else if (_T_13[0]) begin // @[vga.scala 29:107]
      rdwrPort <= 24'hffffff; // @[vga.scala 30:17]
    end else begin
      rdwrPort <= 24'h0; // @[vga.scala 32:17]
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_0 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h0 == index) begin // @[vga.scala 25:23]
          ram_0 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1 == index) begin // @[vga.scala 25:23]
          ram_1 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2 == index) begin // @[vga.scala 25:23]
          ram_2 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_3 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3 == index) begin // @[vga.scala 25:23]
          ram_3 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_4 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4 == index) begin // @[vga.scala 25:23]
          ram_4 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_5 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5 == index) begin // @[vga.scala 25:23]
          ram_5 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_6 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6 == index) begin // @[vga.scala 25:23]
          ram_6 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_7 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7 == index) begin // @[vga.scala 25:23]
          ram_7 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_8 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8 == index) begin // @[vga.scala 25:23]
          ram_8 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_9 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9 == index) begin // @[vga.scala 25:23]
          ram_9 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_10 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha == index) begin // @[vga.scala 25:23]
          ram_10 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_11 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb == index) begin // @[vga.scala 25:23]
          ram_11 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_12 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc == index) begin // @[vga.scala 25:23]
          ram_12 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_13 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd == index) begin // @[vga.scala 25:23]
          ram_13 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_14 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he == index) begin // @[vga.scala 25:23]
          ram_14 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_15 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf == index) begin // @[vga.scala 25:23]
          ram_15 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_16 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h10 == index) begin // @[vga.scala 25:23]
          ram_16 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_17 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h11 == index) begin // @[vga.scala 25:23]
          ram_17 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_18 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h12 == index) begin // @[vga.scala 25:23]
          ram_18 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_19 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h13 == index) begin // @[vga.scala 25:23]
          ram_19 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_20 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h14 == index) begin // @[vga.scala 25:23]
          ram_20 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_21 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h15 == index) begin // @[vga.scala 25:23]
          ram_21 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_22 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h16 == index) begin // @[vga.scala 25:23]
          ram_22 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_23 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h17 == index) begin // @[vga.scala 25:23]
          ram_23 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_24 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h18 == index) begin // @[vga.scala 25:23]
          ram_24 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_25 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h19 == index) begin // @[vga.scala 25:23]
          ram_25 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_26 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1a == index) begin // @[vga.scala 25:23]
          ram_26 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_27 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1b == index) begin // @[vga.scala 25:23]
          ram_27 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_28 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1c == index) begin // @[vga.scala 25:23]
          ram_28 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_29 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1d == index) begin // @[vga.scala 25:23]
          ram_29 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_30 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1e == index) begin // @[vga.scala 25:23]
          ram_30 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_31 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h1f == index) begin // @[vga.scala 25:23]
          ram_31 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_32 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h20 == index) begin // @[vga.scala 25:23]
          ram_32 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_33 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h21 == index) begin // @[vga.scala 25:23]
          ram_33 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_34 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h22 == index) begin // @[vga.scala 25:23]
          ram_34 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_35 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h23 == index) begin // @[vga.scala 25:23]
          ram_35 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_36 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h24 == index) begin // @[vga.scala 25:23]
          ram_36 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_37 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h25 == index) begin // @[vga.scala 25:23]
          ram_37 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_38 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h26 == index) begin // @[vga.scala 25:23]
          ram_38 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_39 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h27 == index) begin // @[vga.scala 25:23]
          ram_39 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_40 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h28 == index) begin // @[vga.scala 25:23]
          ram_40 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_41 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h29 == index) begin // @[vga.scala 25:23]
          ram_41 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_42 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2a == index) begin // @[vga.scala 25:23]
          ram_42 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_43 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2b == index) begin // @[vga.scala 25:23]
          ram_43 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_44 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2c == index) begin // @[vga.scala 25:23]
          ram_44 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_45 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2d == index) begin // @[vga.scala 25:23]
          ram_45 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_46 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2e == index) begin // @[vga.scala 25:23]
          ram_46 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_47 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h2f == index) begin // @[vga.scala 25:23]
          ram_47 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_48 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h30 == index) begin // @[vga.scala 25:23]
          ram_48 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_49 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h31 == index) begin // @[vga.scala 25:23]
          ram_49 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_50 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h32 == index) begin // @[vga.scala 25:23]
          ram_50 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_51 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h33 == index) begin // @[vga.scala 25:23]
          ram_51 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_52 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h34 == index) begin // @[vga.scala 25:23]
          ram_52 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_53 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h35 == index) begin // @[vga.scala 25:23]
          ram_53 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_54 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h36 == index) begin // @[vga.scala 25:23]
          ram_54 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_55 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h37 == index) begin // @[vga.scala 25:23]
          ram_55 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_56 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h38 == index) begin // @[vga.scala 25:23]
          ram_56 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_57 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h39 == index) begin // @[vga.scala 25:23]
          ram_57 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_58 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3a == index) begin // @[vga.scala 25:23]
          ram_58 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_59 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3b == index) begin // @[vga.scala 25:23]
          ram_59 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_60 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3c == index) begin // @[vga.scala 25:23]
          ram_60 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_61 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3d == index) begin // @[vga.scala 25:23]
          ram_61 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_62 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3e == index) begin // @[vga.scala 25:23]
          ram_62 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_63 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h3f == index) begin // @[vga.scala 25:23]
          ram_63 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_64 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h40 == index) begin // @[vga.scala 25:23]
          ram_64 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_65 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h41 == index) begin // @[vga.scala 25:23]
          ram_65 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_66 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h42 == index) begin // @[vga.scala 25:23]
          ram_66 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_67 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h43 == index) begin // @[vga.scala 25:23]
          ram_67 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_68 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h44 == index) begin // @[vga.scala 25:23]
          ram_68 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_69 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h45 == index) begin // @[vga.scala 25:23]
          ram_69 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_70 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h46 == index) begin // @[vga.scala 25:23]
          ram_70 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_71 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h47 == index) begin // @[vga.scala 25:23]
          ram_71 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_72 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h48 == index) begin // @[vga.scala 25:23]
          ram_72 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_73 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h49 == index) begin // @[vga.scala 25:23]
          ram_73 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_74 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4a == index) begin // @[vga.scala 25:23]
          ram_74 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_75 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4b == index) begin // @[vga.scala 25:23]
          ram_75 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_76 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4c == index) begin // @[vga.scala 25:23]
          ram_76 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_77 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4d == index) begin // @[vga.scala 25:23]
          ram_77 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_78 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4e == index) begin // @[vga.scala 25:23]
          ram_78 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_79 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h4f == index) begin // @[vga.scala 25:23]
          ram_79 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_80 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h50 == index) begin // @[vga.scala 25:23]
          ram_80 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_81 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h51 == index) begin // @[vga.scala 25:23]
          ram_81 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_82 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h52 == index) begin // @[vga.scala 25:23]
          ram_82 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_83 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h53 == index) begin // @[vga.scala 25:23]
          ram_83 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_84 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h54 == index) begin // @[vga.scala 25:23]
          ram_84 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_85 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h55 == index) begin // @[vga.scala 25:23]
          ram_85 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_86 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h56 == index) begin // @[vga.scala 25:23]
          ram_86 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_87 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h57 == index) begin // @[vga.scala 25:23]
          ram_87 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_88 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h58 == index) begin // @[vga.scala 25:23]
          ram_88 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_89 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h59 == index) begin // @[vga.scala 25:23]
          ram_89 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_90 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5a == index) begin // @[vga.scala 25:23]
          ram_90 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_91 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5b == index) begin // @[vga.scala 25:23]
          ram_91 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_92 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5c == index) begin // @[vga.scala 25:23]
          ram_92 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_93 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5d == index) begin // @[vga.scala 25:23]
          ram_93 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_94 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5e == index) begin // @[vga.scala 25:23]
          ram_94 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_95 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h5f == index) begin // @[vga.scala 25:23]
          ram_95 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_96 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h60 == index) begin // @[vga.scala 25:23]
          ram_96 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_97 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h61 == index) begin // @[vga.scala 25:23]
          ram_97 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_98 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h62 == index) begin // @[vga.scala 25:23]
          ram_98 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_99 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h63 == index) begin // @[vga.scala 25:23]
          ram_99 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_100 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h64 == index) begin // @[vga.scala 25:23]
          ram_100 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_101 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h65 == index) begin // @[vga.scala 25:23]
          ram_101 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_102 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h66 == index) begin // @[vga.scala 25:23]
          ram_102 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_103 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h67 == index) begin // @[vga.scala 25:23]
          ram_103 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_104 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h68 == index) begin // @[vga.scala 25:23]
          ram_104 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_105 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h69 == index) begin // @[vga.scala 25:23]
          ram_105 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_106 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6a == index) begin // @[vga.scala 25:23]
          ram_106 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_107 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6b == index) begin // @[vga.scala 25:23]
          ram_107 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_108 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6c == index) begin // @[vga.scala 25:23]
          ram_108 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_109 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6d == index) begin // @[vga.scala 25:23]
          ram_109 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_110 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6e == index) begin // @[vga.scala 25:23]
          ram_110 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_111 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h6f == index) begin // @[vga.scala 25:23]
          ram_111 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_112 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h70 == index) begin // @[vga.scala 25:23]
          ram_112 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_113 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h71 == index) begin // @[vga.scala 25:23]
          ram_113 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_114 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h72 == index) begin // @[vga.scala 25:23]
          ram_114 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_115 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h73 == index) begin // @[vga.scala 25:23]
          ram_115 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_116 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h74 == index) begin // @[vga.scala 25:23]
          ram_116 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_117 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h75 == index) begin // @[vga.scala 25:23]
          ram_117 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_118 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h76 == index) begin // @[vga.scala 25:23]
          ram_118 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_119 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h77 == index) begin // @[vga.scala 25:23]
          ram_119 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_120 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h78 == index) begin // @[vga.scala 25:23]
          ram_120 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_121 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h79 == index) begin // @[vga.scala 25:23]
          ram_121 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_122 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7a == index) begin // @[vga.scala 25:23]
          ram_122 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_123 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7b == index) begin // @[vga.scala 25:23]
          ram_123 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_124 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7c == index) begin // @[vga.scala 25:23]
          ram_124 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_125 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7d == index) begin // @[vga.scala 25:23]
          ram_125 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_126 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7e == index) begin // @[vga.scala 25:23]
          ram_126 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_127 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h7f == index) begin // @[vga.scala 25:23]
          ram_127 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_128 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h80 == index) begin // @[vga.scala 25:23]
          ram_128 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_129 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h81 == index) begin // @[vga.scala 25:23]
          ram_129 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_130 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h82 == index) begin // @[vga.scala 25:23]
          ram_130 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_131 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h83 == index) begin // @[vga.scala 25:23]
          ram_131 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_132 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h84 == index) begin // @[vga.scala 25:23]
          ram_132 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_133 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h85 == index) begin // @[vga.scala 25:23]
          ram_133 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_134 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h86 == index) begin // @[vga.scala 25:23]
          ram_134 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_135 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h87 == index) begin // @[vga.scala 25:23]
          ram_135 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_136 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h88 == index) begin // @[vga.scala 25:23]
          ram_136 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_137 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h89 == index) begin // @[vga.scala 25:23]
          ram_137 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_138 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8a == index) begin // @[vga.scala 25:23]
          ram_138 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_139 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8b == index) begin // @[vga.scala 25:23]
          ram_139 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_140 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8c == index) begin // @[vga.scala 25:23]
          ram_140 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_141 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8d == index) begin // @[vga.scala 25:23]
          ram_141 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_142 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8e == index) begin // @[vga.scala 25:23]
          ram_142 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_143 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h8f == index) begin // @[vga.scala 25:23]
          ram_143 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_144 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h90 == index) begin // @[vga.scala 25:23]
          ram_144 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_145 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h91 == index) begin // @[vga.scala 25:23]
          ram_145 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_146 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h92 == index) begin // @[vga.scala 25:23]
          ram_146 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_147 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h93 == index) begin // @[vga.scala 25:23]
          ram_147 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_148 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h94 == index) begin // @[vga.scala 25:23]
          ram_148 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_149 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h95 == index) begin // @[vga.scala 25:23]
          ram_149 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_150 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h96 == index) begin // @[vga.scala 25:23]
          ram_150 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_151 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h97 == index) begin // @[vga.scala 25:23]
          ram_151 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_152 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h98 == index) begin // @[vga.scala 25:23]
          ram_152 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_153 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h99 == index) begin // @[vga.scala 25:23]
          ram_153 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_154 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9a == index) begin // @[vga.scala 25:23]
          ram_154 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_155 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9b == index) begin // @[vga.scala 25:23]
          ram_155 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_156 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9c == index) begin // @[vga.scala 25:23]
          ram_156 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_157 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9d == index) begin // @[vga.scala 25:23]
          ram_157 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_158 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9e == index) begin // @[vga.scala 25:23]
          ram_158 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_159 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'h9f == index) begin // @[vga.scala 25:23]
          ram_159 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_160 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha0 == index) begin // @[vga.scala 25:23]
          ram_160 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_161 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha1 == index) begin // @[vga.scala 25:23]
          ram_161 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_162 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha2 == index) begin // @[vga.scala 25:23]
          ram_162 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_163 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha3 == index) begin // @[vga.scala 25:23]
          ram_163 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_164 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha4 == index) begin // @[vga.scala 25:23]
          ram_164 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_165 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha5 == index) begin // @[vga.scala 25:23]
          ram_165 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_166 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha6 == index) begin // @[vga.scala 25:23]
          ram_166 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_167 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha7 == index) begin // @[vga.scala 25:23]
          ram_167 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_168 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha8 == index) begin // @[vga.scala 25:23]
          ram_168 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_169 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'ha9 == index) begin // @[vga.scala 25:23]
          ram_169 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_170 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'haa == index) begin // @[vga.scala 25:23]
          ram_170 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_171 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hab == index) begin // @[vga.scala 25:23]
          ram_171 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_172 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hac == index) begin // @[vga.scala 25:23]
          ram_172 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_173 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'had == index) begin // @[vga.scala 25:23]
          ram_173 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_174 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hae == index) begin // @[vga.scala 25:23]
          ram_174 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_175 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'haf == index) begin // @[vga.scala 25:23]
          ram_175 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_176 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb0 == index) begin // @[vga.scala 25:23]
          ram_176 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_177 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb1 == index) begin // @[vga.scala 25:23]
          ram_177 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_178 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb2 == index) begin // @[vga.scala 25:23]
          ram_178 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_179 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb3 == index) begin // @[vga.scala 25:23]
          ram_179 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_180 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb4 == index) begin // @[vga.scala 25:23]
          ram_180 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_181 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb5 == index) begin // @[vga.scala 25:23]
          ram_181 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_182 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb6 == index) begin // @[vga.scala 25:23]
          ram_182 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_183 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb7 == index) begin // @[vga.scala 25:23]
          ram_183 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_184 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb8 == index) begin // @[vga.scala 25:23]
          ram_184 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_185 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hb9 == index) begin // @[vga.scala 25:23]
          ram_185 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_186 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hba == index) begin // @[vga.scala 25:23]
          ram_186 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_187 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hbb == index) begin // @[vga.scala 25:23]
          ram_187 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_188 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hbc == index) begin // @[vga.scala 25:23]
          ram_188 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_189 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hbd == index) begin // @[vga.scala 25:23]
          ram_189 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_190 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hbe == index) begin // @[vga.scala 25:23]
          ram_190 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_191 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hbf == index) begin // @[vga.scala 25:23]
          ram_191 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_192 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc0 == index) begin // @[vga.scala 25:23]
          ram_192 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_193 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc1 == index) begin // @[vga.scala 25:23]
          ram_193 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_194 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc2 == index) begin // @[vga.scala 25:23]
          ram_194 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_195 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc3 == index) begin // @[vga.scala 25:23]
          ram_195 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_196 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc4 == index) begin // @[vga.scala 25:23]
          ram_196 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_197 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc5 == index) begin // @[vga.scala 25:23]
          ram_197 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_198 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc6 == index) begin // @[vga.scala 25:23]
          ram_198 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_199 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc7 == index) begin // @[vga.scala 25:23]
          ram_199 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_200 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc8 == index) begin // @[vga.scala 25:23]
          ram_200 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_201 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hc9 == index) begin // @[vga.scala 25:23]
          ram_201 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_202 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hca == index) begin // @[vga.scala 25:23]
          ram_202 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_203 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hcb == index) begin // @[vga.scala 25:23]
          ram_203 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_204 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hcc == index) begin // @[vga.scala 25:23]
          ram_204 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_205 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hcd == index) begin // @[vga.scala 25:23]
          ram_205 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_206 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hce == index) begin // @[vga.scala 25:23]
          ram_206 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_207 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hcf == index) begin // @[vga.scala 25:23]
          ram_207 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_208 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd0 == index) begin // @[vga.scala 25:23]
          ram_208 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_209 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd1 == index) begin // @[vga.scala 25:23]
          ram_209 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_210 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd2 == index) begin // @[vga.scala 25:23]
          ram_210 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_211 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd3 == index) begin // @[vga.scala 25:23]
          ram_211 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_212 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd4 == index) begin // @[vga.scala 25:23]
          ram_212 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_213 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd5 == index) begin // @[vga.scala 25:23]
          ram_213 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_214 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd6 == index) begin // @[vga.scala 25:23]
          ram_214 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_215 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd7 == index) begin // @[vga.scala 25:23]
          ram_215 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_216 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd8 == index) begin // @[vga.scala 25:23]
          ram_216 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_217 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hd9 == index) begin // @[vga.scala 25:23]
          ram_217 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_218 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hda == index) begin // @[vga.scala 25:23]
          ram_218 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_219 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hdb == index) begin // @[vga.scala 25:23]
          ram_219 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_220 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hdc == index) begin // @[vga.scala 25:23]
          ram_220 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_221 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hdd == index) begin // @[vga.scala 25:23]
          ram_221 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_222 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hde == index) begin // @[vga.scala 25:23]
          ram_222 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_223 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hdf == index) begin // @[vga.scala 25:23]
          ram_223 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_224 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he0 == index) begin // @[vga.scala 25:23]
          ram_224 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_225 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he1 == index) begin // @[vga.scala 25:23]
          ram_225 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_226 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he2 == index) begin // @[vga.scala 25:23]
          ram_226 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_227 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he3 == index) begin // @[vga.scala 25:23]
          ram_227 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_228 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he4 == index) begin // @[vga.scala 25:23]
          ram_228 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_229 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he5 == index) begin // @[vga.scala 25:23]
          ram_229 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_230 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he6 == index) begin // @[vga.scala 25:23]
          ram_230 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_231 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he7 == index) begin // @[vga.scala 25:23]
          ram_231 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_232 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he8 == index) begin // @[vga.scala 25:23]
          ram_232 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_233 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'he9 == index) begin // @[vga.scala 25:23]
          ram_233 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_234 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hea == index) begin // @[vga.scala 25:23]
          ram_234 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_235 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'heb == index) begin // @[vga.scala 25:23]
          ram_235 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_236 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hec == index) begin // @[vga.scala 25:23]
          ram_236 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_237 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hed == index) begin // @[vga.scala 25:23]
          ram_237 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_238 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hee == index) begin // @[vga.scala 25:23]
          ram_238 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_239 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hef == index) begin // @[vga.scala 25:23]
          ram_239 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_240 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf0 == index) begin // @[vga.scala 25:23]
          ram_240 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_241 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf1 == index) begin // @[vga.scala 25:23]
          ram_241 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_242 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf2 == index) begin // @[vga.scala 25:23]
          ram_242 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_243 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf3 == index) begin // @[vga.scala 25:23]
          ram_243 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_244 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf4 == index) begin // @[vga.scala 25:23]
          ram_244 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_245 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf5 == index) begin // @[vga.scala 25:23]
          ram_245 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_246 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf6 == index) begin // @[vga.scala 25:23]
          ram_246 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_247 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf7 == index) begin // @[vga.scala 25:23]
          ram_247 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_248 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf8 == index) begin // @[vga.scala 25:23]
          ram_248 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_249 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hf9 == index) begin // @[vga.scala 25:23]
          ram_249 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_250 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hfa == index) begin // @[vga.scala 25:23]
          ram_250 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_251 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hfb == index) begin // @[vga.scala 25:23]
          ram_251 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_252 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hfc == index) begin // @[vga.scala 25:23]
          ram_252 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_253 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hfd == index) begin // @[vga.scala 25:23]
          ram_253 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_254 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hfe == index) begin // @[vga.scala 25:23]
          ram_254 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_255 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (8'hff == index) begin // @[vga.scala 25:23]
          ram_255 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_256 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h100 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_256 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_257 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h101 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_257 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_258 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h102 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_258 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_259 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h103 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_259 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_260 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h104 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_260 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_261 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h105 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_261 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_262 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h106 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_262 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_263 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h107 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_263 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_264 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h108 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_264 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_265 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h109 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_265 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_266 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_266 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_267 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_267 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_268 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_268 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_269 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_269 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_270 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_270 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_271 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h10f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_271 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_272 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h110 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_272 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_273 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h111 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_273 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_274 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h112 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_274 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_275 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h113 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_275 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_276 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h114 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_276 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_277 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h115 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_277 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_278 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h116 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_278 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_279 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h117 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_279 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_280 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h118 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_280 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_281 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h119 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_281 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_282 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_282 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_283 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_283 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_284 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_284 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_285 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_285 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_286 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_286 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_287 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h11f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_287 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_288 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h120 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_288 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_289 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h121 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_289 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_290 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h122 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_290 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_291 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h123 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_291 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_292 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h124 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_292 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_293 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h125 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_293 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_294 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h126 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_294 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_295 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h127 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_295 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_296 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h128 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_296 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_297 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h129 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_297 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_298 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_298 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_299 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_299 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_300 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_300 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_301 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_301 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_302 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_302 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_303 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h12f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_303 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_304 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h130 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_304 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_305 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h131 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_305 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_306 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h132 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_306 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_307 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h133 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_307 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_308 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h134 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_308 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_309 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h135 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_309 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_310 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h136 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_310 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_311 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h137 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_311 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_312 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h138 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_312 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_313 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h139 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_313 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_314 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_314 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_315 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_315 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_316 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_316 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_317 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_317 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_318 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_318 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_319 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h13f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_319 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_320 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h140 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_320 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_321 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h141 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_321 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_322 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h142 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_322 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_323 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h143 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_323 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_324 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h144 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_324 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_325 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h145 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_325 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_326 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h146 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_326 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_327 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h147 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_327 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_328 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h148 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_328 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_329 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h149 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_329 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_330 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_330 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_331 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_331 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_332 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_332 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_333 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_333 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_334 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_334 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_335 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h14f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_335 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_336 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h150 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_336 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_337 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h151 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_337 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_338 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h152 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_338 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_339 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h153 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_339 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_340 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h154 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_340 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_341 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h155 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_341 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_342 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h156 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_342 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_343 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h157 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_343 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_344 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h158 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_344 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_345 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h159 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_345 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_346 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_346 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_347 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_347 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_348 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_348 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_349 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_349 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_350 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_350 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_351 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h15f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_351 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_352 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h160 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_352 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_353 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h161 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_353 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_354 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h162 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_354 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_355 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h163 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_355 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_356 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h164 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_356 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_357 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h165 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_357 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_358 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h166 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_358 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_359 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h167 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_359 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_360 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h168 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_360 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_361 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h169 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_361 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_362 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_362 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_363 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_363 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_364 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_364 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_365 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_365 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_366 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_366 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_367 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h16f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_367 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_368 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h170 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_368 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_369 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h171 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_369 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_370 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h172 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_370 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_371 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h173 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_371 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_372 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h174 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_372 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_373 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h175 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_373 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_374 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h176 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_374 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_375 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h177 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_375 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_376 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h178 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_376 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_377 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h179 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_377 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_378 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_378 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_379 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_379 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_380 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_380 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_381 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_381 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_382 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_382 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_383 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h17f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_383 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_384 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h180 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_384 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_385 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h181 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_385 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_386 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h182 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_386 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_387 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h183 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_387 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_388 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h184 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_388 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_389 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h185 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_389 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_390 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h186 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_390 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_391 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h187 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_391 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_392 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h188 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_392 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_393 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h189 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_393 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_394 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_394 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_395 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_395 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_396 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_396 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_397 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_397 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_398 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_398 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_399 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h18f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_399 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_400 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h190 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_400 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_401 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h191 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_401 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_402 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h192 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_402 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_403 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h193 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_403 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_404 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h194 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_404 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_405 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h195 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_405 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_406 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h196 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_406 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_407 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h197 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_407 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_408 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h198 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_408 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_409 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h199 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_409 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_410 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19a == _GEN_8648) begin // @[vga.scala 25:23]
          ram_410 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_411 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19b == _GEN_8648) begin // @[vga.scala 25:23]
          ram_411 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_412 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19c == _GEN_8648) begin // @[vga.scala 25:23]
          ram_412 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_413 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19d == _GEN_8648) begin // @[vga.scala 25:23]
          ram_413 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_414 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19e == _GEN_8648) begin // @[vga.scala 25:23]
          ram_414 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_415 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h19f == _GEN_8648) begin // @[vga.scala 25:23]
          ram_415 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_416 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_416 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_417 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_417 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_418 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_418 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_419 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_419 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_420 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_420 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_421 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_421 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_422 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_422 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_423 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_423 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_424 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_424 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_425 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1a9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_425 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_426 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1aa == _GEN_8648) begin // @[vga.scala 25:23]
          ram_426 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_427 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ab == _GEN_8648) begin // @[vga.scala 25:23]
          ram_427 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_428 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ac == _GEN_8648) begin // @[vga.scala 25:23]
          ram_428 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_429 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ad == _GEN_8648) begin // @[vga.scala 25:23]
          ram_429 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_430 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ae == _GEN_8648) begin // @[vga.scala 25:23]
          ram_430 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_431 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1af == _GEN_8648) begin // @[vga.scala 25:23]
          ram_431 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_432 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_432 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_433 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_433 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_434 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_434 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_435 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_435 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_436 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_436 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_437 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_437 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_438 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_438 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_439 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_439 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_440 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_440 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_441 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1b9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_441 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_442 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ba == _GEN_8648) begin // @[vga.scala 25:23]
          ram_442 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_443 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1bb == _GEN_8648) begin // @[vga.scala 25:23]
          ram_443 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_444 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1bc == _GEN_8648) begin // @[vga.scala 25:23]
          ram_444 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_445 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1bd == _GEN_8648) begin // @[vga.scala 25:23]
          ram_445 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_446 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1be == _GEN_8648) begin // @[vga.scala 25:23]
          ram_446 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_447 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1bf == _GEN_8648) begin // @[vga.scala 25:23]
          ram_447 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_448 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_448 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_449 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_449 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_450 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_450 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_451 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_451 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_452 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_452 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_453 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_453 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_454 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_454 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_455 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_455 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_456 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_456 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_457 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1c9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_457 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_458 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ca == _GEN_8648) begin // @[vga.scala 25:23]
          ram_458 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_459 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1cb == _GEN_8648) begin // @[vga.scala 25:23]
          ram_459 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_460 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1cc == _GEN_8648) begin // @[vga.scala 25:23]
          ram_460 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_461 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1cd == _GEN_8648) begin // @[vga.scala 25:23]
          ram_461 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_462 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ce == _GEN_8648) begin // @[vga.scala 25:23]
          ram_462 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_463 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1cf == _GEN_8648) begin // @[vga.scala 25:23]
          ram_463 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_464 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_464 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_465 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_465 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_466 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_466 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_467 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_467 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_468 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_468 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_469 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_469 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_470 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_470 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_471 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_471 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_472 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_472 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_473 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1d9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_473 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_474 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1da == _GEN_8648) begin // @[vga.scala 25:23]
          ram_474 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_475 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1db == _GEN_8648) begin // @[vga.scala 25:23]
          ram_475 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_476 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1dc == _GEN_8648) begin // @[vga.scala 25:23]
          ram_476 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_477 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1dd == _GEN_8648) begin // @[vga.scala 25:23]
          ram_477 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_478 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1de == _GEN_8648) begin // @[vga.scala 25:23]
          ram_478 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_479 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1df == _GEN_8648) begin // @[vga.scala 25:23]
          ram_479 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_480 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_480 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_481 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_481 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_482 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_482 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_483 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_483 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_484 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_484 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_485 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_485 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_486 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_486 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_487 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_487 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_488 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_488 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_489 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1e9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_489 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_490 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ea == _GEN_8648) begin // @[vga.scala 25:23]
          ram_490 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_491 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1eb == _GEN_8648) begin // @[vga.scala 25:23]
          ram_491 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_492 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ec == _GEN_8648) begin // @[vga.scala 25:23]
          ram_492 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_493 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ed == _GEN_8648) begin // @[vga.scala 25:23]
          ram_493 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_494 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ee == _GEN_8648) begin // @[vga.scala 25:23]
          ram_494 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_495 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ef == _GEN_8648) begin // @[vga.scala 25:23]
          ram_495 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_496 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f0 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_496 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_497 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f1 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_497 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_498 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f2 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_498 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_499 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f3 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_499 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_500 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f4 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_500 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_501 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f5 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_501 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_502 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f6 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_502 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_503 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f7 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_503 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_504 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f8 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_504 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_505 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1f9 == _GEN_8648) begin // @[vga.scala 25:23]
          ram_505 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_506 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1fa == _GEN_8648) begin // @[vga.scala 25:23]
          ram_506 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_507 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1fb == _GEN_8648) begin // @[vga.scala 25:23]
          ram_507 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_508 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1fc == _GEN_8648) begin // @[vga.scala 25:23]
          ram_508 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_509 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1fd == _GEN_8648) begin // @[vga.scala 25:23]
          ram_509 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_510 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1fe == _GEN_8648) begin // @[vga.scala 25:23]
          ram_510 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_511 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (9'h1ff == _GEN_8648) begin // @[vga.scala 25:23]
          ram_511 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_512 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h200 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_512 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_513 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h201 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_513 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_514 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h202 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_514 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_515 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h203 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_515 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_516 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h204 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_516 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_517 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h205 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_517 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_518 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h206 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_518 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_519 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h207 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_519 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_520 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h208 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_520 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_521 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h209 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_521 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_522 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_522 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_523 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_523 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_524 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_524 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_525 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_525 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_526 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_526 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_527 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h20f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_527 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_528 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h210 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_528 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_529 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h211 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_529 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_530 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h212 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_530 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_531 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h213 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_531 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_532 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h214 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_532 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_533 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h215 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_533 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_534 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h216 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_534 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_535 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h217 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_535 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_536 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h218 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_536 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_537 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h219 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_537 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_538 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_538 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_539 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_539 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_540 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_540 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_541 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_541 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_542 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_542 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_543 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h21f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_543 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_544 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h220 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_544 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_545 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h221 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_545 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_546 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h222 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_546 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_547 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h223 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_547 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_548 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h224 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_548 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_549 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h225 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_549 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_550 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h226 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_550 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_551 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h227 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_551 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_552 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h228 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_552 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_553 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h229 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_553 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_554 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_554 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_555 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_555 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_556 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_556 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_557 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_557 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_558 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_558 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_559 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h22f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_559 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_560 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h230 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_560 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_561 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h231 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_561 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_562 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h232 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_562 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_563 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h233 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_563 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_564 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h234 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_564 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_565 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h235 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_565 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_566 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h236 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_566 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_567 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h237 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_567 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_568 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h238 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_568 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_569 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h239 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_569 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_570 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_570 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_571 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_571 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_572 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_572 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_573 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_573 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_574 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_574 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_575 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h23f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_575 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_576 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h240 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_576 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_577 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h241 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_577 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_578 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h242 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_578 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_579 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h243 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_579 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_580 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h244 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_580 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_581 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h245 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_581 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_582 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h246 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_582 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_583 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h247 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_583 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_584 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h248 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_584 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_585 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h249 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_585 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_586 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_586 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_587 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_587 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_588 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_588 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_589 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_589 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_590 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_590 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_591 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h24f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_591 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_592 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h250 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_592 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_593 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h251 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_593 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_594 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h252 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_594 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_595 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h253 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_595 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_596 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h254 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_596 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_597 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h255 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_597 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_598 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h256 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_598 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_599 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h257 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_599 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_600 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h258 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_600 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_601 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h259 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_601 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_602 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_602 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_603 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_603 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_604 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_604 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_605 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_605 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_606 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_606 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_607 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h25f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_607 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_608 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h260 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_608 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_609 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h261 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_609 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_610 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h262 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_610 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_611 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h263 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_611 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_612 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h264 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_612 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_613 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h265 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_613 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_614 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h266 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_614 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_615 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h267 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_615 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_616 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h268 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_616 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_617 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h269 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_617 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_618 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_618 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_619 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_619 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_620 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_620 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_621 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_621 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_622 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_622 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_623 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h26f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_623 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_624 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h270 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_624 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_625 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h271 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_625 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_626 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h272 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_626 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_627 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h273 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_627 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_628 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h274 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_628 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_629 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h275 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_629 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_630 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h276 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_630 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_631 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h277 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_631 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_632 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h278 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_632 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_633 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h279 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_633 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_634 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_634 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_635 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_635 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_636 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_636 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_637 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_637 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_638 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_638 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_639 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h27f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_639 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_640 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h280 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_640 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_641 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h281 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_641 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_642 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h282 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_642 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_643 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h283 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_643 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_644 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h284 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_644 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_645 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h285 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_645 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_646 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h286 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_646 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_647 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h287 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_647 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_648 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h288 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_648 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_649 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h289 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_649 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_650 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_650 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_651 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_651 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_652 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_652 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_653 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_653 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_654 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_654 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_655 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h28f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_655 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_656 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h290 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_656 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_657 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h291 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_657 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_658 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h292 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_658 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_659 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h293 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_659 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_660 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h294 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_660 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_661 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h295 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_661 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_662 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h296 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_662 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_663 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h297 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_663 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_664 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h298 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_664 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_665 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h299 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_665 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_666 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_666 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_667 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_667 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_668 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_668 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_669 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_669 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_670 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_670 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_671 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h29f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_671 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_672 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_672 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_673 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_673 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_674 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_674 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_675 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_675 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_676 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_676 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_677 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_677 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_678 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_678 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_679 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_679 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_680 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_680 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_681 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2a9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_681 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_682 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2aa == _GEN_8904) begin // @[vga.scala 25:23]
          ram_682 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_683 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ab == _GEN_8904) begin // @[vga.scala 25:23]
          ram_683 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_684 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ac == _GEN_8904) begin // @[vga.scala 25:23]
          ram_684 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_685 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ad == _GEN_8904) begin // @[vga.scala 25:23]
          ram_685 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_686 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ae == _GEN_8904) begin // @[vga.scala 25:23]
          ram_686 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_687 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2af == _GEN_8904) begin // @[vga.scala 25:23]
          ram_687 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_688 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_688 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_689 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_689 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_690 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_690 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_691 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_691 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_692 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_692 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_693 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_693 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_694 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_694 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_695 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_695 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_696 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_696 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_697 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2b9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_697 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_698 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ba == _GEN_8904) begin // @[vga.scala 25:23]
          ram_698 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_699 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2bb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_699 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_700 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2bc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_700 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_701 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2bd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_701 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_702 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2be == _GEN_8904) begin // @[vga.scala 25:23]
          ram_702 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_703 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2bf == _GEN_8904) begin // @[vga.scala 25:23]
          ram_703 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_704 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_704 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_705 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_705 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_706 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_706 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_707 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_707 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_708 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_708 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_709 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_709 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_710 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_710 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_711 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_711 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_712 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_712 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_713 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2c9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_713 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_714 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ca == _GEN_8904) begin // @[vga.scala 25:23]
          ram_714 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_715 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2cb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_715 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_716 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2cc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_716 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_717 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2cd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_717 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_718 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ce == _GEN_8904) begin // @[vga.scala 25:23]
          ram_718 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_719 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2cf == _GEN_8904) begin // @[vga.scala 25:23]
          ram_719 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_720 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_720 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_721 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_721 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_722 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_722 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_723 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_723 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_724 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_724 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_725 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_725 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_726 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_726 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_727 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_727 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_728 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_728 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_729 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2d9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_729 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_730 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2da == _GEN_8904) begin // @[vga.scala 25:23]
          ram_730 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_731 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2db == _GEN_8904) begin // @[vga.scala 25:23]
          ram_731 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_732 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2dc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_732 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_733 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2dd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_733 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_734 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2de == _GEN_8904) begin // @[vga.scala 25:23]
          ram_734 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_735 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2df == _GEN_8904) begin // @[vga.scala 25:23]
          ram_735 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_736 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_736 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_737 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_737 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_738 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_738 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_739 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_739 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_740 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_740 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_741 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_741 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_742 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_742 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_743 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_743 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_744 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_744 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_745 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2e9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_745 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_746 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ea == _GEN_8904) begin // @[vga.scala 25:23]
          ram_746 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_747 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2eb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_747 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_748 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ec == _GEN_8904) begin // @[vga.scala 25:23]
          ram_748 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_749 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ed == _GEN_8904) begin // @[vga.scala 25:23]
          ram_749 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_750 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ee == _GEN_8904) begin // @[vga.scala 25:23]
          ram_750 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_751 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ef == _GEN_8904) begin // @[vga.scala 25:23]
          ram_751 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_752 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_752 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_753 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_753 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_754 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_754 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_755 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_755 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_756 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_756 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_757 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_757 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_758 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_758 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_759 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_759 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_760 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_760 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_761 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2f9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_761 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_762 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2fa == _GEN_8904) begin // @[vga.scala 25:23]
          ram_762 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_763 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2fb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_763 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_764 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2fc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_764 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_765 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2fd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_765 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_766 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2fe == _GEN_8904) begin // @[vga.scala 25:23]
          ram_766 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_767 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h2ff == _GEN_8904) begin // @[vga.scala 25:23]
          ram_767 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_768 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h300 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_768 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_769 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h301 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_769 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_770 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h302 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_770 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_771 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h303 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_771 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_772 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h304 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_772 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_773 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h305 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_773 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_774 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h306 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_774 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_775 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h307 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_775 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_776 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h308 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_776 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_777 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h309 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_777 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_778 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_778 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_779 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_779 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_780 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_780 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_781 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_781 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_782 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_782 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_783 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h30f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_783 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_784 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h310 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_784 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_785 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h311 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_785 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_786 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h312 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_786 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_787 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h313 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_787 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_788 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h314 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_788 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_789 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h315 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_789 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_790 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h316 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_790 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_791 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h317 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_791 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_792 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h318 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_792 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_793 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h319 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_793 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_794 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_794 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_795 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_795 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_796 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_796 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_797 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_797 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_798 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_798 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_799 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h31f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_799 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_800 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h320 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_800 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_801 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h321 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_801 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_802 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h322 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_802 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_803 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h323 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_803 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_804 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h324 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_804 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_805 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h325 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_805 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_806 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h326 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_806 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_807 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h327 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_807 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_808 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h328 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_808 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_809 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h329 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_809 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_810 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_810 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_811 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_811 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_812 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_812 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_813 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_813 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_814 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_814 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_815 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h32f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_815 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_816 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h330 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_816 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_817 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h331 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_817 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_818 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h332 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_818 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_819 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h333 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_819 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_820 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h334 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_820 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_821 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h335 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_821 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_822 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h336 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_822 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_823 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h337 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_823 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_824 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h338 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_824 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_825 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h339 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_825 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_826 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_826 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_827 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_827 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_828 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_828 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_829 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_829 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_830 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_830 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_831 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h33f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_831 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_832 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h340 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_832 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_833 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h341 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_833 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_834 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h342 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_834 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_835 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h343 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_835 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_836 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h344 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_836 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_837 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h345 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_837 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_838 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h346 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_838 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_839 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h347 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_839 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_840 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h348 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_840 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_841 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h349 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_841 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_842 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_842 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_843 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_843 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_844 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_844 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_845 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_845 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_846 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_846 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_847 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h34f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_847 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_848 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h350 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_848 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_849 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h351 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_849 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_850 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h352 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_850 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_851 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h353 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_851 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_852 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h354 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_852 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_853 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h355 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_853 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_854 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h356 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_854 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_855 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h357 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_855 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_856 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h358 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_856 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_857 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h359 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_857 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_858 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_858 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_859 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_859 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_860 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_860 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_861 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_861 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_862 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_862 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_863 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h35f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_863 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_864 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h360 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_864 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_865 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h361 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_865 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_866 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h362 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_866 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_867 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h363 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_867 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_868 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h364 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_868 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_869 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h365 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_869 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_870 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h366 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_870 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_871 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h367 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_871 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_872 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h368 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_872 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_873 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h369 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_873 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_874 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_874 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_875 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_875 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_876 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_876 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_877 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_877 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_878 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_878 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_879 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h36f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_879 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_880 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h370 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_880 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_881 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h371 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_881 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_882 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h372 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_882 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_883 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h373 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_883 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_884 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h374 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_884 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_885 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h375 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_885 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_886 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h376 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_886 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_887 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h377 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_887 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_888 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h378 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_888 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_889 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h379 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_889 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_890 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_890 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_891 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_891 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_892 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_892 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_893 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_893 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_894 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_894 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_895 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h37f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_895 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_896 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h380 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_896 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_897 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h381 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_897 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_898 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h382 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_898 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_899 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h383 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_899 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_900 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h384 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_900 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_901 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h385 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_901 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_902 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h386 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_902 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_903 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h387 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_903 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_904 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h388 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_904 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_905 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h389 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_905 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_906 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_906 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_907 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_907 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_908 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_908 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_909 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_909 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_910 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_910 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_911 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h38f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_911 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_912 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h390 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_912 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_913 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h391 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_913 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_914 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h392 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_914 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_915 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h393 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_915 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_916 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h394 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_916 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_917 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h395 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_917 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_918 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h396 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_918 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_919 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h397 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_919 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_920 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h398 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_920 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_921 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h399 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_921 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_922 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39a == _GEN_8904) begin // @[vga.scala 25:23]
          ram_922 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_923 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39b == _GEN_8904) begin // @[vga.scala 25:23]
          ram_923 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_924 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39c == _GEN_8904) begin // @[vga.scala 25:23]
          ram_924 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_925 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39d == _GEN_8904) begin // @[vga.scala 25:23]
          ram_925 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_926 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39e == _GEN_8904) begin // @[vga.scala 25:23]
          ram_926 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_927 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h39f == _GEN_8904) begin // @[vga.scala 25:23]
          ram_927 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_928 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_928 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_929 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_929 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_930 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_930 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_931 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_931 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_932 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_932 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_933 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_933 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_934 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_934 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_935 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_935 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_936 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_936 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_937 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3a9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_937 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_938 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3aa == _GEN_8904) begin // @[vga.scala 25:23]
          ram_938 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_939 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ab == _GEN_8904) begin // @[vga.scala 25:23]
          ram_939 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_940 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ac == _GEN_8904) begin // @[vga.scala 25:23]
          ram_940 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_941 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ad == _GEN_8904) begin // @[vga.scala 25:23]
          ram_941 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_942 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ae == _GEN_8904) begin // @[vga.scala 25:23]
          ram_942 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_943 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3af == _GEN_8904) begin // @[vga.scala 25:23]
          ram_943 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_944 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_944 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_945 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_945 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_946 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_946 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_947 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_947 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_948 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_948 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_949 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_949 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_950 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_950 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_951 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_951 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_952 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_952 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_953 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3b9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_953 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_954 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ba == _GEN_8904) begin // @[vga.scala 25:23]
          ram_954 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_955 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3bb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_955 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_956 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3bc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_956 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_957 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3bd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_957 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_958 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3be == _GEN_8904) begin // @[vga.scala 25:23]
          ram_958 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_959 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3bf == _GEN_8904) begin // @[vga.scala 25:23]
          ram_959 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_960 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_960 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_961 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_961 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_962 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_962 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_963 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_963 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_964 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_964 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_965 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_965 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_966 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_966 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_967 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_967 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_968 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_968 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_969 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3c9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_969 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_970 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ca == _GEN_8904) begin // @[vga.scala 25:23]
          ram_970 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_971 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3cb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_971 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_972 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3cc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_972 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_973 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3cd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_973 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_974 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ce == _GEN_8904) begin // @[vga.scala 25:23]
          ram_974 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_975 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3cf == _GEN_8904) begin // @[vga.scala 25:23]
          ram_975 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_976 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_976 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_977 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_977 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_978 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_978 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_979 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_979 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_980 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_980 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_981 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_981 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_982 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_982 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_983 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_983 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_984 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_984 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_985 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3d9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_985 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_986 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3da == _GEN_8904) begin // @[vga.scala 25:23]
          ram_986 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_987 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3db == _GEN_8904) begin // @[vga.scala 25:23]
          ram_987 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_988 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3dc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_988 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_989 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3dd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_989 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_990 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3de == _GEN_8904) begin // @[vga.scala 25:23]
          ram_990 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_991 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3df == _GEN_8904) begin // @[vga.scala 25:23]
          ram_991 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_992 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_992 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_993 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_993 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_994 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_994 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_995 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_995 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_996 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_996 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_997 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_997 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_998 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_998 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_999 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_999 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1000 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1000 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1001 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3e9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1001 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1002 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ea == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1002 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1003 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3eb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1003 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1004 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ec == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1004 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1005 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ed == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1005 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1006 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ee == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1006 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1007 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ef == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1007 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1008 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f0 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1008 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1009 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f1 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1009 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1010 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f2 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1010 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1011 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f3 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1011 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1012 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f4 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1012 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1013 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f5 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1013 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1014 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f6 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1014 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1015 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f7 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1015 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1016 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f8 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1016 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1017 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3f9 == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1017 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1018 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3fa == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1018 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1019 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3fb == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1019 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1020 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3fc == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1020 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1021 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3fd == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1021 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1022 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3fe == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1022 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1023 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (10'h3ff == _GEN_8904) begin // @[vga.scala 25:23]
          ram_1023 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1024 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h400 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1024 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1025 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h401 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1025 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1026 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h402 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1026 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1027 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h403 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1027 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1028 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h404 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1028 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1029 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h405 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1029 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1030 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h406 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1030 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1031 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h407 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1031 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1032 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h408 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1032 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1033 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h409 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1033 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1034 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1034 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1035 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1035 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1036 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1036 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1037 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1037 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1038 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1038 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1039 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h40f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1039 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1040 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h410 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1040 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1041 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h411 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1041 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1042 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h412 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1042 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1043 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h413 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1043 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1044 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h414 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1044 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1045 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h415 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1045 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1046 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h416 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1046 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1047 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h417 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1047 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1048 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h418 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1048 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1049 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h419 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1049 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1050 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1050 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1051 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1051 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1052 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1052 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1053 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1053 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1054 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1054 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1055 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h41f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1055 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1056 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h420 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1056 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1057 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h421 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1057 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1058 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h422 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1058 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1059 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h423 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1059 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1060 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h424 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1060 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1061 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h425 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1061 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1062 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h426 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1062 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1063 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h427 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1063 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1064 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h428 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1064 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1065 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h429 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1065 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1066 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1066 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1067 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1067 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1068 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1068 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1069 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1069 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1070 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1070 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1071 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h42f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1071 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1072 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h430 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1072 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1073 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h431 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1073 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1074 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h432 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1074 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1075 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h433 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1075 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1076 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h434 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1076 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1077 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h435 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1077 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1078 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h436 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1078 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1079 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h437 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1079 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1080 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h438 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1080 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1081 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h439 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1081 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1082 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1082 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1083 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1083 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1084 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1084 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1085 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1085 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1086 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1086 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1087 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h43f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1087 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1088 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h440 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1088 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1089 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h441 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1089 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1090 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h442 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1090 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1091 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h443 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1091 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1092 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h444 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1092 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1093 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h445 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1093 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1094 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h446 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1094 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1095 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h447 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1095 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1096 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h448 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1096 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1097 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h449 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1097 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1098 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1098 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1099 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1099 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1100 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1100 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1101 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1101 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1102 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1102 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1103 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h44f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1103 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1104 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h450 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1104 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1105 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h451 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1105 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1106 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h452 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1106 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1107 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h453 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1107 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1108 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h454 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1108 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1109 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h455 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1109 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1110 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h456 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1110 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1111 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h457 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1111 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1112 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h458 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1112 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1113 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h459 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1113 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1114 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1114 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1115 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1115 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1116 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1116 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1117 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1117 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1118 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1118 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1119 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h45f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1119 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1120 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h460 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1120 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1121 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h461 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1121 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1122 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h462 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1122 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1123 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h463 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1123 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1124 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h464 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1124 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1125 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h465 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1125 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1126 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h466 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1126 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1127 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h467 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1127 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1128 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h468 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1128 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1129 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h469 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1129 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1130 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1130 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1131 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1131 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1132 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1132 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1133 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1133 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1134 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1134 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1135 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h46f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1135 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1136 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h470 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1136 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1137 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h471 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1137 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1138 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h472 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1138 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1139 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h473 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1139 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1140 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h474 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1140 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1141 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h475 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1141 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1142 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h476 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1142 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1143 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h477 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1143 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1144 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h478 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1144 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1145 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h479 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1145 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1146 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1146 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1147 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1147 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1148 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1148 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1149 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1149 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1150 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1150 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1151 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h47f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1151 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1152 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h480 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1152 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1153 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h481 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1153 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1154 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h482 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1154 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1155 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h483 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1155 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1156 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h484 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1156 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1157 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h485 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1157 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1158 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h486 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1158 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1159 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h487 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1159 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1160 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h488 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1160 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1161 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h489 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1161 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1162 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1162 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1163 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1163 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1164 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1164 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1165 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1165 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1166 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1166 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1167 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h48f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1167 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1168 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h490 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1168 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1169 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h491 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1169 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1170 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h492 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1170 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1171 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h493 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1171 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1172 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h494 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1172 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1173 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h495 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1173 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1174 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h496 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1174 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1175 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h497 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1175 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1176 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h498 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1176 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1177 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h499 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1177 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1178 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1178 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1179 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1179 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1180 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1180 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1181 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1181 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1182 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1182 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1183 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h49f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1183 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1184 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1184 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1185 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1185 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1186 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1186 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1187 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1187 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1188 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1188 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1189 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1189 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1190 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1190 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1191 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1191 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1192 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1192 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1193 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4a9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1193 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1194 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4aa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1194 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1195 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ab == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1195 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1196 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ac == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1196 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1197 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ad == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1197 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1198 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ae == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1198 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1199 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4af == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1199 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1200 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1200 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1201 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1201 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1202 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1202 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1203 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1203 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1204 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1204 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1205 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1205 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1206 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1206 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1207 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1207 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1208 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1208 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1209 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4b9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1209 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1210 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ba == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1210 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1211 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4bb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1211 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1212 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4bc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1212 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1213 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4bd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1213 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1214 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4be == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1214 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1215 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4bf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1215 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1216 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1216 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1217 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1217 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1218 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1218 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1219 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1219 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1220 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1220 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1221 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1221 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1222 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1222 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1223 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1223 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1224 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1224 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1225 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4c9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1225 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1226 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ca == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1226 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1227 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4cb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1227 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1228 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4cc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1228 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1229 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4cd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1229 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1230 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ce == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1230 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1231 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4cf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1231 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1232 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1232 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1233 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1233 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1234 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1234 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1235 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1235 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1236 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1236 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1237 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1237 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1238 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1238 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1239 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1239 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1240 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1240 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1241 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4d9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1241 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1242 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4da == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1242 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1243 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4db == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1243 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1244 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4dc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1244 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1245 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4dd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1245 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1246 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4de == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1246 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1247 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4df == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1247 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1248 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1248 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1249 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1249 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1250 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1250 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1251 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1251 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1252 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1252 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1253 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1253 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1254 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1254 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1255 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1255 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1256 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1256 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1257 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4e9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1257 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1258 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ea == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1258 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1259 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4eb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1259 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1260 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ec == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1260 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1261 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ed == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1261 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1262 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ee == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1262 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1263 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ef == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1263 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1264 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1264 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1265 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1265 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1266 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1266 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1267 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1267 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1268 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1268 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1269 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1269 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1270 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1270 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1271 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1271 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1272 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1272 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1273 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4f9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1273 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1274 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4fa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1274 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1275 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4fb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1275 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1276 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4fc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1276 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1277 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4fd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1277 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1278 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4fe == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1278 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1279 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h4ff == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1279 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1280 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h500 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1280 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1281 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h501 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1281 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1282 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h502 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1282 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1283 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h503 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1283 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1284 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h504 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1284 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1285 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h505 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1285 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1286 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h506 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1286 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1287 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h507 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1287 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1288 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h508 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1288 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1289 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h509 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1289 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1290 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1290 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1291 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1291 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1292 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1292 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1293 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1293 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1294 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1294 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1295 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h50f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1295 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1296 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h510 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1296 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1297 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h511 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1297 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1298 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h512 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1298 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1299 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h513 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1299 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1300 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h514 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1300 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1301 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h515 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1301 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1302 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h516 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1302 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1303 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h517 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1303 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1304 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h518 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1304 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1305 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h519 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1305 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1306 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1306 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1307 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1307 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1308 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1308 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1309 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1309 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1310 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1310 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1311 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h51f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1311 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1312 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h520 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1312 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1313 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h521 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1313 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1314 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h522 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1314 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1315 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h523 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1315 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1316 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h524 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1316 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1317 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h525 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1317 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1318 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h526 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1318 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1319 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h527 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1319 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1320 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h528 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1320 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1321 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h529 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1321 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1322 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1322 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1323 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1323 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1324 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1324 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1325 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1325 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1326 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1326 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1327 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h52f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1327 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1328 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h530 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1328 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1329 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h531 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1329 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1330 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h532 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1330 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1331 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h533 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1331 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1332 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h534 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1332 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1333 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h535 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1333 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1334 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h536 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1334 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1335 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h537 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1335 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1336 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h538 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1336 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1337 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h539 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1337 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1338 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1338 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1339 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1339 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1340 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1340 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1341 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1341 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1342 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1342 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1343 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h53f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1343 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1344 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h540 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1344 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1345 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h541 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1345 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1346 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h542 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1346 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1347 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h543 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1347 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1348 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h544 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1348 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1349 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h545 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1349 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1350 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h546 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1350 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1351 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h547 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1351 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1352 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h548 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1352 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1353 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h549 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1353 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1354 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1354 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1355 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1355 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1356 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1356 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1357 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1357 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1358 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1358 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1359 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h54f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1359 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1360 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h550 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1360 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1361 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h551 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1361 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1362 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h552 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1362 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1363 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h553 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1363 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1364 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h554 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1364 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1365 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h555 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1365 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1366 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h556 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1366 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1367 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h557 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1367 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1368 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h558 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1368 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1369 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h559 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1369 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1370 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1370 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1371 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1371 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1372 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1372 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1373 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1373 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1374 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1374 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1375 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h55f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1375 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1376 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h560 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1376 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1377 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h561 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1377 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1378 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h562 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1378 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1379 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h563 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1379 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1380 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h564 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1380 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1381 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h565 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1381 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1382 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h566 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1382 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1383 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h567 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1383 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1384 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h568 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1384 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1385 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h569 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1385 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1386 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1386 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1387 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1387 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1388 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1388 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1389 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1389 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1390 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1390 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1391 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h56f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1391 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1392 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h570 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1392 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1393 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h571 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1393 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1394 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h572 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1394 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1395 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h573 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1395 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1396 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h574 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1396 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1397 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h575 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1397 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1398 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h576 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1398 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1399 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h577 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1399 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1400 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h578 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1400 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1401 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h579 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1401 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1402 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1402 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1403 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1403 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1404 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1404 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1405 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1405 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1406 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1406 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1407 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h57f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1407 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1408 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h580 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1408 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1409 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h581 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1409 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1410 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h582 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1410 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1411 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h583 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1411 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1412 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h584 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1412 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1413 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h585 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1413 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1414 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h586 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1414 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1415 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h587 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1415 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1416 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h588 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1416 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1417 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h589 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1417 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1418 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1418 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1419 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1419 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1420 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1420 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1421 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1421 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1422 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1422 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1423 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h58f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1423 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1424 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h590 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1424 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1425 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h591 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1425 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1426 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h592 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1426 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1427 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h593 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1427 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1428 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h594 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1428 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1429 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h595 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1429 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1430 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h596 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1430 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1431 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h597 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1431 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1432 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h598 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1432 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1433 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h599 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1433 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1434 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1434 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1435 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1435 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1436 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1436 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1437 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1437 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1438 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1438 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1439 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h59f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1439 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1440 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1440 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1441 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1441 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1442 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1442 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1443 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1443 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1444 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1444 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1445 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1445 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1446 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1446 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1447 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1447 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1448 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1448 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1449 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5a9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1449 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1450 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5aa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1450 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1451 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ab == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1451 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1452 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ac == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1452 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1453 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ad == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1453 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1454 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ae == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1454 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1455 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5af == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1455 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1456 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1456 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1457 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1457 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1458 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1458 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1459 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1459 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1460 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1460 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1461 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1461 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1462 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1462 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1463 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1463 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1464 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1464 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1465 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5b9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1465 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1466 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ba == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1466 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1467 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5bb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1467 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1468 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5bc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1468 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1469 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5bd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1469 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1470 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5be == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1470 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1471 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5bf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1471 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1472 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1472 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1473 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1473 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1474 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1474 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1475 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1475 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1476 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1476 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1477 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1477 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1478 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1478 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1479 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1479 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1480 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1480 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1481 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5c9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1481 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1482 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ca == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1482 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1483 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5cb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1483 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1484 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5cc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1484 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1485 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5cd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1485 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1486 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ce == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1486 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1487 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5cf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1487 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1488 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1488 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1489 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1489 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1490 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1490 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1491 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1491 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1492 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1492 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1493 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1493 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1494 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1494 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1495 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1495 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1496 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1496 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1497 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5d9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1497 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1498 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5da == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1498 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1499 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5db == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1499 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1500 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5dc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1500 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1501 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5dd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1501 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1502 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5de == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1502 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1503 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5df == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1503 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1504 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1504 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1505 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1505 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1506 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1506 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1507 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1507 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1508 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1508 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1509 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1509 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1510 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1510 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1511 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1511 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1512 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1512 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1513 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5e9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1513 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1514 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ea == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1514 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1515 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5eb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1515 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1516 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ec == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1516 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1517 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ed == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1517 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1518 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ee == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1518 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1519 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ef == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1519 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1520 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1520 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1521 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1521 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1522 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1522 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1523 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1523 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1524 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1524 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1525 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1525 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1526 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1526 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1527 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1527 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1528 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1528 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1529 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5f9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1529 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1530 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5fa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1530 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1531 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5fb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1531 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1532 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5fc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1532 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1533 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5fd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1533 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1534 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5fe == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1534 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1535 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h5ff == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1535 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1536 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h600 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1536 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1537 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h601 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1537 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1538 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h602 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1538 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1539 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h603 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1539 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1540 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h604 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1540 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1541 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h605 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1541 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1542 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h606 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1542 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1543 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h607 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1543 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1544 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h608 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1544 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1545 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h609 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1545 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1546 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1546 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1547 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1547 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1548 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1548 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1549 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1549 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1550 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1550 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1551 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h60f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1551 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1552 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h610 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1552 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1553 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h611 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1553 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1554 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h612 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1554 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1555 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h613 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1555 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1556 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h614 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1556 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1557 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h615 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1557 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1558 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h616 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1558 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1559 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h617 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1559 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1560 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h618 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1560 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1561 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h619 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1561 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1562 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1562 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1563 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1563 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1564 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1564 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1565 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1565 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1566 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1566 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1567 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h61f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1567 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1568 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h620 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1568 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1569 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h621 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1569 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1570 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h622 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1570 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1571 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h623 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1571 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1572 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h624 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1572 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1573 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h625 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1573 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1574 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h626 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1574 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1575 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h627 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1575 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1576 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h628 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1576 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1577 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h629 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1577 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1578 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1578 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1579 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1579 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1580 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1580 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1581 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1581 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1582 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1582 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1583 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h62f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1583 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1584 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h630 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1584 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1585 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h631 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1585 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1586 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h632 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1586 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1587 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h633 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1587 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1588 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h634 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1588 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1589 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h635 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1589 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1590 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h636 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1590 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1591 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h637 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1591 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1592 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h638 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1592 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1593 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h639 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1593 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1594 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1594 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1595 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1595 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1596 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1596 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1597 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1597 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1598 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1598 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1599 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h63f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1599 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1600 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h640 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1600 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1601 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h641 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1601 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1602 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h642 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1602 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1603 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h643 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1603 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1604 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h644 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1604 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1605 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h645 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1605 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1606 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h646 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1606 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1607 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h647 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1607 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1608 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h648 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1608 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1609 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h649 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1609 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1610 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1610 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1611 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1611 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1612 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1612 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1613 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1613 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1614 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1614 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1615 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h64f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1615 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1616 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h650 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1616 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1617 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h651 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1617 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1618 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h652 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1618 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1619 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h653 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1619 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1620 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h654 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1620 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1621 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h655 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1621 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1622 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h656 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1622 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1623 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h657 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1623 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1624 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h658 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1624 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1625 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h659 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1625 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1626 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1626 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1627 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1627 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1628 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1628 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1629 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1629 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1630 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1630 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1631 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h65f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1631 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1632 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h660 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1632 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1633 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h661 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1633 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1634 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h662 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1634 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1635 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h663 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1635 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1636 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h664 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1636 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1637 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h665 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1637 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1638 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h666 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1638 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1639 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h667 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1639 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1640 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h668 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1640 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1641 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h669 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1641 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1642 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1642 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1643 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1643 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1644 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1644 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1645 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1645 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1646 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1646 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1647 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h66f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1647 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1648 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h670 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1648 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1649 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h671 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1649 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1650 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h672 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1650 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1651 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h673 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1651 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1652 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h674 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1652 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1653 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h675 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1653 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1654 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h676 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1654 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1655 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h677 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1655 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1656 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h678 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1656 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1657 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h679 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1657 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1658 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1658 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1659 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1659 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1660 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1660 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1661 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1661 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1662 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1662 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1663 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h67f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1663 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1664 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h680 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1664 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1665 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h681 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1665 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1666 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h682 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1666 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1667 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h683 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1667 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1668 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h684 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1668 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1669 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h685 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1669 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1670 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h686 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1670 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1671 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h687 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1671 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1672 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h688 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1672 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1673 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h689 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1673 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1674 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1674 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1675 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1675 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1676 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1676 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1677 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1677 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1678 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1678 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1679 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h68f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1679 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1680 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h690 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1680 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1681 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h691 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1681 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1682 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h692 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1682 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1683 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h693 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1683 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1684 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h694 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1684 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1685 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h695 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1685 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1686 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h696 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1686 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1687 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h697 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1687 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1688 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h698 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1688 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1689 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h699 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1689 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1690 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1690 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1691 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1691 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1692 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1692 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1693 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1693 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1694 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1694 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1695 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h69f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1695 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1696 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1696 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1697 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1697 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1698 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1698 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1699 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1699 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1700 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1700 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1701 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1701 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1702 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1702 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1703 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1703 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1704 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1704 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1705 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6a9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1705 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1706 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6aa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1706 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1707 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ab == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1707 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1708 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ac == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1708 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1709 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ad == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1709 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1710 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ae == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1710 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1711 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6af == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1711 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1712 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1712 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1713 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1713 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1714 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1714 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1715 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1715 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1716 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1716 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1717 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1717 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1718 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1718 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1719 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1719 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1720 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1720 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1721 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6b9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1721 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1722 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ba == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1722 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1723 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6bb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1723 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1724 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6bc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1724 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1725 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6bd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1725 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1726 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6be == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1726 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1727 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6bf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1727 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1728 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1728 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1729 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1729 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1730 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1730 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1731 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1731 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1732 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1732 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1733 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1733 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1734 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1734 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1735 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1735 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1736 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1736 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1737 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6c9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1737 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1738 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ca == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1738 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1739 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6cb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1739 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1740 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6cc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1740 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1741 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6cd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1741 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1742 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ce == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1742 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1743 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6cf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1743 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1744 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1744 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1745 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1745 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1746 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1746 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1747 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1747 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1748 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1748 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1749 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1749 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1750 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1750 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1751 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1751 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1752 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1752 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1753 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6d9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1753 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1754 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6da == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1754 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1755 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6db == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1755 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1756 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6dc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1756 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1757 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6dd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1757 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1758 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6de == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1758 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1759 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6df == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1759 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1760 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1760 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1761 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1761 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1762 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1762 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1763 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1763 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1764 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1764 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1765 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1765 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1766 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1766 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1767 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1767 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1768 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1768 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1769 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6e9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1769 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1770 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ea == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1770 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1771 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6eb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1771 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1772 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ec == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1772 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1773 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ed == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1773 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1774 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ee == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1774 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1775 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ef == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1775 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1776 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1776 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1777 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1777 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1778 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1778 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1779 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1779 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1780 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1780 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1781 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1781 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1782 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1782 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1783 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1783 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1784 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1784 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1785 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6f9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1785 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1786 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6fa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1786 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1787 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6fb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1787 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1788 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6fc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1788 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1789 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6fd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1789 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1790 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6fe == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1790 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1791 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h6ff == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1791 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1792 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h700 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1792 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1793 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h701 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1793 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1794 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h702 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1794 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1795 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h703 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1795 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1796 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h704 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1796 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1797 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h705 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1797 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1798 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h706 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1798 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1799 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h707 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1799 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1800 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h708 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1800 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1801 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h709 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1801 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1802 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1802 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1803 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1803 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1804 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1804 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1805 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1805 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1806 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1806 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1807 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h70f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1807 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1808 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h710 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1808 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1809 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h711 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1809 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1810 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h712 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1810 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1811 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h713 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1811 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1812 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h714 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1812 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1813 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h715 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1813 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1814 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h716 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1814 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1815 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h717 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1815 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1816 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h718 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1816 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1817 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h719 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1817 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1818 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1818 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1819 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1819 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1820 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1820 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1821 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1821 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1822 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1822 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1823 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h71f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1823 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1824 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h720 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1824 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1825 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h721 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1825 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1826 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h722 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1826 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1827 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h723 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1827 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1828 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h724 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1828 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1829 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h725 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1829 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1830 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h726 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1830 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1831 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h727 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1831 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1832 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h728 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1832 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1833 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h729 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1833 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1834 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1834 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1835 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1835 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1836 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1836 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1837 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1837 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1838 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1838 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1839 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h72f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1839 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1840 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h730 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1840 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1841 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h731 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1841 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1842 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h732 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1842 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1843 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h733 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1843 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1844 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h734 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1844 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1845 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h735 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1845 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1846 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h736 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1846 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1847 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h737 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1847 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1848 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h738 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1848 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1849 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h739 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1849 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1850 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1850 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1851 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1851 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1852 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1852 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1853 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1853 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1854 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1854 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1855 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h73f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1855 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1856 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h740 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1856 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1857 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h741 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1857 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1858 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h742 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1858 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1859 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h743 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1859 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1860 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h744 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1860 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1861 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h745 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1861 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1862 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h746 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1862 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1863 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h747 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1863 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1864 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h748 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1864 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1865 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h749 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1865 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1866 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1866 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1867 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1867 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1868 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1868 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1869 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1869 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1870 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1870 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1871 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h74f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1871 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1872 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h750 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1872 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1873 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h751 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1873 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1874 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h752 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1874 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1875 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h753 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1875 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1876 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h754 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1876 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1877 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h755 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1877 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1878 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h756 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1878 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1879 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h757 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1879 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1880 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h758 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1880 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1881 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h759 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1881 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1882 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1882 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1883 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1883 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1884 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1884 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1885 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1885 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1886 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1886 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1887 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h75f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1887 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1888 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h760 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1888 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1889 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h761 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1889 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1890 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h762 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1890 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1891 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h763 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1891 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1892 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h764 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1892 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1893 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h765 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1893 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1894 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h766 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1894 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1895 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h767 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1895 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1896 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h768 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1896 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1897 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h769 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1897 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1898 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1898 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1899 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1899 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1900 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1900 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1901 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1901 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1902 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1902 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1903 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h76f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1903 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1904 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h770 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1904 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1905 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h771 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1905 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1906 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h772 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1906 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1907 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h773 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1907 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1908 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h774 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1908 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1909 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h775 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1909 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1910 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h776 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1910 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1911 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h777 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1911 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1912 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h778 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1912 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1913 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h779 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1913 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1914 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1914 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1915 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1915 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1916 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1916 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1917 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1917 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1918 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1918 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1919 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h77f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1919 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1920 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h780 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1920 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1921 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h781 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1921 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1922 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h782 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1922 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1923 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h783 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1923 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1924 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h784 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1924 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1925 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h785 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1925 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1926 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h786 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1926 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1927 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h787 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1927 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1928 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h788 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1928 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1929 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h789 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1929 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1930 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1930 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1931 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1931 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1932 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1932 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1933 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1933 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1934 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1934 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1935 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h78f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1935 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1936 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h790 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1936 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1937 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h791 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1937 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1938 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h792 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1938 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1939 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h793 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1939 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1940 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h794 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1940 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1941 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h795 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1941 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1942 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h796 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1942 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1943 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h797 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1943 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1944 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h798 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1944 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1945 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h799 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1945 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1946 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79a == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1946 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1947 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79b == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1947 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1948 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79c == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1948 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1949 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79d == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1949 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1950 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79e == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1950 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1951 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h79f == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1951 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1952 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1952 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1953 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1953 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1954 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1954 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1955 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1955 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1956 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1956 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1957 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1957 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1958 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1958 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1959 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1959 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1960 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1960 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1961 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7a9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1961 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1962 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7aa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1962 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1963 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ab == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1963 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1964 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ac == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1964 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1965 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ad == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1965 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1966 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ae == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1966 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1967 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7af == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1967 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1968 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1968 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1969 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1969 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1970 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1970 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1971 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1971 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1972 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1972 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1973 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1973 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1974 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1974 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1975 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1975 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1976 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1976 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1977 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7b9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1977 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1978 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ba == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1978 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1979 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7bb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1979 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1980 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7bc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1980 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1981 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7bd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1981 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1982 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7be == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1982 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1983 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7bf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1983 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1984 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1984 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1985 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1985 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1986 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1986 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1987 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1987 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1988 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1988 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1989 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1989 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1990 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1990 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1991 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1991 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1992 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1992 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1993 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7c9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1993 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1994 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ca == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1994 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1995 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7cb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1995 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1996 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7cc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1996 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1997 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7cd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1997 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1998 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ce == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1998 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_1999 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7cf == _GEN_9416) begin // @[vga.scala 25:23]
          ram_1999 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2000 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2000 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2001 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2001 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2002 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2002 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2003 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2003 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2004 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2004 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2005 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2005 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2006 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2006 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2007 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2007 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2008 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2008 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2009 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7d9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2009 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2010 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7da == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2010 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2011 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7db == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2011 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2012 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7dc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2012 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2013 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7dd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2013 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2014 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7de == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2014 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2015 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7df == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2015 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2016 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2016 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2017 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2017 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2018 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2018 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2019 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2019 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2020 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2020 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2021 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2021 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2022 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2022 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2023 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2023 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2024 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2024 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2025 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7e9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2025 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2026 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ea == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2026 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2027 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7eb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2027 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2028 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ec == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2028 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2029 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ed == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2029 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2030 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ee == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2030 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2031 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ef == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2031 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2032 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f0 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2032 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2033 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f1 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2033 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2034 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f2 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2034 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2035 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f3 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2035 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2036 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f4 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2036 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2037 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f5 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2037 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2038 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f6 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2038 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2039 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f7 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2039 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2040 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f8 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2040 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2041 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7f9 == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2041 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2042 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7fa == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2042 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2043 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7fb == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2043 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2044 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7fc == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2044 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2045 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7fd == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2045 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2046 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7fe == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2046 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2047 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (11'h7ff == _GEN_9416) begin // @[vga.scala 25:23]
          ram_2047 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2048 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h800 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2048 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2049 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h801 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2049 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2050 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h802 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2050 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2051 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h803 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2051 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2052 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h804 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2052 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2053 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h805 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2053 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2054 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h806 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2054 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2055 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h807 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2055 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2056 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h808 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2056 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2057 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h809 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2057 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2058 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2058 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2059 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2059 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2060 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2060 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2061 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2061 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2062 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2062 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2063 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h80f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2063 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2064 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h810 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2064 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2065 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h811 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2065 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2066 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h812 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2066 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2067 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h813 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2067 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2068 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h814 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2068 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2069 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h815 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2069 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2070 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h816 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2070 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2071 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h817 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2071 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2072 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h818 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2072 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2073 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h819 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2073 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2074 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2074 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2075 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2075 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2076 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2076 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2077 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2077 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2078 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2078 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2079 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h81f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2079 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2080 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h820 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2080 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2081 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h821 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2081 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2082 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h822 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2082 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2083 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h823 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2083 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2084 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h824 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2084 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2085 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h825 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2085 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2086 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h826 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2086 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2087 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h827 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2087 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2088 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h828 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2088 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2089 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h829 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2089 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2090 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2090 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2091 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2091 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2092 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2092 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2093 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2093 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2094 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2094 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2095 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h82f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2095 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2096 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h830 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2096 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2097 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h831 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2097 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2098 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h832 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2098 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2099 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h833 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2099 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2100 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h834 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2100 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2101 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h835 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2101 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2102 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h836 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2102 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2103 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h837 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2103 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2104 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h838 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2104 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2105 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h839 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2105 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2106 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2106 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2107 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2107 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2108 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2108 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2109 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2109 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2110 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2110 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2111 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h83f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2111 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2112 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h840 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2112 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2113 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h841 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2113 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2114 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h842 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2114 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2115 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h843 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2115 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2116 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h844 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2116 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2117 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h845 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2117 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2118 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h846 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2118 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2119 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h847 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2119 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2120 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h848 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2120 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2121 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h849 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2121 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2122 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2122 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2123 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2123 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2124 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2124 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2125 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2125 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2126 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2126 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2127 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h84f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2127 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2128 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h850 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2128 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2129 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h851 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2129 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2130 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h852 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2130 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2131 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h853 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2131 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2132 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h854 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2132 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2133 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h855 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2133 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2134 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h856 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2134 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2135 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h857 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2135 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2136 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h858 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2136 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2137 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h859 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2137 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2138 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2138 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2139 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2139 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2140 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2140 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2141 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2141 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2142 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2142 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2143 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h85f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2143 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2144 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h860 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2144 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2145 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h861 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2145 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2146 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h862 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2146 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2147 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h863 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2147 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2148 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h864 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2148 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2149 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h865 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2149 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2150 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h866 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2150 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2151 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h867 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2151 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2152 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h868 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2152 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2153 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h869 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2153 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2154 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86a == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2154 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2155 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86b == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2155 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2156 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86c == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2156 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2157 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86d == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2157 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2158 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86e == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2158 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2159 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h86f == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2159 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 14:20]
      ram_2160 <= 8'h0; // @[vga.scala 14:20]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (!(io_ascii == 8'ha)) begin // @[vga.scala 22:30]
        if (12'h870 == _GEN_10440) begin // @[vga.scala 25:23]
          ram_2160 <= io_ascii; // @[vga.scala 25:23]
        end
      end
    end
    if (reset) begin // @[vga.scala 20:22]
      index <= 8'h0; // @[vga.scala 20:22]
    end else if (io_w_en) begin // @[vga.scala 21:24]
      if (io_ascii == 8'ha) begin // @[vga.scala 22:30]
        index <= _index_T_6; // @[vga.scala 23:18]
      end else begin
        index <= _index_T_8; // @[vga.scala 26:18]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
  integer initvar;
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vga_mem_MPORT_addr_pipe_0 = _RAND_0[11:0];
  _RAND_1 = {1{`RANDOM}};
  rdwrPort = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  ram_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  ram_1 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  ram_2 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  ram_3 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  ram_4 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  ram_5 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  ram_6 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  ram_7 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  ram_8 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  ram_9 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  ram_10 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  ram_11 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  ram_12 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  ram_13 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  ram_14 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  ram_15 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  ram_16 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  ram_17 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  ram_18 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  ram_19 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  ram_20 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  ram_21 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  ram_22 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  ram_23 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  ram_24 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  ram_25 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  ram_26 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  ram_27 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  ram_28 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  ram_29 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  ram_30 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  ram_31 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  ram_32 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  ram_33 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  ram_34 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  ram_35 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  ram_36 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  ram_37 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  ram_38 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  ram_39 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  ram_40 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  ram_41 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  ram_42 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  ram_43 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  ram_44 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  ram_45 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  ram_46 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  ram_47 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  ram_48 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  ram_49 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  ram_50 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  ram_51 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  ram_52 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  ram_53 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  ram_54 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  ram_55 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  ram_56 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  ram_57 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  ram_58 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  ram_59 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  ram_60 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  ram_61 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  ram_62 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  ram_63 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  ram_64 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  ram_65 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  ram_66 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  ram_67 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  ram_68 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  ram_69 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  ram_70 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  ram_71 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  ram_72 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  ram_73 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  ram_74 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  ram_75 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  ram_76 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  ram_77 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  ram_78 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  ram_79 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  ram_80 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  ram_81 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  ram_82 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  ram_83 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  ram_84 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  ram_85 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  ram_86 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  ram_87 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  ram_88 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  ram_89 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  ram_90 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  ram_91 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  ram_92 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  ram_93 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  ram_94 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  ram_95 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  ram_96 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  ram_97 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  ram_98 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  ram_99 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  ram_100 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  ram_101 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  ram_102 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  ram_103 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  ram_104 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  ram_105 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  ram_106 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  ram_107 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  ram_108 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  ram_109 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  ram_110 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  ram_111 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  ram_112 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  ram_113 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  ram_114 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  ram_115 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  ram_116 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  ram_117 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  ram_118 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  ram_119 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  ram_120 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  ram_121 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  ram_122 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  ram_123 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  ram_124 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  ram_125 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  ram_126 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  ram_127 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  ram_128 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  ram_129 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  ram_130 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  ram_131 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  ram_132 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  ram_133 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  ram_134 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  ram_135 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  ram_136 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  ram_137 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  ram_138 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  ram_139 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  ram_140 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  ram_141 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  ram_142 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  ram_143 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  ram_144 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  ram_145 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  ram_146 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  ram_147 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  ram_148 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  ram_149 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  ram_150 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  ram_151 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  ram_152 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  ram_153 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  ram_154 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  ram_155 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  ram_156 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  ram_157 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  ram_158 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  ram_159 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  ram_160 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  ram_161 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  ram_162 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  ram_163 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  ram_164 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  ram_165 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  ram_166 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  ram_167 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  ram_168 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  ram_169 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  ram_170 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  ram_171 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  ram_172 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  ram_173 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  ram_174 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  ram_175 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  ram_176 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  ram_177 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  ram_178 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  ram_179 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ram_180 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ram_181 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  ram_182 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  ram_183 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  ram_184 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  ram_185 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  ram_186 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  ram_187 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  ram_188 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  ram_189 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  ram_190 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  ram_191 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  ram_192 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  ram_193 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  ram_194 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  ram_195 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  ram_196 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  ram_197 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  ram_198 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  ram_199 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  ram_200 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  ram_201 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  ram_202 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  ram_203 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  ram_204 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  ram_205 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  ram_206 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  ram_207 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  ram_208 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  ram_209 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  ram_210 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  ram_211 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  ram_212 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  ram_213 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  ram_214 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  ram_215 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  ram_216 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  ram_217 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  ram_218 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  ram_219 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  ram_220 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  ram_221 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  ram_222 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  ram_223 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  ram_224 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  ram_225 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  ram_226 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  ram_227 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  ram_228 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  ram_229 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  ram_230 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  ram_231 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  ram_232 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  ram_233 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  ram_234 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  ram_235 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  ram_236 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  ram_237 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  ram_238 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  ram_239 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  ram_240 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  ram_241 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  ram_242 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  ram_243 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  ram_244 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  ram_245 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  ram_246 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  ram_247 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  ram_248 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  ram_249 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  ram_250 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  ram_251 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  ram_252 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  ram_253 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  ram_254 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  ram_255 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  ram_256 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  ram_257 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  ram_258 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  ram_259 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  ram_260 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  ram_261 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  ram_262 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  ram_263 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  ram_264 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  ram_265 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  ram_266 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  ram_267 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  ram_268 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  ram_269 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  ram_270 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  ram_271 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  ram_272 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  ram_273 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  ram_274 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  ram_275 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  ram_276 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  ram_277 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  ram_278 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  ram_279 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  ram_280 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  ram_281 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  ram_282 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  ram_283 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  ram_284 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  ram_285 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  ram_286 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  ram_287 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  ram_288 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  ram_289 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  ram_290 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  ram_291 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  ram_292 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  ram_293 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  ram_294 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  ram_295 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  ram_296 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  ram_297 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  ram_298 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  ram_299 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  ram_300 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  ram_301 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  ram_302 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  ram_303 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  ram_304 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  ram_305 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  ram_306 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  ram_307 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  ram_308 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  ram_309 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  ram_310 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  ram_311 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  ram_312 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  ram_313 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  ram_314 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  ram_315 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  ram_316 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  ram_317 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  ram_318 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  ram_319 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  ram_320 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  ram_321 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  ram_322 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  ram_323 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  ram_324 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  ram_325 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  ram_326 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  ram_327 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  ram_328 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  ram_329 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  ram_330 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  ram_331 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  ram_332 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  ram_333 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  ram_334 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  ram_335 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  ram_336 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  ram_337 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  ram_338 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  ram_339 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  ram_340 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  ram_341 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  ram_342 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  ram_343 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  ram_344 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  ram_345 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  ram_346 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  ram_347 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  ram_348 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  ram_349 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  ram_350 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  ram_351 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  ram_352 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  ram_353 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  ram_354 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  ram_355 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  ram_356 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  ram_357 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  ram_358 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  ram_359 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  ram_360 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  ram_361 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  ram_362 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  ram_363 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  ram_364 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  ram_365 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  ram_366 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  ram_367 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  ram_368 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  ram_369 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  ram_370 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  ram_371 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  ram_372 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  ram_373 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  ram_374 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  ram_375 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  ram_376 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  ram_377 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  ram_378 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  ram_379 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  ram_380 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  ram_381 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  ram_382 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  ram_383 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  ram_384 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  ram_385 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  ram_386 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  ram_387 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  ram_388 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  ram_389 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  ram_390 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  ram_391 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  ram_392 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  ram_393 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  ram_394 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  ram_395 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  ram_396 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  ram_397 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  ram_398 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  ram_399 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  ram_400 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  ram_401 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  ram_402 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  ram_403 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  ram_404 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  ram_405 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  ram_406 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  ram_407 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  ram_408 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  ram_409 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  ram_410 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  ram_411 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  ram_412 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  ram_413 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  ram_414 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  ram_415 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  ram_416 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  ram_417 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  ram_418 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  ram_419 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  ram_420 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  ram_421 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  ram_422 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  ram_423 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  ram_424 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  ram_425 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  ram_426 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  ram_427 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  ram_428 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  ram_429 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  ram_430 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  ram_431 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  ram_432 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  ram_433 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  ram_434 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  ram_435 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  ram_436 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  ram_437 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  ram_438 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  ram_439 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  ram_440 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  ram_441 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  ram_442 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  ram_443 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  ram_444 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  ram_445 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  ram_446 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  ram_447 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  ram_448 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  ram_449 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  ram_450 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  ram_451 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  ram_452 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  ram_453 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  ram_454 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  ram_455 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  ram_456 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  ram_457 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  ram_458 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  ram_459 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  ram_460 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  ram_461 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  ram_462 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  ram_463 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  ram_464 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  ram_465 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  ram_466 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  ram_467 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  ram_468 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  ram_469 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  ram_470 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  ram_471 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  ram_472 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  ram_473 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  ram_474 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  ram_475 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  ram_476 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  ram_477 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  ram_478 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  ram_479 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  ram_480 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  ram_481 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  ram_482 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  ram_483 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  ram_484 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  ram_485 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  ram_486 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  ram_487 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  ram_488 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  ram_489 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  ram_490 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  ram_491 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  ram_492 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  ram_493 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  ram_494 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  ram_495 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  ram_496 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  ram_497 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  ram_498 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  ram_499 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  ram_500 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  ram_501 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  ram_502 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  ram_503 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  ram_504 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  ram_505 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  ram_506 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  ram_507 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  ram_508 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  ram_509 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  ram_510 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  ram_511 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  ram_512 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  ram_513 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  ram_514 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  ram_515 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  ram_516 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  ram_517 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  ram_518 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  ram_519 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  ram_520 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  ram_521 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  ram_522 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  ram_523 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  ram_524 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  ram_525 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  ram_526 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  ram_527 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  ram_528 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  ram_529 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  ram_530 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  ram_531 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  ram_532 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  ram_533 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  ram_534 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  ram_535 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  ram_536 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  ram_537 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  ram_538 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  ram_539 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  ram_540 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  ram_541 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  ram_542 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  ram_543 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  ram_544 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  ram_545 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  ram_546 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  ram_547 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  ram_548 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  ram_549 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  ram_550 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  ram_551 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  ram_552 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  ram_553 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  ram_554 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  ram_555 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  ram_556 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  ram_557 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  ram_558 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  ram_559 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  ram_560 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  ram_561 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  ram_562 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  ram_563 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  ram_564 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  ram_565 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  ram_566 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  ram_567 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  ram_568 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  ram_569 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  ram_570 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  ram_571 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  ram_572 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  ram_573 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  ram_574 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  ram_575 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  ram_576 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  ram_577 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  ram_578 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  ram_579 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  ram_580 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  ram_581 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  ram_582 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  ram_583 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  ram_584 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  ram_585 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  ram_586 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  ram_587 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  ram_588 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  ram_589 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  ram_590 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  ram_591 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  ram_592 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  ram_593 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  ram_594 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  ram_595 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  ram_596 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  ram_597 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  ram_598 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  ram_599 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  ram_600 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  ram_601 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  ram_602 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  ram_603 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  ram_604 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  ram_605 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  ram_606 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  ram_607 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  ram_608 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  ram_609 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  ram_610 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  ram_611 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  ram_612 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  ram_613 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  ram_614 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  ram_615 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  ram_616 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  ram_617 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  ram_618 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  ram_619 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  ram_620 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  ram_621 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  ram_622 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  ram_623 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  ram_624 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  ram_625 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  ram_626 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  ram_627 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  ram_628 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  ram_629 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  ram_630 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  ram_631 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  ram_632 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  ram_633 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  ram_634 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  ram_635 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  ram_636 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  ram_637 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  ram_638 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  ram_639 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  ram_640 = _RAND_642[7:0];
  _RAND_643 = {1{`RANDOM}};
  ram_641 = _RAND_643[7:0];
  _RAND_644 = {1{`RANDOM}};
  ram_642 = _RAND_644[7:0];
  _RAND_645 = {1{`RANDOM}};
  ram_643 = _RAND_645[7:0];
  _RAND_646 = {1{`RANDOM}};
  ram_644 = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  ram_645 = _RAND_647[7:0];
  _RAND_648 = {1{`RANDOM}};
  ram_646 = _RAND_648[7:0];
  _RAND_649 = {1{`RANDOM}};
  ram_647 = _RAND_649[7:0];
  _RAND_650 = {1{`RANDOM}};
  ram_648 = _RAND_650[7:0];
  _RAND_651 = {1{`RANDOM}};
  ram_649 = _RAND_651[7:0];
  _RAND_652 = {1{`RANDOM}};
  ram_650 = _RAND_652[7:0];
  _RAND_653 = {1{`RANDOM}};
  ram_651 = _RAND_653[7:0];
  _RAND_654 = {1{`RANDOM}};
  ram_652 = _RAND_654[7:0];
  _RAND_655 = {1{`RANDOM}};
  ram_653 = _RAND_655[7:0];
  _RAND_656 = {1{`RANDOM}};
  ram_654 = _RAND_656[7:0];
  _RAND_657 = {1{`RANDOM}};
  ram_655 = _RAND_657[7:0];
  _RAND_658 = {1{`RANDOM}};
  ram_656 = _RAND_658[7:0];
  _RAND_659 = {1{`RANDOM}};
  ram_657 = _RAND_659[7:0];
  _RAND_660 = {1{`RANDOM}};
  ram_658 = _RAND_660[7:0];
  _RAND_661 = {1{`RANDOM}};
  ram_659 = _RAND_661[7:0];
  _RAND_662 = {1{`RANDOM}};
  ram_660 = _RAND_662[7:0];
  _RAND_663 = {1{`RANDOM}};
  ram_661 = _RAND_663[7:0];
  _RAND_664 = {1{`RANDOM}};
  ram_662 = _RAND_664[7:0];
  _RAND_665 = {1{`RANDOM}};
  ram_663 = _RAND_665[7:0];
  _RAND_666 = {1{`RANDOM}};
  ram_664 = _RAND_666[7:0];
  _RAND_667 = {1{`RANDOM}};
  ram_665 = _RAND_667[7:0];
  _RAND_668 = {1{`RANDOM}};
  ram_666 = _RAND_668[7:0];
  _RAND_669 = {1{`RANDOM}};
  ram_667 = _RAND_669[7:0];
  _RAND_670 = {1{`RANDOM}};
  ram_668 = _RAND_670[7:0];
  _RAND_671 = {1{`RANDOM}};
  ram_669 = _RAND_671[7:0];
  _RAND_672 = {1{`RANDOM}};
  ram_670 = _RAND_672[7:0];
  _RAND_673 = {1{`RANDOM}};
  ram_671 = _RAND_673[7:0];
  _RAND_674 = {1{`RANDOM}};
  ram_672 = _RAND_674[7:0];
  _RAND_675 = {1{`RANDOM}};
  ram_673 = _RAND_675[7:0];
  _RAND_676 = {1{`RANDOM}};
  ram_674 = _RAND_676[7:0];
  _RAND_677 = {1{`RANDOM}};
  ram_675 = _RAND_677[7:0];
  _RAND_678 = {1{`RANDOM}};
  ram_676 = _RAND_678[7:0];
  _RAND_679 = {1{`RANDOM}};
  ram_677 = _RAND_679[7:0];
  _RAND_680 = {1{`RANDOM}};
  ram_678 = _RAND_680[7:0];
  _RAND_681 = {1{`RANDOM}};
  ram_679 = _RAND_681[7:0];
  _RAND_682 = {1{`RANDOM}};
  ram_680 = _RAND_682[7:0];
  _RAND_683 = {1{`RANDOM}};
  ram_681 = _RAND_683[7:0];
  _RAND_684 = {1{`RANDOM}};
  ram_682 = _RAND_684[7:0];
  _RAND_685 = {1{`RANDOM}};
  ram_683 = _RAND_685[7:0];
  _RAND_686 = {1{`RANDOM}};
  ram_684 = _RAND_686[7:0];
  _RAND_687 = {1{`RANDOM}};
  ram_685 = _RAND_687[7:0];
  _RAND_688 = {1{`RANDOM}};
  ram_686 = _RAND_688[7:0];
  _RAND_689 = {1{`RANDOM}};
  ram_687 = _RAND_689[7:0];
  _RAND_690 = {1{`RANDOM}};
  ram_688 = _RAND_690[7:0];
  _RAND_691 = {1{`RANDOM}};
  ram_689 = _RAND_691[7:0];
  _RAND_692 = {1{`RANDOM}};
  ram_690 = _RAND_692[7:0];
  _RAND_693 = {1{`RANDOM}};
  ram_691 = _RAND_693[7:0];
  _RAND_694 = {1{`RANDOM}};
  ram_692 = _RAND_694[7:0];
  _RAND_695 = {1{`RANDOM}};
  ram_693 = _RAND_695[7:0];
  _RAND_696 = {1{`RANDOM}};
  ram_694 = _RAND_696[7:0];
  _RAND_697 = {1{`RANDOM}};
  ram_695 = _RAND_697[7:0];
  _RAND_698 = {1{`RANDOM}};
  ram_696 = _RAND_698[7:0];
  _RAND_699 = {1{`RANDOM}};
  ram_697 = _RAND_699[7:0];
  _RAND_700 = {1{`RANDOM}};
  ram_698 = _RAND_700[7:0];
  _RAND_701 = {1{`RANDOM}};
  ram_699 = _RAND_701[7:0];
  _RAND_702 = {1{`RANDOM}};
  ram_700 = _RAND_702[7:0];
  _RAND_703 = {1{`RANDOM}};
  ram_701 = _RAND_703[7:0];
  _RAND_704 = {1{`RANDOM}};
  ram_702 = _RAND_704[7:0];
  _RAND_705 = {1{`RANDOM}};
  ram_703 = _RAND_705[7:0];
  _RAND_706 = {1{`RANDOM}};
  ram_704 = _RAND_706[7:0];
  _RAND_707 = {1{`RANDOM}};
  ram_705 = _RAND_707[7:0];
  _RAND_708 = {1{`RANDOM}};
  ram_706 = _RAND_708[7:0];
  _RAND_709 = {1{`RANDOM}};
  ram_707 = _RAND_709[7:0];
  _RAND_710 = {1{`RANDOM}};
  ram_708 = _RAND_710[7:0];
  _RAND_711 = {1{`RANDOM}};
  ram_709 = _RAND_711[7:0];
  _RAND_712 = {1{`RANDOM}};
  ram_710 = _RAND_712[7:0];
  _RAND_713 = {1{`RANDOM}};
  ram_711 = _RAND_713[7:0];
  _RAND_714 = {1{`RANDOM}};
  ram_712 = _RAND_714[7:0];
  _RAND_715 = {1{`RANDOM}};
  ram_713 = _RAND_715[7:0];
  _RAND_716 = {1{`RANDOM}};
  ram_714 = _RAND_716[7:0];
  _RAND_717 = {1{`RANDOM}};
  ram_715 = _RAND_717[7:0];
  _RAND_718 = {1{`RANDOM}};
  ram_716 = _RAND_718[7:0];
  _RAND_719 = {1{`RANDOM}};
  ram_717 = _RAND_719[7:0];
  _RAND_720 = {1{`RANDOM}};
  ram_718 = _RAND_720[7:0];
  _RAND_721 = {1{`RANDOM}};
  ram_719 = _RAND_721[7:0];
  _RAND_722 = {1{`RANDOM}};
  ram_720 = _RAND_722[7:0];
  _RAND_723 = {1{`RANDOM}};
  ram_721 = _RAND_723[7:0];
  _RAND_724 = {1{`RANDOM}};
  ram_722 = _RAND_724[7:0];
  _RAND_725 = {1{`RANDOM}};
  ram_723 = _RAND_725[7:0];
  _RAND_726 = {1{`RANDOM}};
  ram_724 = _RAND_726[7:0];
  _RAND_727 = {1{`RANDOM}};
  ram_725 = _RAND_727[7:0];
  _RAND_728 = {1{`RANDOM}};
  ram_726 = _RAND_728[7:0];
  _RAND_729 = {1{`RANDOM}};
  ram_727 = _RAND_729[7:0];
  _RAND_730 = {1{`RANDOM}};
  ram_728 = _RAND_730[7:0];
  _RAND_731 = {1{`RANDOM}};
  ram_729 = _RAND_731[7:0];
  _RAND_732 = {1{`RANDOM}};
  ram_730 = _RAND_732[7:0];
  _RAND_733 = {1{`RANDOM}};
  ram_731 = _RAND_733[7:0];
  _RAND_734 = {1{`RANDOM}};
  ram_732 = _RAND_734[7:0];
  _RAND_735 = {1{`RANDOM}};
  ram_733 = _RAND_735[7:0];
  _RAND_736 = {1{`RANDOM}};
  ram_734 = _RAND_736[7:0];
  _RAND_737 = {1{`RANDOM}};
  ram_735 = _RAND_737[7:0];
  _RAND_738 = {1{`RANDOM}};
  ram_736 = _RAND_738[7:0];
  _RAND_739 = {1{`RANDOM}};
  ram_737 = _RAND_739[7:0];
  _RAND_740 = {1{`RANDOM}};
  ram_738 = _RAND_740[7:0];
  _RAND_741 = {1{`RANDOM}};
  ram_739 = _RAND_741[7:0];
  _RAND_742 = {1{`RANDOM}};
  ram_740 = _RAND_742[7:0];
  _RAND_743 = {1{`RANDOM}};
  ram_741 = _RAND_743[7:0];
  _RAND_744 = {1{`RANDOM}};
  ram_742 = _RAND_744[7:0];
  _RAND_745 = {1{`RANDOM}};
  ram_743 = _RAND_745[7:0];
  _RAND_746 = {1{`RANDOM}};
  ram_744 = _RAND_746[7:0];
  _RAND_747 = {1{`RANDOM}};
  ram_745 = _RAND_747[7:0];
  _RAND_748 = {1{`RANDOM}};
  ram_746 = _RAND_748[7:0];
  _RAND_749 = {1{`RANDOM}};
  ram_747 = _RAND_749[7:0];
  _RAND_750 = {1{`RANDOM}};
  ram_748 = _RAND_750[7:0];
  _RAND_751 = {1{`RANDOM}};
  ram_749 = _RAND_751[7:0];
  _RAND_752 = {1{`RANDOM}};
  ram_750 = _RAND_752[7:0];
  _RAND_753 = {1{`RANDOM}};
  ram_751 = _RAND_753[7:0];
  _RAND_754 = {1{`RANDOM}};
  ram_752 = _RAND_754[7:0];
  _RAND_755 = {1{`RANDOM}};
  ram_753 = _RAND_755[7:0];
  _RAND_756 = {1{`RANDOM}};
  ram_754 = _RAND_756[7:0];
  _RAND_757 = {1{`RANDOM}};
  ram_755 = _RAND_757[7:0];
  _RAND_758 = {1{`RANDOM}};
  ram_756 = _RAND_758[7:0];
  _RAND_759 = {1{`RANDOM}};
  ram_757 = _RAND_759[7:0];
  _RAND_760 = {1{`RANDOM}};
  ram_758 = _RAND_760[7:0];
  _RAND_761 = {1{`RANDOM}};
  ram_759 = _RAND_761[7:0];
  _RAND_762 = {1{`RANDOM}};
  ram_760 = _RAND_762[7:0];
  _RAND_763 = {1{`RANDOM}};
  ram_761 = _RAND_763[7:0];
  _RAND_764 = {1{`RANDOM}};
  ram_762 = _RAND_764[7:0];
  _RAND_765 = {1{`RANDOM}};
  ram_763 = _RAND_765[7:0];
  _RAND_766 = {1{`RANDOM}};
  ram_764 = _RAND_766[7:0];
  _RAND_767 = {1{`RANDOM}};
  ram_765 = _RAND_767[7:0];
  _RAND_768 = {1{`RANDOM}};
  ram_766 = _RAND_768[7:0];
  _RAND_769 = {1{`RANDOM}};
  ram_767 = _RAND_769[7:0];
  _RAND_770 = {1{`RANDOM}};
  ram_768 = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  ram_769 = _RAND_771[7:0];
  _RAND_772 = {1{`RANDOM}};
  ram_770 = _RAND_772[7:0];
  _RAND_773 = {1{`RANDOM}};
  ram_771 = _RAND_773[7:0];
  _RAND_774 = {1{`RANDOM}};
  ram_772 = _RAND_774[7:0];
  _RAND_775 = {1{`RANDOM}};
  ram_773 = _RAND_775[7:0];
  _RAND_776 = {1{`RANDOM}};
  ram_774 = _RAND_776[7:0];
  _RAND_777 = {1{`RANDOM}};
  ram_775 = _RAND_777[7:0];
  _RAND_778 = {1{`RANDOM}};
  ram_776 = _RAND_778[7:0];
  _RAND_779 = {1{`RANDOM}};
  ram_777 = _RAND_779[7:0];
  _RAND_780 = {1{`RANDOM}};
  ram_778 = _RAND_780[7:0];
  _RAND_781 = {1{`RANDOM}};
  ram_779 = _RAND_781[7:0];
  _RAND_782 = {1{`RANDOM}};
  ram_780 = _RAND_782[7:0];
  _RAND_783 = {1{`RANDOM}};
  ram_781 = _RAND_783[7:0];
  _RAND_784 = {1{`RANDOM}};
  ram_782 = _RAND_784[7:0];
  _RAND_785 = {1{`RANDOM}};
  ram_783 = _RAND_785[7:0];
  _RAND_786 = {1{`RANDOM}};
  ram_784 = _RAND_786[7:0];
  _RAND_787 = {1{`RANDOM}};
  ram_785 = _RAND_787[7:0];
  _RAND_788 = {1{`RANDOM}};
  ram_786 = _RAND_788[7:0];
  _RAND_789 = {1{`RANDOM}};
  ram_787 = _RAND_789[7:0];
  _RAND_790 = {1{`RANDOM}};
  ram_788 = _RAND_790[7:0];
  _RAND_791 = {1{`RANDOM}};
  ram_789 = _RAND_791[7:0];
  _RAND_792 = {1{`RANDOM}};
  ram_790 = _RAND_792[7:0];
  _RAND_793 = {1{`RANDOM}};
  ram_791 = _RAND_793[7:0];
  _RAND_794 = {1{`RANDOM}};
  ram_792 = _RAND_794[7:0];
  _RAND_795 = {1{`RANDOM}};
  ram_793 = _RAND_795[7:0];
  _RAND_796 = {1{`RANDOM}};
  ram_794 = _RAND_796[7:0];
  _RAND_797 = {1{`RANDOM}};
  ram_795 = _RAND_797[7:0];
  _RAND_798 = {1{`RANDOM}};
  ram_796 = _RAND_798[7:0];
  _RAND_799 = {1{`RANDOM}};
  ram_797 = _RAND_799[7:0];
  _RAND_800 = {1{`RANDOM}};
  ram_798 = _RAND_800[7:0];
  _RAND_801 = {1{`RANDOM}};
  ram_799 = _RAND_801[7:0];
  _RAND_802 = {1{`RANDOM}};
  ram_800 = _RAND_802[7:0];
  _RAND_803 = {1{`RANDOM}};
  ram_801 = _RAND_803[7:0];
  _RAND_804 = {1{`RANDOM}};
  ram_802 = _RAND_804[7:0];
  _RAND_805 = {1{`RANDOM}};
  ram_803 = _RAND_805[7:0];
  _RAND_806 = {1{`RANDOM}};
  ram_804 = _RAND_806[7:0];
  _RAND_807 = {1{`RANDOM}};
  ram_805 = _RAND_807[7:0];
  _RAND_808 = {1{`RANDOM}};
  ram_806 = _RAND_808[7:0];
  _RAND_809 = {1{`RANDOM}};
  ram_807 = _RAND_809[7:0];
  _RAND_810 = {1{`RANDOM}};
  ram_808 = _RAND_810[7:0];
  _RAND_811 = {1{`RANDOM}};
  ram_809 = _RAND_811[7:0];
  _RAND_812 = {1{`RANDOM}};
  ram_810 = _RAND_812[7:0];
  _RAND_813 = {1{`RANDOM}};
  ram_811 = _RAND_813[7:0];
  _RAND_814 = {1{`RANDOM}};
  ram_812 = _RAND_814[7:0];
  _RAND_815 = {1{`RANDOM}};
  ram_813 = _RAND_815[7:0];
  _RAND_816 = {1{`RANDOM}};
  ram_814 = _RAND_816[7:0];
  _RAND_817 = {1{`RANDOM}};
  ram_815 = _RAND_817[7:0];
  _RAND_818 = {1{`RANDOM}};
  ram_816 = _RAND_818[7:0];
  _RAND_819 = {1{`RANDOM}};
  ram_817 = _RAND_819[7:0];
  _RAND_820 = {1{`RANDOM}};
  ram_818 = _RAND_820[7:0];
  _RAND_821 = {1{`RANDOM}};
  ram_819 = _RAND_821[7:0];
  _RAND_822 = {1{`RANDOM}};
  ram_820 = _RAND_822[7:0];
  _RAND_823 = {1{`RANDOM}};
  ram_821 = _RAND_823[7:0];
  _RAND_824 = {1{`RANDOM}};
  ram_822 = _RAND_824[7:0];
  _RAND_825 = {1{`RANDOM}};
  ram_823 = _RAND_825[7:0];
  _RAND_826 = {1{`RANDOM}};
  ram_824 = _RAND_826[7:0];
  _RAND_827 = {1{`RANDOM}};
  ram_825 = _RAND_827[7:0];
  _RAND_828 = {1{`RANDOM}};
  ram_826 = _RAND_828[7:0];
  _RAND_829 = {1{`RANDOM}};
  ram_827 = _RAND_829[7:0];
  _RAND_830 = {1{`RANDOM}};
  ram_828 = _RAND_830[7:0];
  _RAND_831 = {1{`RANDOM}};
  ram_829 = _RAND_831[7:0];
  _RAND_832 = {1{`RANDOM}};
  ram_830 = _RAND_832[7:0];
  _RAND_833 = {1{`RANDOM}};
  ram_831 = _RAND_833[7:0];
  _RAND_834 = {1{`RANDOM}};
  ram_832 = _RAND_834[7:0];
  _RAND_835 = {1{`RANDOM}};
  ram_833 = _RAND_835[7:0];
  _RAND_836 = {1{`RANDOM}};
  ram_834 = _RAND_836[7:0];
  _RAND_837 = {1{`RANDOM}};
  ram_835 = _RAND_837[7:0];
  _RAND_838 = {1{`RANDOM}};
  ram_836 = _RAND_838[7:0];
  _RAND_839 = {1{`RANDOM}};
  ram_837 = _RAND_839[7:0];
  _RAND_840 = {1{`RANDOM}};
  ram_838 = _RAND_840[7:0];
  _RAND_841 = {1{`RANDOM}};
  ram_839 = _RAND_841[7:0];
  _RAND_842 = {1{`RANDOM}};
  ram_840 = _RAND_842[7:0];
  _RAND_843 = {1{`RANDOM}};
  ram_841 = _RAND_843[7:0];
  _RAND_844 = {1{`RANDOM}};
  ram_842 = _RAND_844[7:0];
  _RAND_845 = {1{`RANDOM}};
  ram_843 = _RAND_845[7:0];
  _RAND_846 = {1{`RANDOM}};
  ram_844 = _RAND_846[7:0];
  _RAND_847 = {1{`RANDOM}};
  ram_845 = _RAND_847[7:0];
  _RAND_848 = {1{`RANDOM}};
  ram_846 = _RAND_848[7:0];
  _RAND_849 = {1{`RANDOM}};
  ram_847 = _RAND_849[7:0];
  _RAND_850 = {1{`RANDOM}};
  ram_848 = _RAND_850[7:0];
  _RAND_851 = {1{`RANDOM}};
  ram_849 = _RAND_851[7:0];
  _RAND_852 = {1{`RANDOM}};
  ram_850 = _RAND_852[7:0];
  _RAND_853 = {1{`RANDOM}};
  ram_851 = _RAND_853[7:0];
  _RAND_854 = {1{`RANDOM}};
  ram_852 = _RAND_854[7:0];
  _RAND_855 = {1{`RANDOM}};
  ram_853 = _RAND_855[7:0];
  _RAND_856 = {1{`RANDOM}};
  ram_854 = _RAND_856[7:0];
  _RAND_857 = {1{`RANDOM}};
  ram_855 = _RAND_857[7:0];
  _RAND_858 = {1{`RANDOM}};
  ram_856 = _RAND_858[7:0];
  _RAND_859 = {1{`RANDOM}};
  ram_857 = _RAND_859[7:0];
  _RAND_860 = {1{`RANDOM}};
  ram_858 = _RAND_860[7:0];
  _RAND_861 = {1{`RANDOM}};
  ram_859 = _RAND_861[7:0];
  _RAND_862 = {1{`RANDOM}};
  ram_860 = _RAND_862[7:0];
  _RAND_863 = {1{`RANDOM}};
  ram_861 = _RAND_863[7:0];
  _RAND_864 = {1{`RANDOM}};
  ram_862 = _RAND_864[7:0];
  _RAND_865 = {1{`RANDOM}};
  ram_863 = _RAND_865[7:0];
  _RAND_866 = {1{`RANDOM}};
  ram_864 = _RAND_866[7:0];
  _RAND_867 = {1{`RANDOM}};
  ram_865 = _RAND_867[7:0];
  _RAND_868 = {1{`RANDOM}};
  ram_866 = _RAND_868[7:0];
  _RAND_869 = {1{`RANDOM}};
  ram_867 = _RAND_869[7:0];
  _RAND_870 = {1{`RANDOM}};
  ram_868 = _RAND_870[7:0];
  _RAND_871 = {1{`RANDOM}};
  ram_869 = _RAND_871[7:0];
  _RAND_872 = {1{`RANDOM}};
  ram_870 = _RAND_872[7:0];
  _RAND_873 = {1{`RANDOM}};
  ram_871 = _RAND_873[7:0];
  _RAND_874 = {1{`RANDOM}};
  ram_872 = _RAND_874[7:0];
  _RAND_875 = {1{`RANDOM}};
  ram_873 = _RAND_875[7:0];
  _RAND_876 = {1{`RANDOM}};
  ram_874 = _RAND_876[7:0];
  _RAND_877 = {1{`RANDOM}};
  ram_875 = _RAND_877[7:0];
  _RAND_878 = {1{`RANDOM}};
  ram_876 = _RAND_878[7:0];
  _RAND_879 = {1{`RANDOM}};
  ram_877 = _RAND_879[7:0];
  _RAND_880 = {1{`RANDOM}};
  ram_878 = _RAND_880[7:0];
  _RAND_881 = {1{`RANDOM}};
  ram_879 = _RAND_881[7:0];
  _RAND_882 = {1{`RANDOM}};
  ram_880 = _RAND_882[7:0];
  _RAND_883 = {1{`RANDOM}};
  ram_881 = _RAND_883[7:0];
  _RAND_884 = {1{`RANDOM}};
  ram_882 = _RAND_884[7:0];
  _RAND_885 = {1{`RANDOM}};
  ram_883 = _RAND_885[7:0];
  _RAND_886 = {1{`RANDOM}};
  ram_884 = _RAND_886[7:0];
  _RAND_887 = {1{`RANDOM}};
  ram_885 = _RAND_887[7:0];
  _RAND_888 = {1{`RANDOM}};
  ram_886 = _RAND_888[7:0];
  _RAND_889 = {1{`RANDOM}};
  ram_887 = _RAND_889[7:0];
  _RAND_890 = {1{`RANDOM}};
  ram_888 = _RAND_890[7:0];
  _RAND_891 = {1{`RANDOM}};
  ram_889 = _RAND_891[7:0];
  _RAND_892 = {1{`RANDOM}};
  ram_890 = _RAND_892[7:0];
  _RAND_893 = {1{`RANDOM}};
  ram_891 = _RAND_893[7:0];
  _RAND_894 = {1{`RANDOM}};
  ram_892 = _RAND_894[7:0];
  _RAND_895 = {1{`RANDOM}};
  ram_893 = _RAND_895[7:0];
  _RAND_896 = {1{`RANDOM}};
  ram_894 = _RAND_896[7:0];
  _RAND_897 = {1{`RANDOM}};
  ram_895 = _RAND_897[7:0];
  _RAND_898 = {1{`RANDOM}};
  ram_896 = _RAND_898[7:0];
  _RAND_899 = {1{`RANDOM}};
  ram_897 = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  ram_898 = _RAND_900[7:0];
  _RAND_901 = {1{`RANDOM}};
  ram_899 = _RAND_901[7:0];
  _RAND_902 = {1{`RANDOM}};
  ram_900 = _RAND_902[7:0];
  _RAND_903 = {1{`RANDOM}};
  ram_901 = _RAND_903[7:0];
  _RAND_904 = {1{`RANDOM}};
  ram_902 = _RAND_904[7:0];
  _RAND_905 = {1{`RANDOM}};
  ram_903 = _RAND_905[7:0];
  _RAND_906 = {1{`RANDOM}};
  ram_904 = _RAND_906[7:0];
  _RAND_907 = {1{`RANDOM}};
  ram_905 = _RAND_907[7:0];
  _RAND_908 = {1{`RANDOM}};
  ram_906 = _RAND_908[7:0];
  _RAND_909 = {1{`RANDOM}};
  ram_907 = _RAND_909[7:0];
  _RAND_910 = {1{`RANDOM}};
  ram_908 = _RAND_910[7:0];
  _RAND_911 = {1{`RANDOM}};
  ram_909 = _RAND_911[7:0];
  _RAND_912 = {1{`RANDOM}};
  ram_910 = _RAND_912[7:0];
  _RAND_913 = {1{`RANDOM}};
  ram_911 = _RAND_913[7:0];
  _RAND_914 = {1{`RANDOM}};
  ram_912 = _RAND_914[7:0];
  _RAND_915 = {1{`RANDOM}};
  ram_913 = _RAND_915[7:0];
  _RAND_916 = {1{`RANDOM}};
  ram_914 = _RAND_916[7:0];
  _RAND_917 = {1{`RANDOM}};
  ram_915 = _RAND_917[7:0];
  _RAND_918 = {1{`RANDOM}};
  ram_916 = _RAND_918[7:0];
  _RAND_919 = {1{`RANDOM}};
  ram_917 = _RAND_919[7:0];
  _RAND_920 = {1{`RANDOM}};
  ram_918 = _RAND_920[7:0];
  _RAND_921 = {1{`RANDOM}};
  ram_919 = _RAND_921[7:0];
  _RAND_922 = {1{`RANDOM}};
  ram_920 = _RAND_922[7:0];
  _RAND_923 = {1{`RANDOM}};
  ram_921 = _RAND_923[7:0];
  _RAND_924 = {1{`RANDOM}};
  ram_922 = _RAND_924[7:0];
  _RAND_925 = {1{`RANDOM}};
  ram_923 = _RAND_925[7:0];
  _RAND_926 = {1{`RANDOM}};
  ram_924 = _RAND_926[7:0];
  _RAND_927 = {1{`RANDOM}};
  ram_925 = _RAND_927[7:0];
  _RAND_928 = {1{`RANDOM}};
  ram_926 = _RAND_928[7:0];
  _RAND_929 = {1{`RANDOM}};
  ram_927 = _RAND_929[7:0];
  _RAND_930 = {1{`RANDOM}};
  ram_928 = _RAND_930[7:0];
  _RAND_931 = {1{`RANDOM}};
  ram_929 = _RAND_931[7:0];
  _RAND_932 = {1{`RANDOM}};
  ram_930 = _RAND_932[7:0];
  _RAND_933 = {1{`RANDOM}};
  ram_931 = _RAND_933[7:0];
  _RAND_934 = {1{`RANDOM}};
  ram_932 = _RAND_934[7:0];
  _RAND_935 = {1{`RANDOM}};
  ram_933 = _RAND_935[7:0];
  _RAND_936 = {1{`RANDOM}};
  ram_934 = _RAND_936[7:0];
  _RAND_937 = {1{`RANDOM}};
  ram_935 = _RAND_937[7:0];
  _RAND_938 = {1{`RANDOM}};
  ram_936 = _RAND_938[7:0];
  _RAND_939 = {1{`RANDOM}};
  ram_937 = _RAND_939[7:0];
  _RAND_940 = {1{`RANDOM}};
  ram_938 = _RAND_940[7:0];
  _RAND_941 = {1{`RANDOM}};
  ram_939 = _RAND_941[7:0];
  _RAND_942 = {1{`RANDOM}};
  ram_940 = _RAND_942[7:0];
  _RAND_943 = {1{`RANDOM}};
  ram_941 = _RAND_943[7:0];
  _RAND_944 = {1{`RANDOM}};
  ram_942 = _RAND_944[7:0];
  _RAND_945 = {1{`RANDOM}};
  ram_943 = _RAND_945[7:0];
  _RAND_946 = {1{`RANDOM}};
  ram_944 = _RAND_946[7:0];
  _RAND_947 = {1{`RANDOM}};
  ram_945 = _RAND_947[7:0];
  _RAND_948 = {1{`RANDOM}};
  ram_946 = _RAND_948[7:0];
  _RAND_949 = {1{`RANDOM}};
  ram_947 = _RAND_949[7:0];
  _RAND_950 = {1{`RANDOM}};
  ram_948 = _RAND_950[7:0];
  _RAND_951 = {1{`RANDOM}};
  ram_949 = _RAND_951[7:0];
  _RAND_952 = {1{`RANDOM}};
  ram_950 = _RAND_952[7:0];
  _RAND_953 = {1{`RANDOM}};
  ram_951 = _RAND_953[7:0];
  _RAND_954 = {1{`RANDOM}};
  ram_952 = _RAND_954[7:0];
  _RAND_955 = {1{`RANDOM}};
  ram_953 = _RAND_955[7:0];
  _RAND_956 = {1{`RANDOM}};
  ram_954 = _RAND_956[7:0];
  _RAND_957 = {1{`RANDOM}};
  ram_955 = _RAND_957[7:0];
  _RAND_958 = {1{`RANDOM}};
  ram_956 = _RAND_958[7:0];
  _RAND_959 = {1{`RANDOM}};
  ram_957 = _RAND_959[7:0];
  _RAND_960 = {1{`RANDOM}};
  ram_958 = _RAND_960[7:0];
  _RAND_961 = {1{`RANDOM}};
  ram_959 = _RAND_961[7:0];
  _RAND_962 = {1{`RANDOM}};
  ram_960 = _RAND_962[7:0];
  _RAND_963 = {1{`RANDOM}};
  ram_961 = _RAND_963[7:0];
  _RAND_964 = {1{`RANDOM}};
  ram_962 = _RAND_964[7:0];
  _RAND_965 = {1{`RANDOM}};
  ram_963 = _RAND_965[7:0];
  _RAND_966 = {1{`RANDOM}};
  ram_964 = _RAND_966[7:0];
  _RAND_967 = {1{`RANDOM}};
  ram_965 = _RAND_967[7:0];
  _RAND_968 = {1{`RANDOM}};
  ram_966 = _RAND_968[7:0];
  _RAND_969 = {1{`RANDOM}};
  ram_967 = _RAND_969[7:0];
  _RAND_970 = {1{`RANDOM}};
  ram_968 = _RAND_970[7:0];
  _RAND_971 = {1{`RANDOM}};
  ram_969 = _RAND_971[7:0];
  _RAND_972 = {1{`RANDOM}};
  ram_970 = _RAND_972[7:0];
  _RAND_973 = {1{`RANDOM}};
  ram_971 = _RAND_973[7:0];
  _RAND_974 = {1{`RANDOM}};
  ram_972 = _RAND_974[7:0];
  _RAND_975 = {1{`RANDOM}};
  ram_973 = _RAND_975[7:0];
  _RAND_976 = {1{`RANDOM}};
  ram_974 = _RAND_976[7:0];
  _RAND_977 = {1{`RANDOM}};
  ram_975 = _RAND_977[7:0];
  _RAND_978 = {1{`RANDOM}};
  ram_976 = _RAND_978[7:0];
  _RAND_979 = {1{`RANDOM}};
  ram_977 = _RAND_979[7:0];
  _RAND_980 = {1{`RANDOM}};
  ram_978 = _RAND_980[7:0];
  _RAND_981 = {1{`RANDOM}};
  ram_979 = _RAND_981[7:0];
  _RAND_982 = {1{`RANDOM}};
  ram_980 = _RAND_982[7:0];
  _RAND_983 = {1{`RANDOM}};
  ram_981 = _RAND_983[7:0];
  _RAND_984 = {1{`RANDOM}};
  ram_982 = _RAND_984[7:0];
  _RAND_985 = {1{`RANDOM}};
  ram_983 = _RAND_985[7:0];
  _RAND_986 = {1{`RANDOM}};
  ram_984 = _RAND_986[7:0];
  _RAND_987 = {1{`RANDOM}};
  ram_985 = _RAND_987[7:0];
  _RAND_988 = {1{`RANDOM}};
  ram_986 = _RAND_988[7:0];
  _RAND_989 = {1{`RANDOM}};
  ram_987 = _RAND_989[7:0];
  _RAND_990 = {1{`RANDOM}};
  ram_988 = _RAND_990[7:0];
  _RAND_991 = {1{`RANDOM}};
  ram_989 = _RAND_991[7:0];
  _RAND_992 = {1{`RANDOM}};
  ram_990 = _RAND_992[7:0];
  _RAND_993 = {1{`RANDOM}};
  ram_991 = _RAND_993[7:0];
  _RAND_994 = {1{`RANDOM}};
  ram_992 = _RAND_994[7:0];
  _RAND_995 = {1{`RANDOM}};
  ram_993 = _RAND_995[7:0];
  _RAND_996 = {1{`RANDOM}};
  ram_994 = _RAND_996[7:0];
  _RAND_997 = {1{`RANDOM}};
  ram_995 = _RAND_997[7:0];
  _RAND_998 = {1{`RANDOM}};
  ram_996 = _RAND_998[7:0];
  _RAND_999 = {1{`RANDOM}};
  ram_997 = _RAND_999[7:0];
  _RAND_1000 = {1{`RANDOM}};
  ram_998 = _RAND_1000[7:0];
  _RAND_1001 = {1{`RANDOM}};
  ram_999 = _RAND_1001[7:0];
  _RAND_1002 = {1{`RANDOM}};
  ram_1000 = _RAND_1002[7:0];
  _RAND_1003 = {1{`RANDOM}};
  ram_1001 = _RAND_1003[7:0];
  _RAND_1004 = {1{`RANDOM}};
  ram_1002 = _RAND_1004[7:0];
  _RAND_1005 = {1{`RANDOM}};
  ram_1003 = _RAND_1005[7:0];
  _RAND_1006 = {1{`RANDOM}};
  ram_1004 = _RAND_1006[7:0];
  _RAND_1007 = {1{`RANDOM}};
  ram_1005 = _RAND_1007[7:0];
  _RAND_1008 = {1{`RANDOM}};
  ram_1006 = _RAND_1008[7:0];
  _RAND_1009 = {1{`RANDOM}};
  ram_1007 = _RAND_1009[7:0];
  _RAND_1010 = {1{`RANDOM}};
  ram_1008 = _RAND_1010[7:0];
  _RAND_1011 = {1{`RANDOM}};
  ram_1009 = _RAND_1011[7:0];
  _RAND_1012 = {1{`RANDOM}};
  ram_1010 = _RAND_1012[7:0];
  _RAND_1013 = {1{`RANDOM}};
  ram_1011 = _RAND_1013[7:0];
  _RAND_1014 = {1{`RANDOM}};
  ram_1012 = _RAND_1014[7:0];
  _RAND_1015 = {1{`RANDOM}};
  ram_1013 = _RAND_1015[7:0];
  _RAND_1016 = {1{`RANDOM}};
  ram_1014 = _RAND_1016[7:0];
  _RAND_1017 = {1{`RANDOM}};
  ram_1015 = _RAND_1017[7:0];
  _RAND_1018 = {1{`RANDOM}};
  ram_1016 = _RAND_1018[7:0];
  _RAND_1019 = {1{`RANDOM}};
  ram_1017 = _RAND_1019[7:0];
  _RAND_1020 = {1{`RANDOM}};
  ram_1018 = _RAND_1020[7:0];
  _RAND_1021 = {1{`RANDOM}};
  ram_1019 = _RAND_1021[7:0];
  _RAND_1022 = {1{`RANDOM}};
  ram_1020 = _RAND_1022[7:0];
  _RAND_1023 = {1{`RANDOM}};
  ram_1021 = _RAND_1023[7:0];
  _RAND_1024 = {1{`RANDOM}};
  ram_1022 = _RAND_1024[7:0];
  _RAND_1025 = {1{`RANDOM}};
  ram_1023 = _RAND_1025[7:0];
  _RAND_1026 = {1{`RANDOM}};
  ram_1024 = _RAND_1026[7:0];
  _RAND_1027 = {1{`RANDOM}};
  ram_1025 = _RAND_1027[7:0];
  _RAND_1028 = {1{`RANDOM}};
  ram_1026 = _RAND_1028[7:0];
  _RAND_1029 = {1{`RANDOM}};
  ram_1027 = _RAND_1029[7:0];
  _RAND_1030 = {1{`RANDOM}};
  ram_1028 = _RAND_1030[7:0];
  _RAND_1031 = {1{`RANDOM}};
  ram_1029 = _RAND_1031[7:0];
  _RAND_1032 = {1{`RANDOM}};
  ram_1030 = _RAND_1032[7:0];
  _RAND_1033 = {1{`RANDOM}};
  ram_1031 = _RAND_1033[7:0];
  _RAND_1034 = {1{`RANDOM}};
  ram_1032 = _RAND_1034[7:0];
  _RAND_1035 = {1{`RANDOM}};
  ram_1033 = _RAND_1035[7:0];
  _RAND_1036 = {1{`RANDOM}};
  ram_1034 = _RAND_1036[7:0];
  _RAND_1037 = {1{`RANDOM}};
  ram_1035 = _RAND_1037[7:0];
  _RAND_1038 = {1{`RANDOM}};
  ram_1036 = _RAND_1038[7:0];
  _RAND_1039 = {1{`RANDOM}};
  ram_1037 = _RAND_1039[7:0];
  _RAND_1040 = {1{`RANDOM}};
  ram_1038 = _RAND_1040[7:0];
  _RAND_1041 = {1{`RANDOM}};
  ram_1039 = _RAND_1041[7:0];
  _RAND_1042 = {1{`RANDOM}};
  ram_1040 = _RAND_1042[7:0];
  _RAND_1043 = {1{`RANDOM}};
  ram_1041 = _RAND_1043[7:0];
  _RAND_1044 = {1{`RANDOM}};
  ram_1042 = _RAND_1044[7:0];
  _RAND_1045 = {1{`RANDOM}};
  ram_1043 = _RAND_1045[7:0];
  _RAND_1046 = {1{`RANDOM}};
  ram_1044 = _RAND_1046[7:0];
  _RAND_1047 = {1{`RANDOM}};
  ram_1045 = _RAND_1047[7:0];
  _RAND_1048 = {1{`RANDOM}};
  ram_1046 = _RAND_1048[7:0];
  _RAND_1049 = {1{`RANDOM}};
  ram_1047 = _RAND_1049[7:0];
  _RAND_1050 = {1{`RANDOM}};
  ram_1048 = _RAND_1050[7:0];
  _RAND_1051 = {1{`RANDOM}};
  ram_1049 = _RAND_1051[7:0];
  _RAND_1052 = {1{`RANDOM}};
  ram_1050 = _RAND_1052[7:0];
  _RAND_1053 = {1{`RANDOM}};
  ram_1051 = _RAND_1053[7:0];
  _RAND_1054 = {1{`RANDOM}};
  ram_1052 = _RAND_1054[7:0];
  _RAND_1055 = {1{`RANDOM}};
  ram_1053 = _RAND_1055[7:0];
  _RAND_1056 = {1{`RANDOM}};
  ram_1054 = _RAND_1056[7:0];
  _RAND_1057 = {1{`RANDOM}};
  ram_1055 = _RAND_1057[7:0];
  _RAND_1058 = {1{`RANDOM}};
  ram_1056 = _RAND_1058[7:0];
  _RAND_1059 = {1{`RANDOM}};
  ram_1057 = _RAND_1059[7:0];
  _RAND_1060 = {1{`RANDOM}};
  ram_1058 = _RAND_1060[7:0];
  _RAND_1061 = {1{`RANDOM}};
  ram_1059 = _RAND_1061[7:0];
  _RAND_1062 = {1{`RANDOM}};
  ram_1060 = _RAND_1062[7:0];
  _RAND_1063 = {1{`RANDOM}};
  ram_1061 = _RAND_1063[7:0];
  _RAND_1064 = {1{`RANDOM}};
  ram_1062 = _RAND_1064[7:0];
  _RAND_1065 = {1{`RANDOM}};
  ram_1063 = _RAND_1065[7:0];
  _RAND_1066 = {1{`RANDOM}};
  ram_1064 = _RAND_1066[7:0];
  _RAND_1067 = {1{`RANDOM}};
  ram_1065 = _RAND_1067[7:0];
  _RAND_1068 = {1{`RANDOM}};
  ram_1066 = _RAND_1068[7:0];
  _RAND_1069 = {1{`RANDOM}};
  ram_1067 = _RAND_1069[7:0];
  _RAND_1070 = {1{`RANDOM}};
  ram_1068 = _RAND_1070[7:0];
  _RAND_1071 = {1{`RANDOM}};
  ram_1069 = _RAND_1071[7:0];
  _RAND_1072 = {1{`RANDOM}};
  ram_1070 = _RAND_1072[7:0];
  _RAND_1073 = {1{`RANDOM}};
  ram_1071 = _RAND_1073[7:0];
  _RAND_1074 = {1{`RANDOM}};
  ram_1072 = _RAND_1074[7:0];
  _RAND_1075 = {1{`RANDOM}};
  ram_1073 = _RAND_1075[7:0];
  _RAND_1076 = {1{`RANDOM}};
  ram_1074 = _RAND_1076[7:0];
  _RAND_1077 = {1{`RANDOM}};
  ram_1075 = _RAND_1077[7:0];
  _RAND_1078 = {1{`RANDOM}};
  ram_1076 = _RAND_1078[7:0];
  _RAND_1079 = {1{`RANDOM}};
  ram_1077 = _RAND_1079[7:0];
  _RAND_1080 = {1{`RANDOM}};
  ram_1078 = _RAND_1080[7:0];
  _RAND_1081 = {1{`RANDOM}};
  ram_1079 = _RAND_1081[7:0];
  _RAND_1082 = {1{`RANDOM}};
  ram_1080 = _RAND_1082[7:0];
  _RAND_1083 = {1{`RANDOM}};
  ram_1081 = _RAND_1083[7:0];
  _RAND_1084 = {1{`RANDOM}};
  ram_1082 = _RAND_1084[7:0];
  _RAND_1085 = {1{`RANDOM}};
  ram_1083 = _RAND_1085[7:0];
  _RAND_1086 = {1{`RANDOM}};
  ram_1084 = _RAND_1086[7:0];
  _RAND_1087 = {1{`RANDOM}};
  ram_1085 = _RAND_1087[7:0];
  _RAND_1088 = {1{`RANDOM}};
  ram_1086 = _RAND_1088[7:0];
  _RAND_1089 = {1{`RANDOM}};
  ram_1087 = _RAND_1089[7:0];
  _RAND_1090 = {1{`RANDOM}};
  ram_1088 = _RAND_1090[7:0];
  _RAND_1091 = {1{`RANDOM}};
  ram_1089 = _RAND_1091[7:0];
  _RAND_1092 = {1{`RANDOM}};
  ram_1090 = _RAND_1092[7:0];
  _RAND_1093 = {1{`RANDOM}};
  ram_1091 = _RAND_1093[7:0];
  _RAND_1094 = {1{`RANDOM}};
  ram_1092 = _RAND_1094[7:0];
  _RAND_1095 = {1{`RANDOM}};
  ram_1093 = _RAND_1095[7:0];
  _RAND_1096 = {1{`RANDOM}};
  ram_1094 = _RAND_1096[7:0];
  _RAND_1097 = {1{`RANDOM}};
  ram_1095 = _RAND_1097[7:0];
  _RAND_1098 = {1{`RANDOM}};
  ram_1096 = _RAND_1098[7:0];
  _RAND_1099 = {1{`RANDOM}};
  ram_1097 = _RAND_1099[7:0];
  _RAND_1100 = {1{`RANDOM}};
  ram_1098 = _RAND_1100[7:0];
  _RAND_1101 = {1{`RANDOM}};
  ram_1099 = _RAND_1101[7:0];
  _RAND_1102 = {1{`RANDOM}};
  ram_1100 = _RAND_1102[7:0];
  _RAND_1103 = {1{`RANDOM}};
  ram_1101 = _RAND_1103[7:0];
  _RAND_1104 = {1{`RANDOM}};
  ram_1102 = _RAND_1104[7:0];
  _RAND_1105 = {1{`RANDOM}};
  ram_1103 = _RAND_1105[7:0];
  _RAND_1106 = {1{`RANDOM}};
  ram_1104 = _RAND_1106[7:0];
  _RAND_1107 = {1{`RANDOM}};
  ram_1105 = _RAND_1107[7:0];
  _RAND_1108 = {1{`RANDOM}};
  ram_1106 = _RAND_1108[7:0];
  _RAND_1109 = {1{`RANDOM}};
  ram_1107 = _RAND_1109[7:0];
  _RAND_1110 = {1{`RANDOM}};
  ram_1108 = _RAND_1110[7:0];
  _RAND_1111 = {1{`RANDOM}};
  ram_1109 = _RAND_1111[7:0];
  _RAND_1112 = {1{`RANDOM}};
  ram_1110 = _RAND_1112[7:0];
  _RAND_1113 = {1{`RANDOM}};
  ram_1111 = _RAND_1113[7:0];
  _RAND_1114 = {1{`RANDOM}};
  ram_1112 = _RAND_1114[7:0];
  _RAND_1115 = {1{`RANDOM}};
  ram_1113 = _RAND_1115[7:0];
  _RAND_1116 = {1{`RANDOM}};
  ram_1114 = _RAND_1116[7:0];
  _RAND_1117 = {1{`RANDOM}};
  ram_1115 = _RAND_1117[7:0];
  _RAND_1118 = {1{`RANDOM}};
  ram_1116 = _RAND_1118[7:0];
  _RAND_1119 = {1{`RANDOM}};
  ram_1117 = _RAND_1119[7:0];
  _RAND_1120 = {1{`RANDOM}};
  ram_1118 = _RAND_1120[7:0];
  _RAND_1121 = {1{`RANDOM}};
  ram_1119 = _RAND_1121[7:0];
  _RAND_1122 = {1{`RANDOM}};
  ram_1120 = _RAND_1122[7:0];
  _RAND_1123 = {1{`RANDOM}};
  ram_1121 = _RAND_1123[7:0];
  _RAND_1124 = {1{`RANDOM}};
  ram_1122 = _RAND_1124[7:0];
  _RAND_1125 = {1{`RANDOM}};
  ram_1123 = _RAND_1125[7:0];
  _RAND_1126 = {1{`RANDOM}};
  ram_1124 = _RAND_1126[7:0];
  _RAND_1127 = {1{`RANDOM}};
  ram_1125 = _RAND_1127[7:0];
  _RAND_1128 = {1{`RANDOM}};
  ram_1126 = _RAND_1128[7:0];
  _RAND_1129 = {1{`RANDOM}};
  ram_1127 = _RAND_1129[7:0];
  _RAND_1130 = {1{`RANDOM}};
  ram_1128 = _RAND_1130[7:0];
  _RAND_1131 = {1{`RANDOM}};
  ram_1129 = _RAND_1131[7:0];
  _RAND_1132 = {1{`RANDOM}};
  ram_1130 = _RAND_1132[7:0];
  _RAND_1133 = {1{`RANDOM}};
  ram_1131 = _RAND_1133[7:0];
  _RAND_1134 = {1{`RANDOM}};
  ram_1132 = _RAND_1134[7:0];
  _RAND_1135 = {1{`RANDOM}};
  ram_1133 = _RAND_1135[7:0];
  _RAND_1136 = {1{`RANDOM}};
  ram_1134 = _RAND_1136[7:0];
  _RAND_1137 = {1{`RANDOM}};
  ram_1135 = _RAND_1137[7:0];
  _RAND_1138 = {1{`RANDOM}};
  ram_1136 = _RAND_1138[7:0];
  _RAND_1139 = {1{`RANDOM}};
  ram_1137 = _RAND_1139[7:0];
  _RAND_1140 = {1{`RANDOM}};
  ram_1138 = _RAND_1140[7:0];
  _RAND_1141 = {1{`RANDOM}};
  ram_1139 = _RAND_1141[7:0];
  _RAND_1142 = {1{`RANDOM}};
  ram_1140 = _RAND_1142[7:0];
  _RAND_1143 = {1{`RANDOM}};
  ram_1141 = _RAND_1143[7:0];
  _RAND_1144 = {1{`RANDOM}};
  ram_1142 = _RAND_1144[7:0];
  _RAND_1145 = {1{`RANDOM}};
  ram_1143 = _RAND_1145[7:0];
  _RAND_1146 = {1{`RANDOM}};
  ram_1144 = _RAND_1146[7:0];
  _RAND_1147 = {1{`RANDOM}};
  ram_1145 = _RAND_1147[7:0];
  _RAND_1148 = {1{`RANDOM}};
  ram_1146 = _RAND_1148[7:0];
  _RAND_1149 = {1{`RANDOM}};
  ram_1147 = _RAND_1149[7:0];
  _RAND_1150 = {1{`RANDOM}};
  ram_1148 = _RAND_1150[7:0];
  _RAND_1151 = {1{`RANDOM}};
  ram_1149 = _RAND_1151[7:0];
  _RAND_1152 = {1{`RANDOM}};
  ram_1150 = _RAND_1152[7:0];
  _RAND_1153 = {1{`RANDOM}};
  ram_1151 = _RAND_1153[7:0];
  _RAND_1154 = {1{`RANDOM}};
  ram_1152 = _RAND_1154[7:0];
  _RAND_1155 = {1{`RANDOM}};
  ram_1153 = _RAND_1155[7:0];
  _RAND_1156 = {1{`RANDOM}};
  ram_1154 = _RAND_1156[7:0];
  _RAND_1157 = {1{`RANDOM}};
  ram_1155 = _RAND_1157[7:0];
  _RAND_1158 = {1{`RANDOM}};
  ram_1156 = _RAND_1158[7:0];
  _RAND_1159 = {1{`RANDOM}};
  ram_1157 = _RAND_1159[7:0];
  _RAND_1160 = {1{`RANDOM}};
  ram_1158 = _RAND_1160[7:0];
  _RAND_1161 = {1{`RANDOM}};
  ram_1159 = _RAND_1161[7:0];
  _RAND_1162 = {1{`RANDOM}};
  ram_1160 = _RAND_1162[7:0];
  _RAND_1163 = {1{`RANDOM}};
  ram_1161 = _RAND_1163[7:0];
  _RAND_1164 = {1{`RANDOM}};
  ram_1162 = _RAND_1164[7:0];
  _RAND_1165 = {1{`RANDOM}};
  ram_1163 = _RAND_1165[7:0];
  _RAND_1166 = {1{`RANDOM}};
  ram_1164 = _RAND_1166[7:0];
  _RAND_1167 = {1{`RANDOM}};
  ram_1165 = _RAND_1167[7:0];
  _RAND_1168 = {1{`RANDOM}};
  ram_1166 = _RAND_1168[7:0];
  _RAND_1169 = {1{`RANDOM}};
  ram_1167 = _RAND_1169[7:0];
  _RAND_1170 = {1{`RANDOM}};
  ram_1168 = _RAND_1170[7:0];
  _RAND_1171 = {1{`RANDOM}};
  ram_1169 = _RAND_1171[7:0];
  _RAND_1172 = {1{`RANDOM}};
  ram_1170 = _RAND_1172[7:0];
  _RAND_1173 = {1{`RANDOM}};
  ram_1171 = _RAND_1173[7:0];
  _RAND_1174 = {1{`RANDOM}};
  ram_1172 = _RAND_1174[7:0];
  _RAND_1175 = {1{`RANDOM}};
  ram_1173 = _RAND_1175[7:0];
  _RAND_1176 = {1{`RANDOM}};
  ram_1174 = _RAND_1176[7:0];
  _RAND_1177 = {1{`RANDOM}};
  ram_1175 = _RAND_1177[7:0];
  _RAND_1178 = {1{`RANDOM}};
  ram_1176 = _RAND_1178[7:0];
  _RAND_1179 = {1{`RANDOM}};
  ram_1177 = _RAND_1179[7:0];
  _RAND_1180 = {1{`RANDOM}};
  ram_1178 = _RAND_1180[7:0];
  _RAND_1181 = {1{`RANDOM}};
  ram_1179 = _RAND_1181[7:0];
  _RAND_1182 = {1{`RANDOM}};
  ram_1180 = _RAND_1182[7:0];
  _RAND_1183 = {1{`RANDOM}};
  ram_1181 = _RAND_1183[7:0];
  _RAND_1184 = {1{`RANDOM}};
  ram_1182 = _RAND_1184[7:0];
  _RAND_1185 = {1{`RANDOM}};
  ram_1183 = _RAND_1185[7:0];
  _RAND_1186 = {1{`RANDOM}};
  ram_1184 = _RAND_1186[7:0];
  _RAND_1187 = {1{`RANDOM}};
  ram_1185 = _RAND_1187[7:0];
  _RAND_1188 = {1{`RANDOM}};
  ram_1186 = _RAND_1188[7:0];
  _RAND_1189 = {1{`RANDOM}};
  ram_1187 = _RAND_1189[7:0];
  _RAND_1190 = {1{`RANDOM}};
  ram_1188 = _RAND_1190[7:0];
  _RAND_1191 = {1{`RANDOM}};
  ram_1189 = _RAND_1191[7:0];
  _RAND_1192 = {1{`RANDOM}};
  ram_1190 = _RAND_1192[7:0];
  _RAND_1193 = {1{`RANDOM}};
  ram_1191 = _RAND_1193[7:0];
  _RAND_1194 = {1{`RANDOM}};
  ram_1192 = _RAND_1194[7:0];
  _RAND_1195 = {1{`RANDOM}};
  ram_1193 = _RAND_1195[7:0];
  _RAND_1196 = {1{`RANDOM}};
  ram_1194 = _RAND_1196[7:0];
  _RAND_1197 = {1{`RANDOM}};
  ram_1195 = _RAND_1197[7:0];
  _RAND_1198 = {1{`RANDOM}};
  ram_1196 = _RAND_1198[7:0];
  _RAND_1199 = {1{`RANDOM}};
  ram_1197 = _RAND_1199[7:0];
  _RAND_1200 = {1{`RANDOM}};
  ram_1198 = _RAND_1200[7:0];
  _RAND_1201 = {1{`RANDOM}};
  ram_1199 = _RAND_1201[7:0];
  _RAND_1202 = {1{`RANDOM}};
  ram_1200 = _RAND_1202[7:0];
  _RAND_1203 = {1{`RANDOM}};
  ram_1201 = _RAND_1203[7:0];
  _RAND_1204 = {1{`RANDOM}};
  ram_1202 = _RAND_1204[7:0];
  _RAND_1205 = {1{`RANDOM}};
  ram_1203 = _RAND_1205[7:0];
  _RAND_1206 = {1{`RANDOM}};
  ram_1204 = _RAND_1206[7:0];
  _RAND_1207 = {1{`RANDOM}};
  ram_1205 = _RAND_1207[7:0];
  _RAND_1208 = {1{`RANDOM}};
  ram_1206 = _RAND_1208[7:0];
  _RAND_1209 = {1{`RANDOM}};
  ram_1207 = _RAND_1209[7:0];
  _RAND_1210 = {1{`RANDOM}};
  ram_1208 = _RAND_1210[7:0];
  _RAND_1211 = {1{`RANDOM}};
  ram_1209 = _RAND_1211[7:0];
  _RAND_1212 = {1{`RANDOM}};
  ram_1210 = _RAND_1212[7:0];
  _RAND_1213 = {1{`RANDOM}};
  ram_1211 = _RAND_1213[7:0];
  _RAND_1214 = {1{`RANDOM}};
  ram_1212 = _RAND_1214[7:0];
  _RAND_1215 = {1{`RANDOM}};
  ram_1213 = _RAND_1215[7:0];
  _RAND_1216 = {1{`RANDOM}};
  ram_1214 = _RAND_1216[7:0];
  _RAND_1217 = {1{`RANDOM}};
  ram_1215 = _RAND_1217[7:0];
  _RAND_1218 = {1{`RANDOM}};
  ram_1216 = _RAND_1218[7:0];
  _RAND_1219 = {1{`RANDOM}};
  ram_1217 = _RAND_1219[7:0];
  _RAND_1220 = {1{`RANDOM}};
  ram_1218 = _RAND_1220[7:0];
  _RAND_1221 = {1{`RANDOM}};
  ram_1219 = _RAND_1221[7:0];
  _RAND_1222 = {1{`RANDOM}};
  ram_1220 = _RAND_1222[7:0];
  _RAND_1223 = {1{`RANDOM}};
  ram_1221 = _RAND_1223[7:0];
  _RAND_1224 = {1{`RANDOM}};
  ram_1222 = _RAND_1224[7:0];
  _RAND_1225 = {1{`RANDOM}};
  ram_1223 = _RAND_1225[7:0];
  _RAND_1226 = {1{`RANDOM}};
  ram_1224 = _RAND_1226[7:0];
  _RAND_1227 = {1{`RANDOM}};
  ram_1225 = _RAND_1227[7:0];
  _RAND_1228 = {1{`RANDOM}};
  ram_1226 = _RAND_1228[7:0];
  _RAND_1229 = {1{`RANDOM}};
  ram_1227 = _RAND_1229[7:0];
  _RAND_1230 = {1{`RANDOM}};
  ram_1228 = _RAND_1230[7:0];
  _RAND_1231 = {1{`RANDOM}};
  ram_1229 = _RAND_1231[7:0];
  _RAND_1232 = {1{`RANDOM}};
  ram_1230 = _RAND_1232[7:0];
  _RAND_1233 = {1{`RANDOM}};
  ram_1231 = _RAND_1233[7:0];
  _RAND_1234 = {1{`RANDOM}};
  ram_1232 = _RAND_1234[7:0];
  _RAND_1235 = {1{`RANDOM}};
  ram_1233 = _RAND_1235[7:0];
  _RAND_1236 = {1{`RANDOM}};
  ram_1234 = _RAND_1236[7:0];
  _RAND_1237 = {1{`RANDOM}};
  ram_1235 = _RAND_1237[7:0];
  _RAND_1238 = {1{`RANDOM}};
  ram_1236 = _RAND_1238[7:0];
  _RAND_1239 = {1{`RANDOM}};
  ram_1237 = _RAND_1239[7:0];
  _RAND_1240 = {1{`RANDOM}};
  ram_1238 = _RAND_1240[7:0];
  _RAND_1241 = {1{`RANDOM}};
  ram_1239 = _RAND_1241[7:0];
  _RAND_1242 = {1{`RANDOM}};
  ram_1240 = _RAND_1242[7:0];
  _RAND_1243 = {1{`RANDOM}};
  ram_1241 = _RAND_1243[7:0];
  _RAND_1244 = {1{`RANDOM}};
  ram_1242 = _RAND_1244[7:0];
  _RAND_1245 = {1{`RANDOM}};
  ram_1243 = _RAND_1245[7:0];
  _RAND_1246 = {1{`RANDOM}};
  ram_1244 = _RAND_1246[7:0];
  _RAND_1247 = {1{`RANDOM}};
  ram_1245 = _RAND_1247[7:0];
  _RAND_1248 = {1{`RANDOM}};
  ram_1246 = _RAND_1248[7:0];
  _RAND_1249 = {1{`RANDOM}};
  ram_1247 = _RAND_1249[7:0];
  _RAND_1250 = {1{`RANDOM}};
  ram_1248 = _RAND_1250[7:0];
  _RAND_1251 = {1{`RANDOM}};
  ram_1249 = _RAND_1251[7:0];
  _RAND_1252 = {1{`RANDOM}};
  ram_1250 = _RAND_1252[7:0];
  _RAND_1253 = {1{`RANDOM}};
  ram_1251 = _RAND_1253[7:0];
  _RAND_1254 = {1{`RANDOM}};
  ram_1252 = _RAND_1254[7:0];
  _RAND_1255 = {1{`RANDOM}};
  ram_1253 = _RAND_1255[7:0];
  _RAND_1256 = {1{`RANDOM}};
  ram_1254 = _RAND_1256[7:0];
  _RAND_1257 = {1{`RANDOM}};
  ram_1255 = _RAND_1257[7:0];
  _RAND_1258 = {1{`RANDOM}};
  ram_1256 = _RAND_1258[7:0];
  _RAND_1259 = {1{`RANDOM}};
  ram_1257 = _RAND_1259[7:0];
  _RAND_1260 = {1{`RANDOM}};
  ram_1258 = _RAND_1260[7:0];
  _RAND_1261 = {1{`RANDOM}};
  ram_1259 = _RAND_1261[7:0];
  _RAND_1262 = {1{`RANDOM}};
  ram_1260 = _RAND_1262[7:0];
  _RAND_1263 = {1{`RANDOM}};
  ram_1261 = _RAND_1263[7:0];
  _RAND_1264 = {1{`RANDOM}};
  ram_1262 = _RAND_1264[7:0];
  _RAND_1265 = {1{`RANDOM}};
  ram_1263 = _RAND_1265[7:0];
  _RAND_1266 = {1{`RANDOM}};
  ram_1264 = _RAND_1266[7:0];
  _RAND_1267 = {1{`RANDOM}};
  ram_1265 = _RAND_1267[7:0];
  _RAND_1268 = {1{`RANDOM}};
  ram_1266 = _RAND_1268[7:0];
  _RAND_1269 = {1{`RANDOM}};
  ram_1267 = _RAND_1269[7:0];
  _RAND_1270 = {1{`RANDOM}};
  ram_1268 = _RAND_1270[7:0];
  _RAND_1271 = {1{`RANDOM}};
  ram_1269 = _RAND_1271[7:0];
  _RAND_1272 = {1{`RANDOM}};
  ram_1270 = _RAND_1272[7:0];
  _RAND_1273 = {1{`RANDOM}};
  ram_1271 = _RAND_1273[7:0];
  _RAND_1274 = {1{`RANDOM}};
  ram_1272 = _RAND_1274[7:0];
  _RAND_1275 = {1{`RANDOM}};
  ram_1273 = _RAND_1275[7:0];
  _RAND_1276 = {1{`RANDOM}};
  ram_1274 = _RAND_1276[7:0];
  _RAND_1277 = {1{`RANDOM}};
  ram_1275 = _RAND_1277[7:0];
  _RAND_1278 = {1{`RANDOM}};
  ram_1276 = _RAND_1278[7:0];
  _RAND_1279 = {1{`RANDOM}};
  ram_1277 = _RAND_1279[7:0];
  _RAND_1280 = {1{`RANDOM}};
  ram_1278 = _RAND_1280[7:0];
  _RAND_1281 = {1{`RANDOM}};
  ram_1279 = _RAND_1281[7:0];
  _RAND_1282 = {1{`RANDOM}};
  ram_1280 = _RAND_1282[7:0];
  _RAND_1283 = {1{`RANDOM}};
  ram_1281 = _RAND_1283[7:0];
  _RAND_1284 = {1{`RANDOM}};
  ram_1282 = _RAND_1284[7:0];
  _RAND_1285 = {1{`RANDOM}};
  ram_1283 = _RAND_1285[7:0];
  _RAND_1286 = {1{`RANDOM}};
  ram_1284 = _RAND_1286[7:0];
  _RAND_1287 = {1{`RANDOM}};
  ram_1285 = _RAND_1287[7:0];
  _RAND_1288 = {1{`RANDOM}};
  ram_1286 = _RAND_1288[7:0];
  _RAND_1289 = {1{`RANDOM}};
  ram_1287 = _RAND_1289[7:0];
  _RAND_1290 = {1{`RANDOM}};
  ram_1288 = _RAND_1290[7:0];
  _RAND_1291 = {1{`RANDOM}};
  ram_1289 = _RAND_1291[7:0];
  _RAND_1292 = {1{`RANDOM}};
  ram_1290 = _RAND_1292[7:0];
  _RAND_1293 = {1{`RANDOM}};
  ram_1291 = _RAND_1293[7:0];
  _RAND_1294 = {1{`RANDOM}};
  ram_1292 = _RAND_1294[7:0];
  _RAND_1295 = {1{`RANDOM}};
  ram_1293 = _RAND_1295[7:0];
  _RAND_1296 = {1{`RANDOM}};
  ram_1294 = _RAND_1296[7:0];
  _RAND_1297 = {1{`RANDOM}};
  ram_1295 = _RAND_1297[7:0];
  _RAND_1298 = {1{`RANDOM}};
  ram_1296 = _RAND_1298[7:0];
  _RAND_1299 = {1{`RANDOM}};
  ram_1297 = _RAND_1299[7:0];
  _RAND_1300 = {1{`RANDOM}};
  ram_1298 = _RAND_1300[7:0];
  _RAND_1301 = {1{`RANDOM}};
  ram_1299 = _RAND_1301[7:0];
  _RAND_1302 = {1{`RANDOM}};
  ram_1300 = _RAND_1302[7:0];
  _RAND_1303 = {1{`RANDOM}};
  ram_1301 = _RAND_1303[7:0];
  _RAND_1304 = {1{`RANDOM}};
  ram_1302 = _RAND_1304[7:0];
  _RAND_1305 = {1{`RANDOM}};
  ram_1303 = _RAND_1305[7:0];
  _RAND_1306 = {1{`RANDOM}};
  ram_1304 = _RAND_1306[7:0];
  _RAND_1307 = {1{`RANDOM}};
  ram_1305 = _RAND_1307[7:0];
  _RAND_1308 = {1{`RANDOM}};
  ram_1306 = _RAND_1308[7:0];
  _RAND_1309 = {1{`RANDOM}};
  ram_1307 = _RAND_1309[7:0];
  _RAND_1310 = {1{`RANDOM}};
  ram_1308 = _RAND_1310[7:0];
  _RAND_1311 = {1{`RANDOM}};
  ram_1309 = _RAND_1311[7:0];
  _RAND_1312 = {1{`RANDOM}};
  ram_1310 = _RAND_1312[7:0];
  _RAND_1313 = {1{`RANDOM}};
  ram_1311 = _RAND_1313[7:0];
  _RAND_1314 = {1{`RANDOM}};
  ram_1312 = _RAND_1314[7:0];
  _RAND_1315 = {1{`RANDOM}};
  ram_1313 = _RAND_1315[7:0];
  _RAND_1316 = {1{`RANDOM}};
  ram_1314 = _RAND_1316[7:0];
  _RAND_1317 = {1{`RANDOM}};
  ram_1315 = _RAND_1317[7:0];
  _RAND_1318 = {1{`RANDOM}};
  ram_1316 = _RAND_1318[7:0];
  _RAND_1319 = {1{`RANDOM}};
  ram_1317 = _RAND_1319[7:0];
  _RAND_1320 = {1{`RANDOM}};
  ram_1318 = _RAND_1320[7:0];
  _RAND_1321 = {1{`RANDOM}};
  ram_1319 = _RAND_1321[7:0];
  _RAND_1322 = {1{`RANDOM}};
  ram_1320 = _RAND_1322[7:0];
  _RAND_1323 = {1{`RANDOM}};
  ram_1321 = _RAND_1323[7:0];
  _RAND_1324 = {1{`RANDOM}};
  ram_1322 = _RAND_1324[7:0];
  _RAND_1325 = {1{`RANDOM}};
  ram_1323 = _RAND_1325[7:0];
  _RAND_1326 = {1{`RANDOM}};
  ram_1324 = _RAND_1326[7:0];
  _RAND_1327 = {1{`RANDOM}};
  ram_1325 = _RAND_1327[7:0];
  _RAND_1328 = {1{`RANDOM}};
  ram_1326 = _RAND_1328[7:0];
  _RAND_1329 = {1{`RANDOM}};
  ram_1327 = _RAND_1329[7:0];
  _RAND_1330 = {1{`RANDOM}};
  ram_1328 = _RAND_1330[7:0];
  _RAND_1331 = {1{`RANDOM}};
  ram_1329 = _RAND_1331[7:0];
  _RAND_1332 = {1{`RANDOM}};
  ram_1330 = _RAND_1332[7:0];
  _RAND_1333 = {1{`RANDOM}};
  ram_1331 = _RAND_1333[7:0];
  _RAND_1334 = {1{`RANDOM}};
  ram_1332 = _RAND_1334[7:0];
  _RAND_1335 = {1{`RANDOM}};
  ram_1333 = _RAND_1335[7:0];
  _RAND_1336 = {1{`RANDOM}};
  ram_1334 = _RAND_1336[7:0];
  _RAND_1337 = {1{`RANDOM}};
  ram_1335 = _RAND_1337[7:0];
  _RAND_1338 = {1{`RANDOM}};
  ram_1336 = _RAND_1338[7:0];
  _RAND_1339 = {1{`RANDOM}};
  ram_1337 = _RAND_1339[7:0];
  _RAND_1340 = {1{`RANDOM}};
  ram_1338 = _RAND_1340[7:0];
  _RAND_1341 = {1{`RANDOM}};
  ram_1339 = _RAND_1341[7:0];
  _RAND_1342 = {1{`RANDOM}};
  ram_1340 = _RAND_1342[7:0];
  _RAND_1343 = {1{`RANDOM}};
  ram_1341 = _RAND_1343[7:0];
  _RAND_1344 = {1{`RANDOM}};
  ram_1342 = _RAND_1344[7:0];
  _RAND_1345 = {1{`RANDOM}};
  ram_1343 = _RAND_1345[7:0];
  _RAND_1346 = {1{`RANDOM}};
  ram_1344 = _RAND_1346[7:0];
  _RAND_1347 = {1{`RANDOM}};
  ram_1345 = _RAND_1347[7:0];
  _RAND_1348 = {1{`RANDOM}};
  ram_1346 = _RAND_1348[7:0];
  _RAND_1349 = {1{`RANDOM}};
  ram_1347 = _RAND_1349[7:0];
  _RAND_1350 = {1{`RANDOM}};
  ram_1348 = _RAND_1350[7:0];
  _RAND_1351 = {1{`RANDOM}};
  ram_1349 = _RAND_1351[7:0];
  _RAND_1352 = {1{`RANDOM}};
  ram_1350 = _RAND_1352[7:0];
  _RAND_1353 = {1{`RANDOM}};
  ram_1351 = _RAND_1353[7:0];
  _RAND_1354 = {1{`RANDOM}};
  ram_1352 = _RAND_1354[7:0];
  _RAND_1355 = {1{`RANDOM}};
  ram_1353 = _RAND_1355[7:0];
  _RAND_1356 = {1{`RANDOM}};
  ram_1354 = _RAND_1356[7:0];
  _RAND_1357 = {1{`RANDOM}};
  ram_1355 = _RAND_1357[7:0];
  _RAND_1358 = {1{`RANDOM}};
  ram_1356 = _RAND_1358[7:0];
  _RAND_1359 = {1{`RANDOM}};
  ram_1357 = _RAND_1359[7:0];
  _RAND_1360 = {1{`RANDOM}};
  ram_1358 = _RAND_1360[7:0];
  _RAND_1361 = {1{`RANDOM}};
  ram_1359 = _RAND_1361[7:0];
  _RAND_1362 = {1{`RANDOM}};
  ram_1360 = _RAND_1362[7:0];
  _RAND_1363 = {1{`RANDOM}};
  ram_1361 = _RAND_1363[7:0];
  _RAND_1364 = {1{`RANDOM}};
  ram_1362 = _RAND_1364[7:0];
  _RAND_1365 = {1{`RANDOM}};
  ram_1363 = _RAND_1365[7:0];
  _RAND_1366 = {1{`RANDOM}};
  ram_1364 = _RAND_1366[7:0];
  _RAND_1367 = {1{`RANDOM}};
  ram_1365 = _RAND_1367[7:0];
  _RAND_1368 = {1{`RANDOM}};
  ram_1366 = _RAND_1368[7:0];
  _RAND_1369 = {1{`RANDOM}};
  ram_1367 = _RAND_1369[7:0];
  _RAND_1370 = {1{`RANDOM}};
  ram_1368 = _RAND_1370[7:0];
  _RAND_1371 = {1{`RANDOM}};
  ram_1369 = _RAND_1371[7:0];
  _RAND_1372 = {1{`RANDOM}};
  ram_1370 = _RAND_1372[7:0];
  _RAND_1373 = {1{`RANDOM}};
  ram_1371 = _RAND_1373[7:0];
  _RAND_1374 = {1{`RANDOM}};
  ram_1372 = _RAND_1374[7:0];
  _RAND_1375 = {1{`RANDOM}};
  ram_1373 = _RAND_1375[7:0];
  _RAND_1376 = {1{`RANDOM}};
  ram_1374 = _RAND_1376[7:0];
  _RAND_1377 = {1{`RANDOM}};
  ram_1375 = _RAND_1377[7:0];
  _RAND_1378 = {1{`RANDOM}};
  ram_1376 = _RAND_1378[7:0];
  _RAND_1379 = {1{`RANDOM}};
  ram_1377 = _RAND_1379[7:0];
  _RAND_1380 = {1{`RANDOM}};
  ram_1378 = _RAND_1380[7:0];
  _RAND_1381 = {1{`RANDOM}};
  ram_1379 = _RAND_1381[7:0];
  _RAND_1382 = {1{`RANDOM}};
  ram_1380 = _RAND_1382[7:0];
  _RAND_1383 = {1{`RANDOM}};
  ram_1381 = _RAND_1383[7:0];
  _RAND_1384 = {1{`RANDOM}};
  ram_1382 = _RAND_1384[7:0];
  _RAND_1385 = {1{`RANDOM}};
  ram_1383 = _RAND_1385[7:0];
  _RAND_1386 = {1{`RANDOM}};
  ram_1384 = _RAND_1386[7:0];
  _RAND_1387 = {1{`RANDOM}};
  ram_1385 = _RAND_1387[7:0];
  _RAND_1388 = {1{`RANDOM}};
  ram_1386 = _RAND_1388[7:0];
  _RAND_1389 = {1{`RANDOM}};
  ram_1387 = _RAND_1389[7:0];
  _RAND_1390 = {1{`RANDOM}};
  ram_1388 = _RAND_1390[7:0];
  _RAND_1391 = {1{`RANDOM}};
  ram_1389 = _RAND_1391[7:0];
  _RAND_1392 = {1{`RANDOM}};
  ram_1390 = _RAND_1392[7:0];
  _RAND_1393 = {1{`RANDOM}};
  ram_1391 = _RAND_1393[7:0];
  _RAND_1394 = {1{`RANDOM}};
  ram_1392 = _RAND_1394[7:0];
  _RAND_1395 = {1{`RANDOM}};
  ram_1393 = _RAND_1395[7:0];
  _RAND_1396 = {1{`RANDOM}};
  ram_1394 = _RAND_1396[7:0];
  _RAND_1397 = {1{`RANDOM}};
  ram_1395 = _RAND_1397[7:0];
  _RAND_1398 = {1{`RANDOM}};
  ram_1396 = _RAND_1398[7:0];
  _RAND_1399 = {1{`RANDOM}};
  ram_1397 = _RAND_1399[7:0];
  _RAND_1400 = {1{`RANDOM}};
  ram_1398 = _RAND_1400[7:0];
  _RAND_1401 = {1{`RANDOM}};
  ram_1399 = _RAND_1401[7:0];
  _RAND_1402 = {1{`RANDOM}};
  ram_1400 = _RAND_1402[7:0];
  _RAND_1403 = {1{`RANDOM}};
  ram_1401 = _RAND_1403[7:0];
  _RAND_1404 = {1{`RANDOM}};
  ram_1402 = _RAND_1404[7:0];
  _RAND_1405 = {1{`RANDOM}};
  ram_1403 = _RAND_1405[7:0];
  _RAND_1406 = {1{`RANDOM}};
  ram_1404 = _RAND_1406[7:0];
  _RAND_1407 = {1{`RANDOM}};
  ram_1405 = _RAND_1407[7:0];
  _RAND_1408 = {1{`RANDOM}};
  ram_1406 = _RAND_1408[7:0];
  _RAND_1409 = {1{`RANDOM}};
  ram_1407 = _RAND_1409[7:0];
  _RAND_1410 = {1{`RANDOM}};
  ram_1408 = _RAND_1410[7:0];
  _RAND_1411 = {1{`RANDOM}};
  ram_1409 = _RAND_1411[7:0];
  _RAND_1412 = {1{`RANDOM}};
  ram_1410 = _RAND_1412[7:0];
  _RAND_1413 = {1{`RANDOM}};
  ram_1411 = _RAND_1413[7:0];
  _RAND_1414 = {1{`RANDOM}};
  ram_1412 = _RAND_1414[7:0];
  _RAND_1415 = {1{`RANDOM}};
  ram_1413 = _RAND_1415[7:0];
  _RAND_1416 = {1{`RANDOM}};
  ram_1414 = _RAND_1416[7:0];
  _RAND_1417 = {1{`RANDOM}};
  ram_1415 = _RAND_1417[7:0];
  _RAND_1418 = {1{`RANDOM}};
  ram_1416 = _RAND_1418[7:0];
  _RAND_1419 = {1{`RANDOM}};
  ram_1417 = _RAND_1419[7:0];
  _RAND_1420 = {1{`RANDOM}};
  ram_1418 = _RAND_1420[7:0];
  _RAND_1421 = {1{`RANDOM}};
  ram_1419 = _RAND_1421[7:0];
  _RAND_1422 = {1{`RANDOM}};
  ram_1420 = _RAND_1422[7:0];
  _RAND_1423 = {1{`RANDOM}};
  ram_1421 = _RAND_1423[7:0];
  _RAND_1424 = {1{`RANDOM}};
  ram_1422 = _RAND_1424[7:0];
  _RAND_1425 = {1{`RANDOM}};
  ram_1423 = _RAND_1425[7:0];
  _RAND_1426 = {1{`RANDOM}};
  ram_1424 = _RAND_1426[7:0];
  _RAND_1427 = {1{`RANDOM}};
  ram_1425 = _RAND_1427[7:0];
  _RAND_1428 = {1{`RANDOM}};
  ram_1426 = _RAND_1428[7:0];
  _RAND_1429 = {1{`RANDOM}};
  ram_1427 = _RAND_1429[7:0];
  _RAND_1430 = {1{`RANDOM}};
  ram_1428 = _RAND_1430[7:0];
  _RAND_1431 = {1{`RANDOM}};
  ram_1429 = _RAND_1431[7:0];
  _RAND_1432 = {1{`RANDOM}};
  ram_1430 = _RAND_1432[7:0];
  _RAND_1433 = {1{`RANDOM}};
  ram_1431 = _RAND_1433[7:0];
  _RAND_1434 = {1{`RANDOM}};
  ram_1432 = _RAND_1434[7:0];
  _RAND_1435 = {1{`RANDOM}};
  ram_1433 = _RAND_1435[7:0];
  _RAND_1436 = {1{`RANDOM}};
  ram_1434 = _RAND_1436[7:0];
  _RAND_1437 = {1{`RANDOM}};
  ram_1435 = _RAND_1437[7:0];
  _RAND_1438 = {1{`RANDOM}};
  ram_1436 = _RAND_1438[7:0];
  _RAND_1439 = {1{`RANDOM}};
  ram_1437 = _RAND_1439[7:0];
  _RAND_1440 = {1{`RANDOM}};
  ram_1438 = _RAND_1440[7:0];
  _RAND_1441 = {1{`RANDOM}};
  ram_1439 = _RAND_1441[7:0];
  _RAND_1442 = {1{`RANDOM}};
  ram_1440 = _RAND_1442[7:0];
  _RAND_1443 = {1{`RANDOM}};
  ram_1441 = _RAND_1443[7:0];
  _RAND_1444 = {1{`RANDOM}};
  ram_1442 = _RAND_1444[7:0];
  _RAND_1445 = {1{`RANDOM}};
  ram_1443 = _RAND_1445[7:0];
  _RAND_1446 = {1{`RANDOM}};
  ram_1444 = _RAND_1446[7:0];
  _RAND_1447 = {1{`RANDOM}};
  ram_1445 = _RAND_1447[7:0];
  _RAND_1448 = {1{`RANDOM}};
  ram_1446 = _RAND_1448[7:0];
  _RAND_1449 = {1{`RANDOM}};
  ram_1447 = _RAND_1449[7:0];
  _RAND_1450 = {1{`RANDOM}};
  ram_1448 = _RAND_1450[7:0];
  _RAND_1451 = {1{`RANDOM}};
  ram_1449 = _RAND_1451[7:0];
  _RAND_1452 = {1{`RANDOM}};
  ram_1450 = _RAND_1452[7:0];
  _RAND_1453 = {1{`RANDOM}};
  ram_1451 = _RAND_1453[7:0];
  _RAND_1454 = {1{`RANDOM}};
  ram_1452 = _RAND_1454[7:0];
  _RAND_1455 = {1{`RANDOM}};
  ram_1453 = _RAND_1455[7:0];
  _RAND_1456 = {1{`RANDOM}};
  ram_1454 = _RAND_1456[7:0];
  _RAND_1457 = {1{`RANDOM}};
  ram_1455 = _RAND_1457[7:0];
  _RAND_1458 = {1{`RANDOM}};
  ram_1456 = _RAND_1458[7:0];
  _RAND_1459 = {1{`RANDOM}};
  ram_1457 = _RAND_1459[7:0];
  _RAND_1460 = {1{`RANDOM}};
  ram_1458 = _RAND_1460[7:0];
  _RAND_1461 = {1{`RANDOM}};
  ram_1459 = _RAND_1461[7:0];
  _RAND_1462 = {1{`RANDOM}};
  ram_1460 = _RAND_1462[7:0];
  _RAND_1463 = {1{`RANDOM}};
  ram_1461 = _RAND_1463[7:0];
  _RAND_1464 = {1{`RANDOM}};
  ram_1462 = _RAND_1464[7:0];
  _RAND_1465 = {1{`RANDOM}};
  ram_1463 = _RAND_1465[7:0];
  _RAND_1466 = {1{`RANDOM}};
  ram_1464 = _RAND_1466[7:0];
  _RAND_1467 = {1{`RANDOM}};
  ram_1465 = _RAND_1467[7:0];
  _RAND_1468 = {1{`RANDOM}};
  ram_1466 = _RAND_1468[7:0];
  _RAND_1469 = {1{`RANDOM}};
  ram_1467 = _RAND_1469[7:0];
  _RAND_1470 = {1{`RANDOM}};
  ram_1468 = _RAND_1470[7:0];
  _RAND_1471 = {1{`RANDOM}};
  ram_1469 = _RAND_1471[7:0];
  _RAND_1472 = {1{`RANDOM}};
  ram_1470 = _RAND_1472[7:0];
  _RAND_1473 = {1{`RANDOM}};
  ram_1471 = _RAND_1473[7:0];
  _RAND_1474 = {1{`RANDOM}};
  ram_1472 = _RAND_1474[7:0];
  _RAND_1475 = {1{`RANDOM}};
  ram_1473 = _RAND_1475[7:0];
  _RAND_1476 = {1{`RANDOM}};
  ram_1474 = _RAND_1476[7:0];
  _RAND_1477 = {1{`RANDOM}};
  ram_1475 = _RAND_1477[7:0];
  _RAND_1478 = {1{`RANDOM}};
  ram_1476 = _RAND_1478[7:0];
  _RAND_1479 = {1{`RANDOM}};
  ram_1477 = _RAND_1479[7:0];
  _RAND_1480 = {1{`RANDOM}};
  ram_1478 = _RAND_1480[7:0];
  _RAND_1481 = {1{`RANDOM}};
  ram_1479 = _RAND_1481[7:0];
  _RAND_1482 = {1{`RANDOM}};
  ram_1480 = _RAND_1482[7:0];
  _RAND_1483 = {1{`RANDOM}};
  ram_1481 = _RAND_1483[7:0];
  _RAND_1484 = {1{`RANDOM}};
  ram_1482 = _RAND_1484[7:0];
  _RAND_1485 = {1{`RANDOM}};
  ram_1483 = _RAND_1485[7:0];
  _RAND_1486 = {1{`RANDOM}};
  ram_1484 = _RAND_1486[7:0];
  _RAND_1487 = {1{`RANDOM}};
  ram_1485 = _RAND_1487[7:0];
  _RAND_1488 = {1{`RANDOM}};
  ram_1486 = _RAND_1488[7:0];
  _RAND_1489 = {1{`RANDOM}};
  ram_1487 = _RAND_1489[7:0];
  _RAND_1490 = {1{`RANDOM}};
  ram_1488 = _RAND_1490[7:0];
  _RAND_1491 = {1{`RANDOM}};
  ram_1489 = _RAND_1491[7:0];
  _RAND_1492 = {1{`RANDOM}};
  ram_1490 = _RAND_1492[7:0];
  _RAND_1493 = {1{`RANDOM}};
  ram_1491 = _RAND_1493[7:0];
  _RAND_1494 = {1{`RANDOM}};
  ram_1492 = _RAND_1494[7:0];
  _RAND_1495 = {1{`RANDOM}};
  ram_1493 = _RAND_1495[7:0];
  _RAND_1496 = {1{`RANDOM}};
  ram_1494 = _RAND_1496[7:0];
  _RAND_1497 = {1{`RANDOM}};
  ram_1495 = _RAND_1497[7:0];
  _RAND_1498 = {1{`RANDOM}};
  ram_1496 = _RAND_1498[7:0];
  _RAND_1499 = {1{`RANDOM}};
  ram_1497 = _RAND_1499[7:0];
  _RAND_1500 = {1{`RANDOM}};
  ram_1498 = _RAND_1500[7:0];
  _RAND_1501 = {1{`RANDOM}};
  ram_1499 = _RAND_1501[7:0];
  _RAND_1502 = {1{`RANDOM}};
  ram_1500 = _RAND_1502[7:0];
  _RAND_1503 = {1{`RANDOM}};
  ram_1501 = _RAND_1503[7:0];
  _RAND_1504 = {1{`RANDOM}};
  ram_1502 = _RAND_1504[7:0];
  _RAND_1505 = {1{`RANDOM}};
  ram_1503 = _RAND_1505[7:0];
  _RAND_1506 = {1{`RANDOM}};
  ram_1504 = _RAND_1506[7:0];
  _RAND_1507 = {1{`RANDOM}};
  ram_1505 = _RAND_1507[7:0];
  _RAND_1508 = {1{`RANDOM}};
  ram_1506 = _RAND_1508[7:0];
  _RAND_1509 = {1{`RANDOM}};
  ram_1507 = _RAND_1509[7:0];
  _RAND_1510 = {1{`RANDOM}};
  ram_1508 = _RAND_1510[7:0];
  _RAND_1511 = {1{`RANDOM}};
  ram_1509 = _RAND_1511[7:0];
  _RAND_1512 = {1{`RANDOM}};
  ram_1510 = _RAND_1512[7:0];
  _RAND_1513 = {1{`RANDOM}};
  ram_1511 = _RAND_1513[7:0];
  _RAND_1514 = {1{`RANDOM}};
  ram_1512 = _RAND_1514[7:0];
  _RAND_1515 = {1{`RANDOM}};
  ram_1513 = _RAND_1515[7:0];
  _RAND_1516 = {1{`RANDOM}};
  ram_1514 = _RAND_1516[7:0];
  _RAND_1517 = {1{`RANDOM}};
  ram_1515 = _RAND_1517[7:0];
  _RAND_1518 = {1{`RANDOM}};
  ram_1516 = _RAND_1518[7:0];
  _RAND_1519 = {1{`RANDOM}};
  ram_1517 = _RAND_1519[7:0];
  _RAND_1520 = {1{`RANDOM}};
  ram_1518 = _RAND_1520[7:0];
  _RAND_1521 = {1{`RANDOM}};
  ram_1519 = _RAND_1521[7:0];
  _RAND_1522 = {1{`RANDOM}};
  ram_1520 = _RAND_1522[7:0];
  _RAND_1523 = {1{`RANDOM}};
  ram_1521 = _RAND_1523[7:0];
  _RAND_1524 = {1{`RANDOM}};
  ram_1522 = _RAND_1524[7:0];
  _RAND_1525 = {1{`RANDOM}};
  ram_1523 = _RAND_1525[7:0];
  _RAND_1526 = {1{`RANDOM}};
  ram_1524 = _RAND_1526[7:0];
  _RAND_1527 = {1{`RANDOM}};
  ram_1525 = _RAND_1527[7:0];
  _RAND_1528 = {1{`RANDOM}};
  ram_1526 = _RAND_1528[7:0];
  _RAND_1529 = {1{`RANDOM}};
  ram_1527 = _RAND_1529[7:0];
  _RAND_1530 = {1{`RANDOM}};
  ram_1528 = _RAND_1530[7:0];
  _RAND_1531 = {1{`RANDOM}};
  ram_1529 = _RAND_1531[7:0];
  _RAND_1532 = {1{`RANDOM}};
  ram_1530 = _RAND_1532[7:0];
  _RAND_1533 = {1{`RANDOM}};
  ram_1531 = _RAND_1533[7:0];
  _RAND_1534 = {1{`RANDOM}};
  ram_1532 = _RAND_1534[7:0];
  _RAND_1535 = {1{`RANDOM}};
  ram_1533 = _RAND_1535[7:0];
  _RAND_1536 = {1{`RANDOM}};
  ram_1534 = _RAND_1536[7:0];
  _RAND_1537 = {1{`RANDOM}};
  ram_1535 = _RAND_1537[7:0];
  _RAND_1538 = {1{`RANDOM}};
  ram_1536 = _RAND_1538[7:0];
  _RAND_1539 = {1{`RANDOM}};
  ram_1537 = _RAND_1539[7:0];
  _RAND_1540 = {1{`RANDOM}};
  ram_1538 = _RAND_1540[7:0];
  _RAND_1541 = {1{`RANDOM}};
  ram_1539 = _RAND_1541[7:0];
  _RAND_1542 = {1{`RANDOM}};
  ram_1540 = _RAND_1542[7:0];
  _RAND_1543 = {1{`RANDOM}};
  ram_1541 = _RAND_1543[7:0];
  _RAND_1544 = {1{`RANDOM}};
  ram_1542 = _RAND_1544[7:0];
  _RAND_1545 = {1{`RANDOM}};
  ram_1543 = _RAND_1545[7:0];
  _RAND_1546 = {1{`RANDOM}};
  ram_1544 = _RAND_1546[7:0];
  _RAND_1547 = {1{`RANDOM}};
  ram_1545 = _RAND_1547[7:0];
  _RAND_1548 = {1{`RANDOM}};
  ram_1546 = _RAND_1548[7:0];
  _RAND_1549 = {1{`RANDOM}};
  ram_1547 = _RAND_1549[7:0];
  _RAND_1550 = {1{`RANDOM}};
  ram_1548 = _RAND_1550[7:0];
  _RAND_1551 = {1{`RANDOM}};
  ram_1549 = _RAND_1551[7:0];
  _RAND_1552 = {1{`RANDOM}};
  ram_1550 = _RAND_1552[7:0];
  _RAND_1553 = {1{`RANDOM}};
  ram_1551 = _RAND_1553[7:0];
  _RAND_1554 = {1{`RANDOM}};
  ram_1552 = _RAND_1554[7:0];
  _RAND_1555 = {1{`RANDOM}};
  ram_1553 = _RAND_1555[7:0];
  _RAND_1556 = {1{`RANDOM}};
  ram_1554 = _RAND_1556[7:0];
  _RAND_1557 = {1{`RANDOM}};
  ram_1555 = _RAND_1557[7:0];
  _RAND_1558 = {1{`RANDOM}};
  ram_1556 = _RAND_1558[7:0];
  _RAND_1559 = {1{`RANDOM}};
  ram_1557 = _RAND_1559[7:0];
  _RAND_1560 = {1{`RANDOM}};
  ram_1558 = _RAND_1560[7:0];
  _RAND_1561 = {1{`RANDOM}};
  ram_1559 = _RAND_1561[7:0];
  _RAND_1562 = {1{`RANDOM}};
  ram_1560 = _RAND_1562[7:0];
  _RAND_1563 = {1{`RANDOM}};
  ram_1561 = _RAND_1563[7:0];
  _RAND_1564 = {1{`RANDOM}};
  ram_1562 = _RAND_1564[7:0];
  _RAND_1565 = {1{`RANDOM}};
  ram_1563 = _RAND_1565[7:0];
  _RAND_1566 = {1{`RANDOM}};
  ram_1564 = _RAND_1566[7:0];
  _RAND_1567 = {1{`RANDOM}};
  ram_1565 = _RAND_1567[7:0];
  _RAND_1568 = {1{`RANDOM}};
  ram_1566 = _RAND_1568[7:0];
  _RAND_1569 = {1{`RANDOM}};
  ram_1567 = _RAND_1569[7:0];
  _RAND_1570 = {1{`RANDOM}};
  ram_1568 = _RAND_1570[7:0];
  _RAND_1571 = {1{`RANDOM}};
  ram_1569 = _RAND_1571[7:0];
  _RAND_1572 = {1{`RANDOM}};
  ram_1570 = _RAND_1572[7:0];
  _RAND_1573 = {1{`RANDOM}};
  ram_1571 = _RAND_1573[7:0];
  _RAND_1574 = {1{`RANDOM}};
  ram_1572 = _RAND_1574[7:0];
  _RAND_1575 = {1{`RANDOM}};
  ram_1573 = _RAND_1575[7:0];
  _RAND_1576 = {1{`RANDOM}};
  ram_1574 = _RAND_1576[7:0];
  _RAND_1577 = {1{`RANDOM}};
  ram_1575 = _RAND_1577[7:0];
  _RAND_1578 = {1{`RANDOM}};
  ram_1576 = _RAND_1578[7:0];
  _RAND_1579 = {1{`RANDOM}};
  ram_1577 = _RAND_1579[7:0];
  _RAND_1580 = {1{`RANDOM}};
  ram_1578 = _RAND_1580[7:0];
  _RAND_1581 = {1{`RANDOM}};
  ram_1579 = _RAND_1581[7:0];
  _RAND_1582 = {1{`RANDOM}};
  ram_1580 = _RAND_1582[7:0];
  _RAND_1583 = {1{`RANDOM}};
  ram_1581 = _RAND_1583[7:0];
  _RAND_1584 = {1{`RANDOM}};
  ram_1582 = _RAND_1584[7:0];
  _RAND_1585 = {1{`RANDOM}};
  ram_1583 = _RAND_1585[7:0];
  _RAND_1586 = {1{`RANDOM}};
  ram_1584 = _RAND_1586[7:0];
  _RAND_1587 = {1{`RANDOM}};
  ram_1585 = _RAND_1587[7:0];
  _RAND_1588 = {1{`RANDOM}};
  ram_1586 = _RAND_1588[7:0];
  _RAND_1589 = {1{`RANDOM}};
  ram_1587 = _RAND_1589[7:0];
  _RAND_1590 = {1{`RANDOM}};
  ram_1588 = _RAND_1590[7:0];
  _RAND_1591 = {1{`RANDOM}};
  ram_1589 = _RAND_1591[7:0];
  _RAND_1592 = {1{`RANDOM}};
  ram_1590 = _RAND_1592[7:0];
  _RAND_1593 = {1{`RANDOM}};
  ram_1591 = _RAND_1593[7:0];
  _RAND_1594 = {1{`RANDOM}};
  ram_1592 = _RAND_1594[7:0];
  _RAND_1595 = {1{`RANDOM}};
  ram_1593 = _RAND_1595[7:0];
  _RAND_1596 = {1{`RANDOM}};
  ram_1594 = _RAND_1596[7:0];
  _RAND_1597 = {1{`RANDOM}};
  ram_1595 = _RAND_1597[7:0];
  _RAND_1598 = {1{`RANDOM}};
  ram_1596 = _RAND_1598[7:0];
  _RAND_1599 = {1{`RANDOM}};
  ram_1597 = _RAND_1599[7:0];
  _RAND_1600 = {1{`RANDOM}};
  ram_1598 = _RAND_1600[7:0];
  _RAND_1601 = {1{`RANDOM}};
  ram_1599 = _RAND_1601[7:0];
  _RAND_1602 = {1{`RANDOM}};
  ram_1600 = _RAND_1602[7:0];
  _RAND_1603 = {1{`RANDOM}};
  ram_1601 = _RAND_1603[7:0];
  _RAND_1604 = {1{`RANDOM}};
  ram_1602 = _RAND_1604[7:0];
  _RAND_1605 = {1{`RANDOM}};
  ram_1603 = _RAND_1605[7:0];
  _RAND_1606 = {1{`RANDOM}};
  ram_1604 = _RAND_1606[7:0];
  _RAND_1607 = {1{`RANDOM}};
  ram_1605 = _RAND_1607[7:0];
  _RAND_1608 = {1{`RANDOM}};
  ram_1606 = _RAND_1608[7:0];
  _RAND_1609 = {1{`RANDOM}};
  ram_1607 = _RAND_1609[7:0];
  _RAND_1610 = {1{`RANDOM}};
  ram_1608 = _RAND_1610[7:0];
  _RAND_1611 = {1{`RANDOM}};
  ram_1609 = _RAND_1611[7:0];
  _RAND_1612 = {1{`RANDOM}};
  ram_1610 = _RAND_1612[7:0];
  _RAND_1613 = {1{`RANDOM}};
  ram_1611 = _RAND_1613[7:0];
  _RAND_1614 = {1{`RANDOM}};
  ram_1612 = _RAND_1614[7:0];
  _RAND_1615 = {1{`RANDOM}};
  ram_1613 = _RAND_1615[7:0];
  _RAND_1616 = {1{`RANDOM}};
  ram_1614 = _RAND_1616[7:0];
  _RAND_1617 = {1{`RANDOM}};
  ram_1615 = _RAND_1617[7:0];
  _RAND_1618 = {1{`RANDOM}};
  ram_1616 = _RAND_1618[7:0];
  _RAND_1619 = {1{`RANDOM}};
  ram_1617 = _RAND_1619[7:0];
  _RAND_1620 = {1{`RANDOM}};
  ram_1618 = _RAND_1620[7:0];
  _RAND_1621 = {1{`RANDOM}};
  ram_1619 = _RAND_1621[7:0];
  _RAND_1622 = {1{`RANDOM}};
  ram_1620 = _RAND_1622[7:0];
  _RAND_1623 = {1{`RANDOM}};
  ram_1621 = _RAND_1623[7:0];
  _RAND_1624 = {1{`RANDOM}};
  ram_1622 = _RAND_1624[7:0];
  _RAND_1625 = {1{`RANDOM}};
  ram_1623 = _RAND_1625[7:0];
  _RAND_1626 = {1{`RANDOM}};
  ram_1624 = _RAND_1626[7:0];
  _RAND_1627 = {1{`RANDOM}};
  ram_1625 = _RAND_1627[7:0];
  _RAND_1628 = {1{`RANDOM}};
  ram_1626 = _RAND_1628[7:0];
  _RAND_1629 = {1{`RANDOM}};
  ram_1627 = _RAND_1629[7:0];
  _RAND_1630 = {1{`RANDOM}};
  ram_1628 = _RAND_1630[7:0];
  _RAND_1631 = {1{`RANDOM}};
  ram_1629 = _RAND_1631[7:0];
  _RAND_1632 = {1{`RANDOM}};
  ram_1630 = _RAND_1632[7:0];
  _RAND_1633 = {1{`RANDOM}};
  ram_1631 = _RAND_1633[7:0];
  _RAND_1634 = {1{`RANDOM}};
  ram_1632 = _RAND_1634[7:0];
  _RAND_1635 = {1{`RANDOM}};
  ram_1633 = _RAND_1635[7:0];
  _RAND_1636 = {1{`RANDOM}};
  ram_1634 = _RAND_1636[7:0];
  _RAND_1637 = {1{`RANDOM}};
  ram_1635 = _RAND_1637[7:0];
  _RAND_1638 = {1{`RANDOM}};
  ram_1636 = _RAND_1638[7:0];
  _RAND_1639 = {1{`RANDOM}};
  ram_1637 = _RAND_1639[7:0];
  _RAND_1640 = {1{`RANDOM}};
  ram_1638 = _RAND_1640[7:0];
  _RAND_1641 = {1{`RANDOM}};
  ram_1639 = _RAND_1641[7:0];
  _RAND_1642 = {1{`RANDOM}};
  ram_1640 = _RAND_1642[7:0];
  _RAND_1643 = {1{`RANDOM}};
  ram_1641 = _RAND_1643[7:0];
  _RAND_1644 = {1{`RANDOM}};
  ram_1642 = _RAND_1644[7:0];
  _RAND_1645 = {1{`RANDOM}};
  ram_1643 = _RAND_1645[7:0];
  _RAND_1646 = {1{`RANDOM}};
  ram_1644 = _RAND_1646[7:0];
  _RAND_1647 = {1{`RANDOM}};
  ram_1645 = _RAND_1647[7:0];
  _RAND_1648 = {1{`RANDOM}};
  ram_1646 = _RAND_1648[7:0];
  _RAND_1649 = {1{`RANDOM}};
  ram_1647 = _RAND_1649[7:0];
  _RAND_1650 = {1{`RANDOM}};
  ram_1648 = _RAND_1650[7:0];
  _RAND_1651 = {1{`RANDOM}};
  ram_1649 = _RAND_1651[7:0];
  _RAND_1652 = {1{`RANDOM}};
  ram_1650 = _RAND_1652[7:0];
  _RAND_1653 = {1{`RANDOM}};
  ram_1651 = _RAND_1653[7:0];
  _RAND_1654 = {1{`RANDOM}};
  ram_1652 = _RAND_1654[7:0];
  _RAND_1655 = {1{`RANDOM}};
  ram_1653 = _RAND_1655[7:0];
  _RAND_1656 = {1{`RANDOM}};
  ram_1654 = _RAND_1656[7:0];
  _RAND_1657 = {1{`RANDOM}};
  ram_1655 = _RAND_1657[7:0];
  _RAND_1658 = {1{`RANDOM}};
  ram_1656 = _RAND_1658[7:0];
  _RAND_1659 = {1{`RANDOM}};
  ram_1657 = _RAND_1659[7:0];
  _RAND_1660 = {1{`RANDOM}};
  ram_1658 = _RAND_1660[7:0];
  _RAND_1661 = {1{`RANDOM}};
  ram_1659 = _RAND_1661[7:0];
  _RAND_1662 = {1{`RANDOM}};
  ram_1660 = _RAND_1662[7:0];
  _RAND_1663 = {1{`RANDOM}};
  ram_1661 = _RAND_1663[7:0];
  _RAND_1664 = {1{`RANDOM}};
  ram_1662 = _RAND_1664[7:0];
  _RAND_1665 = {1{`RANDOM}};
  ram_1663 = _RAND_1665[7:0];
  _RAND_1666 = {1{`RANDOM}};
  ram_1664 = _RAND_1666[7:0];
  _RAND_1667 = {1{`RANDOM}};
  ram_1665 = _RAND_1667[7:0];
  _RAND_1668 = {1{`RANDOM}};
  ram_1666 = _RAND_1668[7:0];
  _RAND_1669 = {1{`RANDOM}};
  ram_1667 = _RAND_1669[7:0];
  _RAND_1670 = {1{`RANDOM}};
  ram_1668 = _RAND_1670[7:0];
  _RAND_1671 = {1{`RANDOM}};
  ram_1669 = _RAND_1671[7:0];
  _RAND_1672 = {1{`RANDOM}};
  ram_1670 = _RAND_1672[7:0];
  _RAND_1673 = {1{`RANDOM}};
  ram_1671 = _RAND_1673[7:0];
  _RAND_1674 = {1{`RANDOM}};
  ram_1672 = _RAND_1674[7:0];
  _RAND_1675 = {1{`RANDOM}};
  ram_1673 = _RAND_1675[7:0];
  _RAND_1676 = {1{`RANDOM}};
  ram_1674 = _RAND_1676[7:0];
  _RAND_1677 = {1{`RANDOM}};
  ram_1675 = _RAND_1677[7:0];
  _RAND_1678 = {1{`RANDOM}};
  ram_1676 = _RAND_1678[7:0];
  _RAND_1679 = {1{`RANDOM}};
  ram_1677 = _RAND_1679[7:0];
  _RAND_1680 = {1{`RANDOM}};
  ram_1678 = _RAND_1680[7:0];
  _RAND_1681 = {1{`RANDOM}};
  ram_1679 = _RAND_1681[7:0];
  _RAND_1682 = {1{`RANDOM}};
  ram_1680 = _RAND_1682[7:0];
  _RAND_1683 = {1{`RANDOM}};
  ram_1681 = _RAND_1683[7:0];
  _RAND_1684 = {1{`RANDOM}};
  ram_1682 = _RAND_1684[7:0];
  _RAND_1685 = {1{`RANDOM}};
  ram_1683 = _RAND_1685[7:0];
  _RAND_1686 = {1{`RANDOM}};
  ram_1684 = _RAND_1686[7:0];
  _RAND_1687 = {1{`RANDOM}};
  ram_1685 = _RAND_1687[7:0];
  _RAND_1688 = {1{`RANDOM}};
  ram_1686 = _RAND_1688[7:0];
  _RAND_1689 = {1{`RANDOM}};
  ram_1687 = _RAND_1689[7:0];
  _RAND_1690 = {1{`RANDOM}};
  ram_1688 = _RAND_1690[7:0];
  _RAND_1691 = {1{`RANDOM}};
  ram_1689 = _RAND_1691[7:0];
  _RAND_1692 = {1{`RANDOM}};
  ram_1690 = _RAND_1692[7:0];
  _RAND_1693 = {1{`RANDOM}};
  ram_1691 = _RAND_1693[7:0];
  _RAND_1694 = {1{`RANDOM}};
  ram_1692 = _RAND_1694[7:0];
  _RAND_1695 = {1{`RANDOM}};
  ram_1693 = _RAND_1695[7:0];
  _RAND_1696 = {1{`RANDOM}};
  ram_1694 = _RAND_1696[7:0];
  _RAND_1697 = {1{`RANDOM}};
  ram_1695 = _RAND_1697[7:0];
  _RAND_1698 = {1{`RANDOM}};
  ram_1696 = _RAND_1698[7:0];
  _RAND_1699 = {1{`RANDOM}};
  ram_1697 = _RAND_1699[7:0];
  _RAND_1700 = {1{`RANDOM}};
  ram_1698 = _RAND_1700[7:0];
  _RAND_1701 = {1{`RANDOM}};
  ram_1699 = _RAND_1701[7:0];
  _RAND_1702 = {1{`RANDOM}};
  ram_1700 = _RAND_1702[7:0];
  _RAND_1703 = {1{`RANDOM}};
  ram_1701 = _RAND_1703[7:0];
  _RAND_1704 = {1{`RANDOM}};
  ram_1702 = _RAND_1704[7:0];
  _RAND_1705 = {1{`RANDOM}};
  ram_1703 = _RAND_1705[7:0];
  _RAND_1706 = {1{`RANDOM}};
  ram_1704 = _RAND_1706[7:0];
  _RAND_1707 = {1{`RANDOM}};
  ram_1705 = _RAND_1707[7:0];
  _RAND_1708 = {1{`RANDOM}};
  ram_1706 = _RAND_1708[7:0];
  _RAND_1709 = {1{`RANDOM}};
  ram_1707 = _RAND_1709[7:0];
  _RAND_1710 = {1{`RANDOM}};
  ram_1708 = _RAND_1710[7:0];
  _RAND_1711 = {1{`RANDOM}};
  ram_1709 = _RAND_1711[7:0];
  _RAND_1712 = {1{`RANDOM}};
  ram_1710 = _RAND_1712[7:0];
  _RAND_1713 = {1{`RANDOM}};
  ram_1711 = _RAND_1713[7:0];
  _RAND_1714 = {1{`RANDOM}};
  ram_1712 = _RAND_1714[7:0];
  _RAND_1715 = {1{`RANDOM}};
  ram_1713 = _RAND_1715[7:0];
  _RAND_1716 = {1{`RANDOM}};
  ram_1714 = _RAND_1716[7:0];
  _RAND_1717 = {1{`RANDOM}};
  ram_1715 = _RAND_1717[7:0];
  _RAND_1718 = {1{`RANDOM}};
  ram_1716 = _RAND_1718[7:0];
  _RAND_1719 = {1{`RANDOM}};
  ram_1717 = _RAND_1719[7:0];
  _RAND_1720 = {1{`RANDOM}};
  ram_1718 = _RAND_1720[7:0];
  _RAND_1721 = {1{`RANDOM}};
  ram_1719 = _RAND_1721[7:0];
  _RAND_1722 = {1{`RANDOM}};
  ram_1720 = _RAND_1722[7:0];
  _RAND_1723 = {1{`RANDOM}};
  ram_1721 = _RAND_1723[7:0];
  _RAND_1724 = {1{`RANDOM}};
  ram_1722 = _RAND_1724[7:0];
  _RAND_1725 = {1{`RANDOM}};
  ram_1723 = _RAND_1725[7:0];
  _RAND_1726 = {1{`RANDOM}};
  ram_1724 = _RAND_1726[7:0];
  _RAND_1727 = {1{`RANDOM}};
  ram_1725 = _RAND_1727[7:0];
  _RAND_1728 = {1{`RANDOM}};
  ram_1726 = _RAND_1728[7:0];
  _RAND_1729 = {1{`RANDOM}};
  ram_1727 = _RAND_1729[7:0];
  _RAND_1730 = {1{`RANDOM}};
  ram_1728 = _RAND_1730[7:0];
  _RAND_1731 = {1{`RANDOM}};
  ram_1729 = _RAND_1731[7:0];
  _RAND_1732 = {1{`RANDOM}};
  ram_1730 = _RAND_1732[7:0];
  _RAND_1733 = {1{`RANDOM}};
  ram_1731 = _RAND_1733[7:0];
  _RAND_1734 = {1{`RANDOM}};
  ram_1732 = _RAND_1734[7:0];
  _RAND_1735 = {1{`RANDOM}};
  ram_1733 = _RAND_1735[7:0];
  _RAND_1736 = {1{`RANDOM}};
  ram_1734 = _RAND_1736[7:0];
  _RAND_1737 = {1{`RANDOM}};
  ram_1735 = _RAND_1737[7:0];
  _RAND_1738 = {1{`RANDOM}};
  ram_1736 = _RAND_1738[7:0];
  _RAND_1739 = {1{`RANDOM}};
  ram_1737 = _RAND_1739[7:0];
  _RAND_1740 = {1{`RANDOM}};
  ram_1738 = _RAND_1740[7:0];
  _RAND_1741 = {1{`RANDOM}};
  ram_1739 = _RAND_1741[7:0];
  _RAND_1742 = {1{`RANDOM}};
  ram_1740 = _RAND_1742[7:0];
  _RAND_1743 = {1{`RANDOM}};
  ram_1741 = _RAND_1743[7:0];
  _RAND_1744 = {1{`RANDOM}};
  ram_1742 = _RAND_1744[7:0];
  _RAND_1745 = {1{`RANDOM}};
  ram_1743 = _RAND_1745[7:0];
  _RAND_1746 = {1{`RANDOM}};
  ram_1744 = _RAND_1746[7:0];
  _RAND_1747 = {1{`RANDOM}};
  ram_1745 = _RAND_1747[7:0];
  _RAND_1748 = {1{`RANDOM}};
  ram_1746 = _RAND_1748[7:0];
  _RAND_1749 = {1{`RANDOM}};
  ram_1747 = _RAND_1749[7:0];
  _RAND_1750 = {1{`RANDOM}};
  ram_1748 = _RAND_1750[7:0];
  _RAND_1751 = {1{`RANDOM}};
  ram_1749 = _RAND_1751[7:0];
  _RAND_1752 = {1{`RANDOM}};
  ram_1750 = _RAND_1752[7:0];
  _RAND_1753 = {1{`RANDOM}};
  ram_1751 = _RAND_1753[7:0];
  _RAND_1754 = {1{`RANDOM}};
  ram_1752 = _RAND_1754[7:0];
  _RAND_1755 = {1{`RANDOM}};
  ram_1753 = _RAND_1755[7:0];
  _RAND_1756 = {1{`RANDOM}};
  ram_1754 = _RAND_1756[7:0];
  _RAND_1757 = {1{`RANDOM}};
  ram_1755 = _RAND_1757[7:0];
  _RAND_1758 = {1{`RANDOM}};
  ram_1756 = _RAND_1758[7:0];
  _RAND_1759 = {1{`RANDOM}};
  ram_1757 = _RAND_1759[7:0];
  _RAND_1760 = {1{`RANDOM}};
  ram_1758 = _RAND_1760[7:0];
  _RAND_1761 = {1{`RANDOM}};
  ram_1759 = _RAND_1761[7:0];
  _RAND_1762 = {1{`RANDOM}};
  ram_1760 = _RAND_1762[7:0];
  _RAND_1763 = {1{`RANDOM}};
  ram_1761 = _RAND_1763[7:0];
  _RAND_1764 = {1{`RANDOM}};
  ram_1762 = _RAND_1764[7:0];
  _RAND_1765 = {1{`RANDOM}};
  ram_1763 = _RAND_1765[7:0];
  _RAND_1766 = {1{`RANDOM}};
  ram_1764 = _RAND_1766[7:0];
  _RAND_1767 = {1{`RANDOM}};
  ram_1765 = _RAND_1767[7:0];
  _RAND_1768 = {1{`RANDOM}};
  ram_1766 = _RAND_1768[7:0];
  _RAND_1769 = {1{`RANDOM}};
  ram_1767 = _RAND_1769[7:0];
  _RAND_1770 = {1{`RANDOM}};
  ram_1768 = _RAND_1770[7:0];
  _RAND_1771 = {1{`RANDOM}};
  ram_1769 = _RAND_1771[7:0];
  _RAND_1772 = {1{`RANDOM}};
  ram_1770 = _RAND_1772[7:0];
  _RAND_1773 = {1{`RANDOM}};
  ram_1771 = _RAND_1773[7:0];
  _RAND_1774 = {1{`RANDOM}};
  ram_1772 = _RAND_1774[7:0];
  _RAND_1775 = {1{`RANDOM}};
  ram_1773 = _RAND_1775[7:0];
  _RAND_1776 = {1{`RANDOM}};
  ram_1774 = _RAND_1776[7:0];
  _RAND_1777 = {1{`RANDOM}};
  ram_1775 = _RAND_1777[7:0];
  _RAND_1778 = {1{`RANDOM}};
  ram_1776 = _RAND_1778[7:0];
  _RAND_1779 = {1{`RANDOM}};
  ram_1777 = _RAND_1779[7:0];
  _RAND_1780 = {1{`RANDOM}};
  ram_1778 = _RAND_1780[7:0];
  _RAND_1781 = {1{`RANDOM}};
  ram_1779 = _RAND_1781[7:0];
  _RAND_1782 = {1{`RANDOM}};
  ram_1780 = _RAND_1782[7:0];
  _RAND_1783 = {1{`RANDOM}};
  ram_1781 = _RAND_1783[7:0];
  _RAND_1784 = {1{`RANDOM}};
  ram_1782 = _RAND_1784[7:0];
  _RAND_1785 = {1{`RANDOM}};
  ram_1783 = _RAND_1785[7:0];
  _RAND_1786 = {1{`RANDOM}};
  ram_1784 = _RAND_1786[7:0];
  _RAND_1787 = {1{`RANDOM}};
  ram_1785 = _RAND_1787[7:0];
  _RAND_1788 = {1{`RANDOM}};
  ram_1786 = _RAND_1788[7:0];
  _RAND_1789 = {1{`RANDOM}};
  ram_1787 = _RAND_1789[7:0];
  _RAND_1790 = {1{`RANDOM}};
  ram_1788 = _RAND_1790[7:0];
  _RAND_1791 = {1{`RANDOM}};
  ram_1789 = _RAND_1791[7:0];
  _RAND_1792 = {1{`RANDOM}};
  ram_1790 = _RAND_1792[7:0];
  _RAND_1793 = {1{`RANDOM}};
  ram_1791 = _RAND_1793[7:0];
  _RAND_1794 = {1{`RANDOM}};
  ram_1792 = _RAND_1794[7:0];
  _RAND_1795 = {1{`RANDOM}};
  ram_1793 = _RAND_1795[7:0];
  _RAND_1796 = {1{`RANDOM}};
  ram_1794 = _RAND_1796[7:0];
  _RAND_1797 = {1{`RANDOM}};
  ram_1795 = _RAND_1797[7:0];
  _RAND_1798 = {1{`RANDOM}};
  ram_1796 = _RAND_1798[7:0];
  _RAND_1799 = {1{`RANDOM}};
  ram_1797 = _RAND_1799[7:0];
  _RAND_1800 = {1{`RANDOM}};
  ram_1798 = _RAND_1800[7:0];
  _RAND_1801 = {1{`RANDOM}};
  ram_1799 = _RAND_1801[7:0];
  _RAND_1802 = {1{`RANDOM}};
  ram_1800 = _RAND_1802[7:0];
  _RAND_1803 = {1{`RANDOM}};
  ram_1801 = _RAND_1803[7:0];
  _RAND_1804 = {1{`RANDOM}};
  ram_1802 = _RAND_1804[7:0];
  _RAND_1805 = {1{`RANDOM}};
  ram_1803 = _RAND_1805[7:0];
  _RAND_1806 = {1{`RANDOM}};
  ram_1804 = _RAND_1806[7:0];
  _RAND_1807 = {1{`RANDOM}};
  ram_1805 = _RAND_1807[7:0];
  _RAND_1808 = {1{`RANDOM}};
  ram_1806 = _RAND_1808[7:0];
  _RAND_1809 = {1{`RANDOM}};
  ram_1807 = _RAND_1809[7:0];
  _RAND_1810 = {1{`RANDOM}};
  ram_1808 = _RAND_1810[7:0];
  _RAND_1811 = {1{`RANDOM}};
  ram_1809 = _RAND_1811[7:0];
  _RAND_1812 = {1{`RANDOM}};
  ram_1810 = _RAND_1812[7:0];
  _RAND_1813 = {1{`RANDOM}};
  ram_1811 = _RAND_1813[7:0];
  _RAND_1814 = {1{`RANDOM}};
  ram_1812 = _RAND_1814[7:0];
  _RAND_1815 = {1{`RANDOM}};
  ram_1813 = _RAND_1815[7:0];
  _RAND_1816 = {1{`RANDOM}};
  ram_1814 = _RAND_1816[7:0];
  _RAND_1817 = {1{`RANDOM}};
  ram_1815 = _RAND_1817[7:0];
  _RAND_1818 = {1{`RANDOM}};
  ram_1816 = _RAND_1818[7:0];
  _RAND_1819 = {1{`RANDOM}};
  ram_1817 = _RAND_1819[7:0];
  _RAND_1820 = {1{`RANDOM}};
  ram_1818 = _RAND_1820[7:0];
  _RAND_1821 = {1{`RANDOM}};
  ram_1819 = _RAND_1821[7:0];
  _RAND_1822 = {1{`RANDOM}};
  ram_1820 = _RAND_1822[7:0];
  _RAND_1823 = {1{`RANDOM}};
  ram_1821 = _RAND_1823[7:0];
  _RAND_1824 = {1{`RANDOM}};
  ram_1822 = _RAND_1824[7:0];
  _RAND_1825 = {1{`RANDOM}};
  ram_1823 = _RAND_1825[7:0];
  _RAND_1826 = {1{`RANDOM}};
  ram_1824 = _RAND_1826[7:0];
  _RAND_1827 = {1{`RANDOM}};
  ram_1825 = _RAND_1827[7:0];
  _RAND_1828 = {1{`RANDOM}};
  ram_1826 = _RAND_1828[7:0];
  _RAND_1829 = {1{`RANDOM}};
  ram_1827 = _RAND_1829[7:0];
  _RAND_1830 = {1{`RANDOM}};
  ram_1828 = _RAND_1830[7:0];
  _RAND_1831 = {1{`RANDOM}};
  ram_1829 = _RAND_1831[7:0];
  _RAND_1832 = {1{`RANDOM}};
  ram_1830 = _RAND_1832[7:0];
  _RAND_1833 = {1{`RANDOM}};
  ram_1831 = _RAND_1833[7:0];
  _RAND_1834 = {1{`RANDOM}};
  ram_1832 = _RAND_1834[7:0];
  _RAND_1835 = {1{`RANDOM}};
  ram_1833 = _RAND_1835[7:0];
  _RAND_1836 = {1{`RANDOM}};
  ram_1834 = _RAND_1836[7:0];
  _RAND_1837 = {1{`RANDOM}};
  ram_1835 = _RAND_1837[7:0];
  _RAND_1838 = {1{`RANDOM}};
  ram_1836 = _RAND_1838[7:0];
  _RAND_1839 = {1{`RANDOM}};
  ram_1837 = _RAND_1839[7:0];
  _RAND_1840 = {1{`RANDOM}};
  ram_1838 = _RAND_1840[7:0];
  _RAND_1841 = {1{`RANDOM}};
  ram_1839 = _RAND_1841[7:0];
  _RAND_1842 = {1{`RANDOM}};
  ram_1840 = _RAND_1842[7:0];
  _RAND_1843 = {1{`RANDOM}};
  ram_1841 = _RAND_1843[7:0];
  _RAND_1844 = {1{`RANDOM}};
  ram_1842 = _RAND_1844[7:0];
  _RAND_1845 = {1{`RANDOM}};
  ram_1843 = _RAND_1845[7:0];
  _RAND_1846 = {1{`RANDOM}};
  ram_1844 = _RAND_1846[7:0];
  _RAND_1847 = {1{`RANDOM}};
  ram_1845 = _RAND_1847[7:0];
  _RAND_1848 = {1{`RANDOM}};
  ram_1846 = _RAND_1848[7:0];
  _RAND_1849 = {1{`RANDOM}};
  ram_1847 = _RAND_1849[7:0];
  _RAND_1850 = {1{`RANDOM}};
  ram_1848 = _RAND_1850[7:0];
  _RAND_1851 = {1{`RANDOM}};
  ram_1849 = _RAND_1851[7:0];
  _RAND_1852 = {1{`RANDOM}};
  ram_1850 = _RAND_1852[7:0];
  _RAND_1853 = {1{`RANDOM}};
  ram_1851 = _RAND_1853[7:0];
  _RAND_1854 = {1{`RANDOM}};
  ram_1852 = _RAND_1854[7:0];
  _RAND_1855 = {1{`RANDOM}};
  ram_1853 = _RAND_1855[7:0];
  _RAND_1856 = {1{`RANDOM}};
  ram_1854 = _RAND_1856[7:0];
  _RAND_1857 = {1{`RANDOM}};
  ram_1855 = _RAND_1857[7:0];
  _RAND_1858 = {1{`RANDOM}};
  ram_1856 = _RAND_1858[7:0];
  _RAND_1859 = {1{`RANDOM}};
  ram_1857 = _RAND_1859[7:0];
  _RAND_1860 = {1{`RANDOM}};
  ram_1858 = _RAND_1860[7:0];
  _RAND_1861 = {1{`RANDOM}};
  ram_1859 = _RAND_1861[7:0];
  _RAND_1862 = {1{`RANDOM}};
  ram_1860 = _RAND_1862[7:0];
  _RAND_1863 = {1{`RANDOM}};
  ram_1861 = _RAND_1863[7:0];
  _RAND_1864 = {1{`RANDOM}};
  ram_1862 = _RAND_1864[7:0];
  _RAND_1865 = {1{`RANDOM}};
  ram_1863 = _RAND_1865[7:0];
  _RAND_1866 = {1{`RANDOM}};
  ram_1864 = _RAND_1866[7:0];
  _RAND_1867 = {1{`RANDOM}};
  ram_1865 = _RAND_1867[7:0];
  _RAND_1868 = {1{`RANDOM}};
  ram_1866 = _RAND_1868[7:0];
  _RAND_1869 = {1{`RANDOM}};
  ram_1867 = _RAND_1869[7:0];
  _RAND_1870 = {1{`RANDOM}};
  ram_1868 = _RAND_1870[7:0];
  _RAND_1871 = {1{`RANDOM}};
  ram_1869 = _RAND_1871[7:0];
  _RAND_1872 = {1{`RANDOM}};
  ram_1870 = _RAND_1872[7:0];
  _RAND_1873 = {1{`RANDOM}};
  ram_1871 = _RAND_1873[7:0];
  _RAND_1874 = {1{`RANDOM}};
  ram_1872 = _RAND_1874[7:0];
  _RAND_1875 = {1{`RANDOM}};
  ram_1873 = _RAND_1875[7:0];
  _RAND_1876 = {1{`RANDOM}};
  ram_1874 = _RAND_1876[7:0];
  _RAND_1877 = {1{`RANDOM}};
  ram_1875 = _RAND_1877[7:0];
  _RAND_1878 = {1{`RANDOM}};
  ram_1876 = _RAND_1878[7:0];
  _RAND_1879 = {1{`RANDOM}};
  ram_1877 = _RAND_1879[7:0];
  _RAND_1880 = {1{`RANDOM}};
  ram_1878 = _RAND_1880[7:0];
  _RAND_1881 = {1{`RANDOM}};
  ram_1879 = _RAND_1881[7:0];
  _RAND_1882 = {1{`RANDOM}};
  ram_1880 = _RAND_1882[7:0];
  _RAND_1883 = {1{`RANDOM}};
  ram_1881 = _RAND_1883[7:0];
  _RAND_1884 = {1{`RANDOM}};
  ram_1882 = _RAND_1884[7:0];
  _RAND_1885 = {1{`RANDOM}};
  ram_1883 = _RAND_1885[7:0];
  _RAND_1886 = {1{`RANDOM}};
  ram_1884 = _RAND_1886[7:0];
  _RAND_1887 = {1{`RANDOM}};
  ram_1885 = _RAND_1887[7:0];
  _RAND_1888 = {1{`RANDOM}};
  ram_1886 = _RAND_1888[7:0];
  _RAND_1889 = {1{`RANDOM}};
  ram_1887 = _RAND_1889[7:0];
  _RAND_1890 = {1{`RANDOM}};
  ram_1888 = _RAND_1890[7:0];
  _RAND_1891 = {1{`RANDOM}};
  ram_1889 = _RAND_1891[7:0];
  _RAND_1892 = {1{`RANDOM}};
  ram_1890 = _RAND_1892[7:0];
  _RAND_1893 = {1{`RANDOM}};
  ram_1891 = _RAND_1893[7:0];
  _RAND_1894 = {1{`RANDOM}};
  ram_1892 = _RAND_1894[7:0];
  _RAND_1895 = {1{`RANDOM}};
  ram_1893 = _RAND_1895[7:0];
  _RAND_1896 = {1{`RANDOM}};
  ram_1894 = _RAND_1896[7:0];
  _RAND_1897 = {1{`RANDOM}};
  ram_1895 = _RAND_1897[7:0];
  _RAND_1898 = {1{`RANDOM}};
  ram_1896 = _RAND_1898[7:0];
  _RAND_1899 = {1{`RANDOM}};
  ram_1897 = _RAND_1899[7:0];
  _RAND_1900 = {1{`RANDOM}};
  ram_1898 = _RAND_1900[7:0];
  _RAND_1901 = {1{`RANDOM}};
  ram_1899 = _RAND_1901[7:0];
  _RAND_1902 = {1{`RANDOM}};
  ram_1900 = _RAND_1902[7:0];
  _RAND_1903 = {1{`RANDOM}};
  ram_1901 = _RAND_1903[7:0];
  _RAND_1904 = {1{`RANDOM}};
  ram_1902 = _RAND_1904[7:0];
  _RAND_1905 = {1{`RANDOM}};
  ram_1903 = _RAND_1905[7:0];
  _RAND_1906 = {1{`RANDOM}};
  ram_1904 = _RAND_1906[7:0];
  _RAND_1907 = {1{`RANDOM}};
  ram_1905 = _RAND_1907[7:0];
  _RAND_1908 = {1{`RANDOM}};
  ram_1906 = _RAND_1908[7:0];
  _RAND_1909 = {1{`RANDOM}};
  ram_1907 = _RAND_1909[7:0];
  _RAND_1910 = {1{`RANDOM}};
  ram_1908 = _RAND_1910[7:0];
  _RAND_1911 = {1{`RANDOM}};
  ram_1909 = _RAND_1911[7:0];
  _RAND_1912 = {1{`RANDOM}};
  ram_1910 = _RAND_1912[7:0];
  _RAND_1913 = {1{`RANDOM}};
  ram_1911 = _RAND_1913[7:0];
  _RAND_1914 = {1{`RANDOM}};
  ram_1912 = _RAND_1914[7:0];
  _RAND_1915 = {1{`RANDOM}};
  ram_1913 = _RAND_1915[7:0];
  _RAND_1916 = {1{`RANDOM}};
  ram_1914 = _RAND_1916[7:0];
  _RAND_1917 = {1{`RANDOM}};
  ram_1915 = _RAND_1917[7:0];
  _RAND_1918 = {1{`RANDOM}};
  ram_1916 = _RAND_1918[7:0];
  _RAND_1919 = {1{`RANDOM}};
  ram_1917 = _RAND_1919[7:0];
  _RAND_1920 = {1{`RANDOM}};
  ram_1918 = _RAND_1920[7:0];
  _RAND_1921 = {1{`RANDOM}};
  ram_1919 = _RAND_1921[7:0];
  _RAND_1922 = {1{`RANDOM}};
  ram_1920 = _RAND_1922[7:0];
  _RAND_1923 = {1{`RANDOM}};
  ram_1921 = _RAND_1923[7:0];
  _RAND_1924 = {1{`RANDOM}};
  ram_1922 = _RAND_1924[7:0];
  _RAND_1925 = {1{`RANDOM}};
  ram_1923 = _RAND_1925[7:0];
  _RAND_1926 = {1{`RANDOM}};
  ram_1924 = _RAND_1926[7:0];
  _RAND_1927 = {1{`RANDOM}};
  ram_1925 = _RAND_1927[7:0];
  _RAND_1928 = {1{`RANDOM}};
  ram_1926 = _RAND_1928[7:0];
  _RAND_1929 = {1{`RANDOM}};
  ram_1927 = _RAND_1929[7:0];
  _RAND_1930 = {1{`RANDOM}};
  ram_1928 = _RAND_1930[7:0];
  _RAND_1931 = {1{`RANDOM}};
  ram_1929 = _RAND_1931[7:0];
  _RAND_1932 = {1{`RANDOM}};
  ram_1930 = _RAND_1932[7:0];
  _RAND_1933 = {1{`RANDOM}};
  ram_1931 = _RAND_1933[7:0];
  _RAND_1934 = {1{`RANDOM}};
  ram_1932 = _RAND_1934[7:0];
  _RAND_1935 = {1{`RANDOM}};
  ram_1933 = _RAND_1935[7:0];
  _RAND_1936 = {1{`RANDOM}};
  ram_1934 = _RAND_1936[7:0];
  _RAND_1937 = {1{`RANDOM}};
  ram_1935 = _RAND_1937[7:0];
  _RAND_1938 = {1{`RANDOM}};
  ram_1936 = _RAND_1938[7:0];
  _RAND_1939 = {1{`RANDOM}};
  ram_1937 = _RAND_1939[7:0];
  _RAND_1940 = {1{`RANDOM}};
  ram_1938 = _RAND_1940[7:0];
  _RAND_1941 = {1{`RANDOM}};
  ram_1939 = _RAND_1941[7:0];
  _RAND_1942 = {1{`RANDOM}};
  ram_1940 = _RAND_1942[7:0];
  _RAND_1943 = {1{`RANDOM}};
  ram_1941 = _RAND_1943[7:0];
  _RAND_1944 = {1{`RANDOM}};
  ram_1942 = _RAND_1944[7:0];
  _RAND_1945 = {1{`RANDOM}};
  ram_1943 = _RAND_1945[7:0];
  _RAND_1946 = {1{`RANDOM}};
  ram_1944 = _RAND_1946[7:0];
  _RAND_1947 = {1{`RANDOM}};
  ram_1945 = _RAND_1947[7:0];
  _RAND_1948 = {1{`RANDOM}};
  ram_1946 = _RAND_1948[7:0];
  _RAND_1949 = {1{`RANDOM}};
  ram_1947 = _RAND_1949[7:0];
  _RAND_1950 = {1{`RANDOM}};
  ram_1948 = _RAND_1950[7:0];
  _RAND_1951 = {1{`RANDOM}};
  ram_1949 = _RAND_1951[7:0];
  _RAND_1952 = {1{`RANDOM}};
  ram_1950 = _RAND_1952[7:0];
  _RAND_1953 = {1{`RANDOM}};
  ram_1951 = _RAND_1953[7:0];
  _RAND_1954 = {1{`RANDOM}};
  ram_1952 = _RAND_1954[7:0];
  _RAND_1955 = {1{`RANDOM}};
  ram_1953 = _RAND_1955[7:0];
  _RAND_1956 = {1{`RANDOM}};
  ram_1954 = _RAND_1956[7:0];
  _RAND_1957 = {1{`RANDOM}};
  ram_1955 = _RAND_1957[7:0];
  _RAND_1958 = {1{`RANDOM}};
  ram_1956 = _RAND_1958[7:0];
  _RAND_1959 = {1{`RANDOM}};
  ram_1957 = _RAND_1959[7:0];
  _RAND_1960 = {1{`RANDOM}};
  ram_1958 = _RAND_1960[7:0];
  _RAND_1961 = {1{`RANDOM}};
  ram_1959 = _RAND_1961[7:0];
  _RAND_1962 = {1{`RANDOM}};
  ram_1960 = _RAND_1962[7:0];
  _RAND_1963 = {1{`RANDOM}};
  ram_1961 = _RAND_1963[7:0];
  _RAND_1964 = {1{`RANDOM}};
  ram_1962 = _RAND_1964[7:0];
  _RAND_1965 = {1{`RANDOM}};
  ram_1963 = _RAND_1965[7:0];
  _RAND_1966 = {1{`RANDOM}};
  ram_1964 = _RAND_1966[7:0];
  _RAND_1967 = {1{`RANDOM}};
  ram_1965 = _RAND_1967[7:0];
  _RAND_1968 = {1{`RANDOM}};
  ram_1966 = _RAND_1968[7:0];
  _RAND_1969 = {1{`RANDOM}};
  ram_1967 = _RAND_1969[7:0];
  _RAND_1970 = {1{`RANDOM}};
  ram_1968 = _RAND_1970[7:0];
  _RAND_1971 = {1{`RANDOM}};
  ram_1969 = _RAND_1971[7:0];
  _RAND_1972 = {1{`RANDOM}};
  ram_1970 = _RAND_1972[7:0];
  _RAND_1973 = {1{`RANDOM}};
  ram_1971 = _RAND_1973[7:0];
  _RAND_1974 = {1{`RANDOM}};
  ram_1972 = _RAND_1974[7:0];
  _RAND_1975 = {1{`RANDOM}};
  ram_1973 = _RAND_1975[7:0];
  _RAND_1976 = {1{`RANDOM}};
  ram_1974 = _RAND_1976[7:0];
  _RAND_1977 = {1{`RANDOM}};
  ram_1975 = _RAND_1977[7:0];
  _RAND_1978 = {1{`RANDOM}};
  ram_1976 = _RAND_1978[7:0];
  _RAND_1979 = {1{`RANDOM}};
  ram_1977 = _RAND_1979[7:0];
  _RAND_1980 = {1{`RANDOM}};
  ram_1978 = _RAND_1980[7:0];
  _RAND_1981 = {1{`RANDOM}};
  ram_1979 = _RAND_1981[7:0];
  _RAND_1982 = {1{`RANDOM}};
  ram_1980 = _RAND_1982[7:0];
  _RAND_1983 = {1{`RANDOM}};
  ram_1981 = _RAND_1983[7:0];
  _RAND_1984 = {1{`RANDOM}};
  ram_1982 = _RAND_1984[7:0];
  _RAND_1985 = {1{`RANDOM}};
  ram_1983 = _RAND_1985[7:0];
  _RAND_1986 = {1{`RANDOM}};
  ram_1984 = _RAND_1986[7:0];
  _RAND_1987 = {1{`RANDOM}};
  ram_1985 = _RAND_1987[7:0];
  _RAND_1988 = {1{`RANDOM}};
  ram_1986 = _RAND_1988[7:0];
  _RAND_1989 = {1{`RANDOM}};
  ram_1987 = _RAND_1989[7:0];
  _RAND_1990 = {1{`RANDOM}};
  ram_1988 = _RAND_1990[7:0];
  _RAND_1991 = {1{`RANDOM}};
  ram_1989 = _RAND_1991[7:0];
  _RAND_1992 = {1{`RANDOM}};
  ram_1990 = _RAND_1992[7:0];
  _RAND_1993 = {1{`RANDOM}};
  ram_1991 = _RAND_1993[7:0];
  _RAND_1994 = {1{`RANDOM}};
  ram_1992 = _RAND_1994[7:0];
  _RAND_1995 = {1{`RANDOM}};
  ram_1993 = _RAND_1995[7:0];
  _RAND_1996 = {1{`RANDOM}};
  ram_1994 = _RAND_1996[7:0];
  _RAND_1997 = {1{`RANDOM}};
  ram_1995 = _RAND_1997[7:0];
  _RAND_1998 = {1{`RANDOM}};
  ram_1996 = _RAND_1998[7:0];
  _RAND_1999 = {1{`RANDOM}};
  ram_1997 = _RAND_1999[7:0];
  _RAND_2000 = {1{`RANDOM}};
  ram_1998 = _RAND_2000[7:0];
  _RAND_2001 = {1{`RANDOM}};
  ram_1999 = _RAND_2001[7:0];
  _RAND_2002 = {1{`RANDOM}};
  ram_2000 = _RAND_2002[7:0];
  _RAND_2003 = {1{`RANDOM}};
  ram_2001 = _RAND_2003[7:0];
  _RAND_2004 = {1{`RANDOM}};
  ram_2002 = _RAND_2004[7:0];
  _RAND_2005 = {1{`RANDOM}};
  ram_2003 = _RAND_2005[7:0];
  _RAND_2006 = {1{`RANDOM}};
  ram_2004 = _RAND_2006[7:0];
  _RAND_2007 = {1{`RANDOM}};
  ram_2005 = _RAND_2007[7:0];
  _RAND_2008 = {1{`RANDOM}};
  ram_2006 = _RAND_2008[7:0];
  _RAND_2009 = {1{`RANDOM}};
  ram_2007 = _RAND_2009[7:0];
  _RAND_2010 = {1{`RANDOM}};
  ram_2008 = _RAND_2010[7:0];
  _RAND_2011 = {1{`RANDOM}};
  ram_2009 = _RAND_2011[7:0];
  _RAND_2012 = {1{`RANDOM}};
  ram_2010 = _RAND_2012[7:0];
  _RAND_2013 = {1{`RANDOM}};
  ram_2011 = _RAND_2013[7:0];
  _RAND_2014 = {1{`RANDOM}};
  ram_2012 = _RAND_2014[7:0];
  _RAND_2015 = {1{`RANDOM}};
  ram_2013 = _RAND_2015[7:0];
  _RAND_2016 = {1{`RANDOM}};
  ram_2014 = _RAND_2016[7:0];
  _RAND_2017 = {1{`RANDOM}};
  ram_2015 = _RAND_2017[7:0];
  _RAND_2018 = {1{`RANDOM}};
  ram_2016 = _RAND_2018[7:0];
  _RAND_2019 = {1{`RANDOM}};
  ram_2017 = _RAND_2019[7:0];
  _RAND_2020 = {1{`RANDOM}};
  ram_2018 = _RAND_2020[7:0];
  _RAND_2021 = {1{`RANDOM}};
  ram_2019 = _RAND_2021[7:0];
  _RAND_2022 = {1{`RANDOM}};
  ram_2020 = _RAND_2022[7:0];
  _RAND_2023 = {1{`RANDOM}};
  ram_2021 = _RAND_2023[7:0];
  _RAND_2024 = {1{`RANDOM}};
  ram_2022 = _RAND_2024[7:0];
  _RAND_2025 = {1{`RANDOM}};
  ram_2023 = _RAND_2025[7:0];
  _RAND_2026 = {1{`RANDOM}};
  ram_2024 = _RAND_2026[7:0];
  _RAND_2027 = {1{`RANDOM}};
  ram_2025 = _RAND_2027[7:0];
  _RAND_2028 = {1{`RANDOM}};
  ram_2026 = _RAND_2028[7:0];
  _RAND_2029 = {1{`RANDOM}};
  ram_2027 = _RAND_2029[7:0];
  _RAND_2030 = {1{`RANDOM}};
  ram_2028 = _RAND_2030[7:0];
  _RAND_2031 = {1{`RANDOM}};
  ram_2029 = _RAND_2031[7:0];
  _RAND_2032 = {1{`RANDOM}};
  ram_2030 = _RAND_2032[7:0];
  _RAND_2033 = {1{`RANDOM}};
  ram_2031 = _RAND_2033[7:0];
  _RAND_2034 = {1{`RANDOM}};
  ram_2032 = _RAND_2034[7:0];
  _RAND_2035 = {1{`RANDOM}};
  ram_2033 = _RAND_2035[7:0];
  _RAND_2036 = {1{`RANDOM}};
  ram_2034 = _RAND_2036[7:0];
  _RAND_2037 = {1{`RANDOM}};
  ram_2035 = _RAND_2037[7:0];
  _RAND_2038 = {1{`RANDOM}};
  ram_2036 = _RAND_2038[7:0];
  _RAND_2039 = {1{`RANDOM}};
  ram_2037 = _RAND_2039[7:0];
  _RAND_2040 = {1{`RANDOM}};
  ram_2038 = _RAND_2040[7:0];
  _RAND_2041 = {1{`RANDOM}};
  ram_2039 = _RAND_2041[7:0];
  _RAND_2042 = {1{`RANDOM}};
  ram_2040 = _RAND_2042[7:0];
  _RAND_2043 = {1{`RANDOM}};
  ram_2041 = _RAND_2043[7:0];
  _RAND_2044 = {1{`RANDOM}};
  ram_2042 = _RAND_2044[7:0];
  _RAND_2045 = {1{`RANDOM}};
  ram_2043 = _RAND_2045[7:0];
  _RAND_2046 = {1{`RANDOM}};
  ram_2044 = _RAND_2046[7:0];
  _RAND_2047 = {1{`RANDOM}};
  ram_2045 = _RAND_2047[7:0];
  _RAND_2048 = {1{`RANDOM}};
  ram_2046 = _RAND_2048[7:0];
  _RAND_2049 = {1{`RANDOM}};
  ram_2047 = _RAND_2049[7:0];
  _RAND_2050 = {1{`RANDOM}};
  ram_2048 = _RAND_2050[7:0];
  _RAND_2051 = {1{`RANDOM}};
  ram_2049 = _RAND_2051[7:0];
  _RAND_2052 = {1{`RANDOM}};
  ram_2050 = _RAND_2052[7:0];
  _RAND_2053 = {1{`RANDOM}};
  ram_2051 = _RAND_2053[7:0];
  _RAND_2054 = {1{`RANDOM}};
  ram_2052 = _RAND_2054[7:0];
  _RAND_2055 = {1{`RANDOM}};
  ram_2053 = _RAND_2055[7:0];
  _RAND_2056 = {1{`RANDOM}};
  ram_2054 = _RAND_2056[7:0];
  _RAND_2057 = {1{`RANDOM}};
  ram_2055 = _RAND_2057[7:0];
  _RAND_2058 = {1{`RANDOM}};
  ram_2056 = _RAND_2058[7:0];
  _RAND_2059 = {1{`RANDOM}};
  ram_2057 = _RAND_2059[7:0];
  _RAND_2060 = {1{`RANDOM}};
  ram_2058 = _RAND_2060[7:0];
  _RAND_2061 = {1{`RANDOM}};
  ram_2059 = _RAND_2061[7:0];
  _RAND_2062 = {1{`RANDOM}};
  ram_2060 = _RAND_2062[7:0];
  _RAND_2063 = {1{`RANDOM}};
  ram_2061 = _RAND_2063[7:0];
  _RAND_2064 = {1{`RANDOM}};
  ram_2062 = _RAND_2064[7:0];
  _RAND_2065 = {1{`RANDOM}};
  ram_2063 = _RAND_2065[7:0];
  _RAND_2066 = {1{`RANDOM}};
  ram_2064 = _RAND_2066[7:0];
  _RAND_2067 = {1{`RANDOM}};
  ram_2065 = _RAND_2067[7:0];
  _RAND_2068 = {1{`RANDOM}};
  ram_2066 = _RAND_2068[7:0];
  _RAND_2069 = {1{`RANDOM}};
  ram_2067 = _RAND_2069[7:0];
  _RAND_2070 = {1{`RANDOM}};
  ram_2068 = _RAND_2070[7:0];
  _RAND_2071 = {1{`RANDOM}};
  ram_2069 = _RAND_2071[7:0];
  _RAND_2072 = {1{`RANDOM}};
  ram_2070 = _RAND_2072[7:0];
  _RAND_2073 = {1{`RANDOM}};
  ram_2071 = _RAND_2073[7:0];
  _RAND_2074 = {1{`RANDOM}};
  ram_2072 = _RAND_2074[7:0];
  _RAND_2075 = {1{`RANDOM}};
  ram_2073 = _RAND_2075[7:0];
  _RAND_2076 = {1{`RANDOM}};
  ram_2074 = _RAND_2076[7:0];
  _RAND_2077 = {1{`RANDOM}};
  ram_2075 = _RAND_2077[7:0];
  _RAND_2078 = {1{`RANDOM}};
  ram_2076 = _RAND_2078[7:0];
  _RAND_2079 = {1{`RANDOM}};
  ram_2077 = _RAND_2079[7:0];
  _RAND_2080 = {1{`RANDOM}};
  ram_2078 = _RAND_2080[7:0];
  _RAND_2081 = {1{`RANDOM}};
  ram_2079 = _RAND_2081[7:0];
  _RAND_2082 = {1{`RANDOM}};
  ram_2080 = _RAND_2082[7:0];
  _RAND_2083 = {1{`RANDOM}};
  ram_2081 = _RAND_2083[7:0];
  _RAND_2084 = {1{`RANDOM}};
  ram_2082 = _RAND_2084[7:0];
  _RAND_2085 = {1{`RANDOM}};
  ram_2083 = _RAND_2085[7:0];
  _RAND_2086 = {1{`RANDOM}};
  ram_2084 = _RAND_2086[7:0];
  _RAND_2087 = {1{`RANDOM}};
  ram_2085 = _RAND_2087[7:0];
  _RAND_2088 = {1{`RANDOM}};
  ram_2086 = _RAND_2088[7:0];
  _RAND_2089 = {1{`RANDOM}};
  ram_2087 = _RAND_2089[7:0];
  _RAND_2090 = {1{`RANDOM}};
  ram_2088 = _RAND_2090[7:0];
  _RAND_2091 = {1{`RANDOM}};
  ram_2089 = _RAND_2091[7:0];
  _RAND_2092 = {1{`RANDOM}};
  ram_2090 = _RAND_2092[7:0];
  _RAND_2093 = {1{`RANDOM}};
  ram_2091 = _RAND_2093[7:0];
  _RAND_2094 = {1{`RANDOM}};
  ram_2092 = _RAND_2094[7:0];
  _RAND_2095 = {1{`RANDOM}};
  ram_2093 = _RAND_2095[7:0];
  _RAND_2096 = {1{`RANDOM}};
  ram_2094 = _RAND_2096[7:0];
  _RAND_2097 = {1{`RANDOM}};
  ram_2095 = _RAND_2097[7:0];
  _RAND_2098 = {1{`RANDOM}};
  ram_2096 = _RAND_2098[7:0];
  _RAND_2099 = {1{`RANDOM}};
  ram_2097 = _RAND_2099[7:0];
  _RAND_2100 = {1{`RANDOM}};
  ram_2098 = _RAND_2100[7:0];
  _RAND_2101 = {1{`RANDOM}};
  ram_2099 = _RAND_2101[7:0];
  _RAND_2102 = {1{`RANDOM}};
  ram_2100 = _RAND_2102[7:0];
  _RAND_2103 = {1{`RANDOM}};
  ram_2101 = _RAND_2103[7:0];
  _RAND_2104 = {1{`RANDOM}};
  ram_2102 = _RAND_2104[7:0];
  _RAND_2105 = {1{`RANDOM}};
  ram_2103 = _RAND_2105[7:0];
  _RAND_2106 = {1{`RANDOM}};
  ram_2104 = _RAND_2106[7:0];
  _RAND_2107 = {1{`RANDOM}};
  ram_2105 = _RAND_2107[7:0];
  _RAND_2108 = {1{`RANDOM}};
  ram_2106 = _RAND_2108[7:0];
  _RAND_2109 = {1{`RANDOM}};
  ram_2107 = _RAND_2109[7:0];
  _RAND_2110 = {1{`RANDOM}};
  ram_2108 = _RAND_2110[7:0];
  _RAND_2111 = {1{`RANDOM}};
  ram_2109 = _RAND_2111[7:0];
  _RAND_2112 = {1{`RANDOM}};
  ram_2110 = _RAND_2112[7:0];
  _RAND_2113 = {1{`RANDOM}};
  ram_2111 = _RAND_2113[7:0];
  _RAND_2114 = {1{`RANDOM}};
  ram_2112 = _RAND_2114[7:0];
  _RAND_2115 = {1{`RANDOM}};
  ram_2113 = _RAND_2115[7:0];
  _RAND_2116 = {1{`RANDOM}};
  ram_2114 = _RAND_2116[7:0];
  _RAND_2117 = {1{`RANDOM}};
  ram_2115 = _RAND_2117[7:0];
  _RAND_2118 = {1{`RANDOM}};
  ram_2116 = _RAND_2118[7:0];
  _RAND_2119 = {1{`RANDOM}};
  ram_2117 = _RAND_2119[7:0];
  _RAND_2120 = {1{`RANDOM}};
  ram_2118 = _RAND_2120[7:0];
  _RAND_2121 = {1{`RANDOM}};
  ram_2119 = _RAND_2121[7:0];
  _RAND_2122 = {1{`RANDOM}};
  ram_2120 = _RAND_2122[7:0];
  _RAND_2123 = {1{`RANDOM}};
  ram_2121 = _RAND_2123[7:0];
  _RAND_2124 = {1{`RANDOM}};
  ram_2122 = _RAND_2124[7:0];
  _RAND_2125 = {1{`RANDOM}};
  ram_2123 = _RAND_2125[7:0];
  _RAND_2126 = {1{`RANDOM}};
  ram_2124 = _RAND_2126[7:0];
  _RAND_2127 = {1{`RANDOM}};
  ram_2125 = _RAND_2127[7:0];
  _RAND_2128 = {1{`RANDOM}};
  ram_2126 = _RAND_2128[7:0];
  _RAND_2129 = {1{`RANDOM}};
  ram_2127 = _RAND_2129[7:0];
  _RAND_2130 = {1{`RANDOM}};
  ram_2128 = _RAND_2130[7:0];
  _RAND_2131 = {1{`RANDOM}};
  ram_2129 = _RAND_2131[7:0];
  _RAND_2132 = {1{`RANDOM}};
  ram_2130 = _RAND_2132[7:0];
  _RAND_2133 = {1{`RANDOM}};
  ram_2131 = _RAND_2133[7:0];
  _RAND_2134 = {1{`RANDOM}};
  ram_2132 = _RAND_2134[7:0];
  _RAND_2135 = {1{`RANDOM}};
  ram_2133 = _RAND_2135[7:0];
  _RAND_2136 = {1{`RANDOM}};
  ram_2134 = _RAND_2136[7:0];
  _RAND_2137 = {1{`RANDOM}};
  ram_2135 = _RAND_2137[7:0];
  _RAND_2138 = {1{`RANDOM}};
  ram_2136 = _RAND_2138[7:0];
  _RAND_2139 = {1{`RANDOM}};
  ram_2137 = _RAND_2139[7:0];
  _RAND_2140 = {1{`RANDOM}};
  ram_2138 = _RAND_2140[7:0];
  _RAND_2141 = {1{`RANDOM}};
  ram_2139 = _RAND_2141[7:0];
  _RAND_2142 = {1{`RANDOM}};
  ram_2140 = _RAND_2142[7:0];
  _RAND_2143 = {1{`RANDOM}};
  ram_2141 = _RAND_2143[7:0];
  _RAND_2144 = {1{`RANDOM}};
  ram_2142 = _RAND_2144[7:0];
  _RAND_2145 = {1{`RANDOM}};
  ram_2143 = _RAND_2145[7:0];
  _RAND_2146 = {1{`RANDOM}};
  ram_2144 = _RAND_2146[7:0];
  _RAND_2147 = {1{`RANDOM}};
  ram_2145 = _RAND_2147[7:0];
  _RAND_2148 = {1{`RANDOM}};
  ram_2146 = _RAND_2148[7:0];
  _RAND_2149 = {1{`RANDOM}};
  ram_2147 = _RAND_2149[7:0];
  _RAND_2150 = {1{`RANDOM}};
  ram_2148 = _RAND_2150[7:0];
  _RAND_2151 = {1{`RANDOM}};
  ram_2149 = _RAND_2151[7:0];
  _RAND_2152 = {1{`RANDOM}};
  ram_2150 = _RAND_2152[7:0];
  _RAND_2153 = {1{`RANDOM}};
  ram_2151 = _RAND_2153[7:0];
  _RAND_2154 = {1{`RANDOM}};
  ram_2152 = _RAND_2154[7:0];
  _RAND_2155 = {1{`RANDOM}};
  ram_2153 = _RAND_2155[7:0];
  _RAND_2156 = {1{`RANDOM}};
  ram_2154 = _RAND_2156[7:0];
  _RAND_2157 = {1{`RANDOM}};
  ram_2155 = _RAND_2157[7:0];
  _RAND_2158 = {1{`RANDOM}};
  ram_2156 = _RAND_2158[7:0];
  _RAND_2159 = {1{`RANDOM}};
  ram_2157 = _RAND_2159[7:0];
  _RAND_2160 = {1{`RANDOM}};
  ram_2158 = _RAND_2160[7:0];
  _RAND_2161 = {1{`RANDOM}};
  ram_2159 = _RAND_2161[7:0];
  _RAND_2162 = {1{`RANDOM}};
  ram_2160 = _RAND_2162[7:0];
  _RAND_2163 = {1{`RANDOM}};
  index = _RAND_2163[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
  $readmemh("resource/vga_font.txt", vga_mem);
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vga_ctrl(
  input         clock,
  input         reset,
  input  [23:0] io_vga_data,
  output [9:0]  io_h_addr,
  output [9:0]  io_v_addr,
  output        io_hsync,
  output        io_vsync,
  output        io_valid,
  output [7:0]  io_vga_r,
  output [7:0]  io_vga_g,
  output [7:0]  io_vga_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] x_cnt; // @[vga.scala 60:22]
  reg [9:0] y_cnt; // @[vga.scala 61:22]
  wire  _T = x_cnt == 10'h320; // @[vga.scala 63:15]
  wire [9:0] _x_cnt_T_1 = x_cnt + 10'h1; // @[vga.scala 66:21]
  wire [9:0] _y_cnt_T_1 = y_cnt + 10'h1; // @[vga.scala 71:21]
  wire  h_valid = x_cnt > 10'h90 & x_cnt <= 10'h310; // @[vga.scala 75:39]
  wire  v_valid = y_cnt > 10'h23 & y_cnt <= 10'h203; // @[vga.scala 76:39]
  wire [9:0] _io_h_addr_T_1 = x_cnt - 10'h91; // @[vga.scala 78:33]
  wire [9:0] _io_v_addr_T_1 = y_cnt - 10'h24; // @[vga.scala 79:33]
  assign io_h_addr = h_valid ? _io_h_addr_T_1 : 10'h0; // @[vga.scala 78:19]
  assign io_v_addr = v_valid ? _io_v_addr_T_1 : 10'h0; // @[vga.scala 79:19]
  assign io_hsync = x_cnt > 10'h60; // @[vga.scala 73:21]
  assign io_vsync = y_cnt > 10'h2; // @[vga.scala 74:21]
  assign io_valid = h_valid & v_valid; // @[vga.scala 77:23]
  assign io_vga_r = io_vga_data[23:16]; // @[vga.scala 80:26]
  assign io_vga_g = io_vga_data[15:8]; // @[vga.scala 81:26]
  assign io_vga_b = io_vga_data[7:0]; // @[vga.scala 82:26]
  always @(posedge clock) begin
    if (reset) begin // @[vga.scala 60:22]
      x_cnt <= 10'h1; // @[vga.scala 60:22]
    end else if (x_cnt == 10'h320) begin // @[vga.scala 63:26]
      x_cnt <= 10'h1; // @[vga.scala 64:14]
    end else begin
      x_cnt <= _x_cnt_T_1; // @[vga.scala 66:14]
    end
    if (reset) begin // @[vga.scala 61:22]
      y_cnt <= 10'h1; // @[vga.scala 61:22]
    end else if (y_cnt == 10'h20d & _T) begin // @[vga.scala 68:47]
      y_cnt <= 10'h1; // @[vga.scala 69:14]
    end else if (_T) begin // @[vga.scala 70:32]
      y_cnt <= _y_cnt_T_1; // @[vga.scala 71:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_cnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  y_cnt = _RAND_1[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input        clock,
  input        reset,
  input        io_ps2_clk,
  input        io_ps2_data,
  output       io_VGA_HSYNC,
  output       io_VGA_VSYNC,
  output       io_VGA_BLANK_N,
  output [7:0] io_VGA_R,
  output [7:0] io_VGA_G,
  output [7:0] io_VGA_B,
  output [7:0] io_bcd8seg_0,
  output [7:0] io_bcd8seg_1,
  output [7:0] io_bcd8seg_2,
  output [7:0] io_bcd8seg_3,
  output [7:0] io_bcd8seg_4,
  output [7:0] io_bcd8seg_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  PS2_clock; // @[top.scala 19:19]
  wire  PS2_reset; // @[top.scala 19:19]
  wire  PS2_io_ps2_clk; // @[top.scala 19:19]
  wire  PS2_io_ps2_data; // @[top.scala 19:19]
  wire [7:0] PS2_io_ascii; // @[top.scala 19:19]
  wire  PS2_io_ready; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_0; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_1; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_2; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_3; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_4; // @[top.scala 19:19]
  wire [7:0] PS2_io_bcd8seg_5; // @[top.scala 19:19]
  wire  vm_clock; // @[top.scala 25:18]
  wire  vm_reset; // @[top.scala 25:18]
  wire [9:0] vm_io_h_addr; // @[top.scala 25:18]
  wire [8:0] vm_io_v_addr; // @[top.scala 25:18]
  wire [7:0] vm_io_ascii; // @[top.scala 25:18]
  wire  vm_io_w_en; // @[top.scala 25:18]
  wire [23:0] vm_io_vga_data; // @[top.scala 25:18]
  wire  vc_clock; // @[top.scala 26:18]
  wire  vc_reset; // @[top.scala 26:18]
  wire [23:0] vc_io_vga_data; // @[top.scala 26:18]
  wire [9:0] vc_io_h_addr; // @[top.scala 26:18]
  wire [9:0] vc_io_v_addr; // @[top.scala 26:18]
  wire  vc_io_hsync; // @[top.scala 26:18]
  wire  vc_io_vsync; // @[top.scala 26:18]
  wire  vc_io_valid; // @[top.scala 26:18]
  wire [7:0] vc_io_vga_r; // @[top.scala 26:18]
  wire [7:0] vc_io_vga_g; // @[top.scala 26:18]
  wire [7:0] vc_io_vga_b; // @[top.scala 26:18]
  reg [7:0] ascii; // @[top.scala 17:22]
  reg  ready; // @[top.scala 18:22]
  ps2 PS2 ( // @[top.scala 19:19]
    .clock(PS2_clock),
    .reset(PS2_reset),
    .io_ps2_clk(PS2_io_ps2_clk),
    .io_ps2_data(PS2_io_ps2_data),
    .io_ascii(PS2_io_ascii),
    .io_ready(PS2_io_ready),
    .io_bcd8seg_0(PS2_io_bcd8seg_0),
    .io_bcd8seg_1(PS2_io_bcd8seg_1),
    .io_bcd8seg_2(PS2_io_bcd8seg_2),
    .io_bcd8seg_3(PS2_io_bcd8seg_3),
    .io_bcd8seg_4(PS2_io_bcd8seg_4),
    .io_bcd8seg_5(PS2_io_bcd8seg_5)
  );
  vmem vm ( // @[top.scala 25:18]
    .clock(vm_clock),
    .reset(vm_reset),
    .io_h_addr(vm_io_h_addr),
    .io_v_addr(vm_io_v_addr),
    .io_ascii(vm_io_ascii),
    .io_w_en(vm_io_w_en),
    .io_vga_data(vm_io_vga_data)
  );
  vga_ctrl vc ( // @[top.scala 26:18]
    .clock(vc_clock),
    .reset(vc_reset),
    .io_vga_data(vc_io_vga_data),
    .io_h_addr(vc_io_h_addr),
    .io_v_addr(vc_io_v_addr),
    .io_hsync(vc_io_hsync),
    .io_vsync(vc_io_vsync),
    .io_valid(vc_io_valid),
    .io_vga_r(vc_io_vga_r),
    .io_vga_g(vc_io_vga_g),
    .io_vga_b(vc_io_vga_b)
  );
  assign io_VGA_HSYNC = vc_io_hsync; // @[top.scala 32:17]
  assign io_VGA_VSYNC = vc_io_vsync; // @[top.scala 33:17]
  assign io_VGA_BLANK_N = vc_io_valid; // @[top.scala 37:19]
  assign io_VGA_R = vc_io_vga_r; // @[top.scala 34:13]
  assign io_VGA_G = vc_io_vga_g; // @[top.scala 35:13]
  assign io_VGA_B = vc_io_vga_b; // @[top.scala 36:13]
  assign io_bcd8seg_0 = PS2_io_bcd8seg_0; // @[top.scala 24:15]
  assign io_bcd8seg_1 = PS2_io_bcd8seg_1; // @[top.scala 24:15]
  assign io_bcd8seg_2 = PS2_io_bcd8seg_2; // @[top.scala 24:15]
  assign io_bcd8seg_3 = PS2_io_bcd8seg_3; // @[top.scala 24:15]
  assign io_bcd8seg_4 = PS2_io_bcd8seg_4; // @[top.scala 24:15]
  assign io_bcd8seg_5 = PS2_io_bcd8seg_5; // @[top.scala 24:15]
  assign PS2_clock = clock;
  assign PS2_reset = reset;
  assign PS2_io_ps2_clk = io_ps2_clk; // @[top.scala 20:19]
  assign PS2_io_ps2_data = io_ps2_data; // @[top.scala 21:20]
  assign vm_clock = clock;
  assign vm_reset = reset;
  assign vm_io_h_addr = vc_io_h_addr; // @[top.scala 29:17]
  assign vm_io_v_addr = vc_io_v_addr[8:0]; // @[top.scala 30:17]
  assign vm_io_ascii = ready ? ascii : 8'h0; // @[top.scala 38:22 top.scala 39:20 top.scala 27:16]
  assign vm_io_w_en = ready; // @[top.scala 38:22 top.scala 40:19 top.scala 28:15]
  assign vc_clock = clock;
  assign vc_reset = reset;
  assign vc_io_vga_data = vm_io_vga_data; // @[top.scala 31:19]
  always @(posedge clock) begin
    if (reset) begin // @[top.scala 17:22]
      ascii <= 8'h0; // @[top.scala 17:22]
    end else begin
      ascii <= PS2_io_ascii; // @[top.scala 22:10]
    end
    if (reset) begin // @[top.scala 18:22]
      ready <= 1'h0; // @[top.scala 18:22]
    end else begin
      ready <= PS2_io_ready; // @[top.scala 23:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ascii = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  ready = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
