module DCache(
  input          clock,
  input          reset,
  output         io_in_ar_ready,
  input          io_in_ar_valid,
  input  [31:0]  io_in_ar_bits_addr,
  output         io_in_r_valid,
  output [63:0]  io_in_r_bits_data,
  output         io_in_aw_ready,
  input          io_in_aw_valid,
  input  [31:0]  io_in_aw_bits_addr,
  output         io_in_w_ready,
  input          io_in_w_valid,
  input  [63:0]  io_in_w_bits_data,
  input  [7:0]   io_in_w_bits_strb,
  output         io_in_b_valid,
  input          io_mem_ar_ready,
  output         io_mem_ar_valid,
  output [31:0]  io_mem_ar_bits_addr,
  output [7:0]   io_mem_ar_bits_len,
  output         io_mem_r_ready,
  input          io_mem_r_valid,
  input  [63:0]  io_mem_r_bits_data,
  input          io_mem_aw_ready,
  output         io_mem_aw_valid,
  output [31:0]  io_mem_aw_bits_addr,
  input          io_mem_w_ready,
  output         io_mem_w_valid,
  output [63:0]  io_mem_w_bits_data,
  output [7:0]   io_mem_w_bits_strb,
  output         io_mem_w_bits_last,
  output         io_mem_b_ready,
  input          io_mem_b_valid,
  input  [127:0] io_ram_bits_Q0,
  input  [127:0] io_ram_bits_Q1,
  output         io_ram_bits_WEN,
  output [127:0] io_ram_bits_BWEN,
  output [6:0]   io_ram_bits_A,
  output [127:0] io_ram_bits_D,
  output         io_ram_bits_WAY,
  input          io_flush,
  output [63:0]  io_hitrate,
  input          io_uncache
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [127:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [63:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
`endif // RANDOMIZE_REG_INIT
  wire  lfsr8_clock; // @[dcache.scala 65:21]
  wire  lfsr8_reset; // @[dcache.scala 65:21]
  wire  lfsr8_io_en; // @[dcache.scala 65:21]
  wire [7:0] lfsr8_io_out; // @[dcache.scala 65:21]
  reg [41:0] cache_tag_0; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_1; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_2; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_3; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_4; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_5; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_6; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_7; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_8; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_9; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_10; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_11; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_12; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_13; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_14; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_15; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_16; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_17; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_18; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_19; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_20; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_21; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_22; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_23; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_24; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_25; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_26; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_27; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_28; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_29; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_30; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_31; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_32; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_33; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_34; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_35; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_36; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_37; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_38; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_39; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_40; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_41; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_42; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_43; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_44; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_45; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_46; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_47; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_48; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_49; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_50; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_51; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_52; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_53; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_54; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_55; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_56; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_57; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_58; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_59; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_60; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_61; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_62; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_63; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_64; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_65; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_66; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_67; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_68; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_69; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_70; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_71; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_72; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_73; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_74; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_75; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_76; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_77; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_78; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_79; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_80; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_81; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_82; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_83; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_84; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_85; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_86; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_87; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_88; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_89; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_90; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_91; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_92; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_93; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_94; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_95; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_96; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_97; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_98; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_99; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_100; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_101; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_102; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_103; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_104; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_105; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_106; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_107; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_108; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_109; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_110; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_111; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_112; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_113; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_114; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_115; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_116; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_117; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_118; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_119; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_120; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_121; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_122; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_123; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_124; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_125; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_126; // @[dcache.scala 29:26]
  reg [41:0] cache_tag_127; // @[dcache.scala 29:26]
  reg  valid_0_0; // @[dcache.scala 30:22]
  reg  valid_0_1; // @[dcache.scala 30:22]
  reg  valid_1_0; // @[dcache.scala 30:22]
  reg  valid_1_1; // @[dcache.scala 30:22]
  reg  valid_2_0; // @[dcache.scala 30:22]
  reg  valid_2_1; // @[dcache.scala 30:22]
  reg  valid_3_0; // @[dcache.scala 30:22]
  reg  valid_3_1; // @[dcache.scala 30:22]
  reg  valid_4_0; // @[dcache.scala 30:22]
  reg  valid_4_1; // @[dcache.scala 30:22]
  reg  valid_5_0; // @[dcache.scala 30:22]
  reg  valid_5_1; // @[dcache.scala 30:22]
  reg  valid_6_0; // @[dcache.scala 30:22]
  reg  valid_6_1; // @[dcache.scala 30:22]
  reg  valid_7_0; // @[dcache.scala 30:22]
  reg  valid_7_1; // @[dcache.scala 30:22]
  reg  valid_8_0; // @[dcache.scala 30:22]
  reg  valid_8_1; // @[dcache.scala 30:22]
  reg  valid_9_0; // @[dcache.scala 30:22]
  reg  valid_9_1; // @[dcache.scala 30:22]
  reg  valid_10_0; // @[dcache.scala 30:22]
  reg  valid_10_1; // @[dcache.scala 30:22]
  reg  valid_11_0; // @[dcache.scala 30:22]
  reg  valid_11_1; // @[dcache.scala 30:22]
  reg  valid_12_0; // @[dcache.scala 30:22]
  reg  valid_12_1; // @[dcache.scala 30:22]
  reg  valid_13_0; // @[dcache.scala 30:22]
  reg  valid_13_1; // @[dcache.scala 30:22]
  reg  valid_14_0; // @[dcache.scala 30:22]
  reg  valid_14_1; // @[dcache.scala 30:22]
  reg  valid_15_0; // @[dcache.scala 30:22]
  reg  valid_15_1; // @[dcache.scala 30:22]
  reg  valid_16_0; // @[dcache.scala 30:22]
  reg  valid_16_1; // @[dcache.scala 30:22]
  reg  valid_17_0; // @[dcache.scala 30:22]
  reg  valid_17_1; // @[dcache.scala 30:22]
  reg  valid_18_0; // @[dcache.scala 30:22]
  reg  valid_18_1; // @[dcache.scala 30:22]
  reg  valid_19_0; // @[dcache.scala 30:22]
  reg  valid_19_1; // @[dcache.scala 30:22]
  reg  valid_20_0; // @[dcache.scala 30:22]
  reg  valid_20_1; // @[dcache.scala 30:22]
  reg  valid_21_0; // @[dcache.scala 30:22]
  reg  valid_21_1; // @[dcache.scala 30:22]
  reg  valid_22_0; // @[dcache.scala 30:22]
  reg  valid_22_1; // @[dcache.scala 30:22]
  reg  valid_23_0; // @[dcache.scala 30:22]
  reg  valid_23_1; // @[dcache.scala 30:22]
  reg  valid_24_0; // @[dcache.scala 30:22]
  reg  valid_24_1; // @[dcache.scala 30:22]
  reg  valid_25_0; // @[dcache.scala 30:22]
  reg  valid_25_1; // @[dcache.scala 30:22]
  reg  valid_26_0; // @[dcache.scala 30:22]
  reg  valid_26_1; // @[dcache.scala 30:22]
  reg  valid_27_0; // @[dcache.scala 30:22]
  reg  valid_27_1; // @[dcache.scala 30:22]
  reg  valid_28_0; // @[dcache.scala 30:22]
  reg  valid_28_1; // @[dcache.scala 30:22]
  reg  valid_29_0; // @[dcache.scala 30:22]
  reg  valid_29_1; // @[dcache.scala 30:22]
  reg  valid_30_0; // @[dcache.scala 30:22]
  reg  valid_30_1; // @[dcache.scala 30:22]
  reg  valid_31_0; // @[dcache.scala 30:22]
  reg  valid_31_1; // @[dcache.scala 30:22]
  reg  valid_32_0; // @[dcache.scala 30:22]
  reg  valid_32_1; // @[dcache.scala 30:22]
  reg  valid_33_0; // @[dcache.scala 30:22]
  reg  valid_33_1; // @[dcache.scala 30:22]
  reg  valid_34_0; // @[dcache.scala 30:22]
  reg  valid_34_1; // @[dcache.scala 30:22]
  reg  valid_35_0; // @[dcache.scala 30:22]
  reg  valid_35_1; // @[dcache.scala 30:22]
  reg  valid_36_0; // @[dcache.scala 30:22]
  reg  valid_36_1; // @[dcache.scala 30:22]
  reg  valid_37_0; // @[dcache.scala 30:22]
  reg  valid_37_1; // @[dcache.scala 30:22]
  reg  valid_38_0; // @[dcache.scala 30:22]
  reg  valid_38_1; // @[dcache.scala 30:22]
  reg  valid_39_0; // @[dcache.scala 30:22]
  reg  valid_39_1; // @[dcache.scala 30:22]
  reg  valid_40_0; // @[dcache.scala 30:22]
  reg  valid_40_1; // @[dcache.scala 30:22]
  reg  valid_41_0; // @[dcache.scala 30:22]
  reg  valid_41_1; // @[dcache.scala 30:22]
  reg  valid_42_0; // @[dcache.scala 30:22]
  reg  valid_42_1; // @[dcache.scala 30:22]
  reg  valid_43_0; // @[dcache.scala 30:22]
  reg  valid_43_1; // @[dcache.scala 30:22]
  reg  valid_44_0; // @[dcache.scala 30:22]
  reg  valid_44_1; // @[dcache.scala 30:22]
  reg  valid_45_0; // @[dcache.scala 30:22]
  reg  valid_45_1; // @[dcache.scala 30:22]
  reg  valid_46_0; // @[dcache.scala 30:22]
  reg  valid_46_1; // @[dcache.scala 30:22]
  reg  valid_47_0; // @[dcache.scala 30:22]
  reg  valid_47_1; // @[dcache.scala 30:22]
  reg  valid_48_0; // @[dcache.scala 30:22]
  reg  valid_48_1; // @[dcache.scala 30:22]
  reg  valid_49_0; // @[dcache.scala 30:22]
  reg  valid_49_1; // @[dcache.scala 30:22]
  reg  valid_50_0; // @[dcache.scala 30:22]
  reg  valid_50_1; // @[dcache.scala 30:22]
  reg  valid_51_0; // @[dcache.scala 30:22]
  reg  valid_51_1; // @[dcache.scala 30:22]
  reg  valid_52_0; // @[dcache.scala 30:22]
  reg  valid_52_1; // @[dcache.scala 30:22]
  reg  valid_53_0; // @[dcache.scala 30:22]
  reg  valid_53_1; // @[dcache.scala 30:22]
  reg  valid_54_0; // @[dcache.scala 30:22]
  reg  valid_54_1; // @[dcache.scala 30:22]
  reg  valid_55_0; // @[dcache.scala 30:22]
  reg  valid_55_1; // @[dcache.scala 30:22]
  reg  valid_56_0; // @[dcache.scala 30:22]
  reg  valid_56_1; // @[dcache.scala 30:22]
  reg  valid_57_0; // @[dcache.scala 30:22]
  reg  valid_57_1; // @[dcache.scala 30:22]
  reg  valid_58_0; // @[dcache.scala 30:22]
  reg  valid_58_1; // @[dcache.scala 30:22]
  reg  valid_59_0; // @[dcache.scala 30:22]
  reg  valid_59_1; // @[dcache.scala 30:22]
  reg  valid_60_0; // @[dcache.scala 30:22]
  reg  valid_60_1; // @[dcache.scala 30:22]
  reg  valid_61_0; // @[dcache.scala 30:22]
  reg  valid_61_1; // @[dcache.scala 30:22]
  reg  valid_62_0; // @[dcache.scala 30:22]
  reg  valid_62_1; // @[dcache.scala 30:22]
  reg  valid_63_0; // @[dcache.scala 30:22]
  reg  valid_63_1; // @[dcache.scala 30:22]
  reg  valid_64_0; // @[dcache.scala 30:22]
  reg  valid_64_1; // @[dcache.scala 30:22]
  reg  valid_65_0; // @[dcache.scala 30:22]
  reg  valid_65_1; // @[dcache.scala 30:22]
  reg  valid_66_0; // @[dcache.scala 30:22]
  reg  valid_66_1; // @[dcache.scala 30:22]
  reg  valid_67_0; // @[dcache.scala 30:22]
  reg  valid_67_1; // @[dcache.scala 30:22]
  reg  valid_68_0; // @[dcache.scala 30:22]
  reg  valid_68_1; // @[dcache.scala 30:22]
  reg  valid_69_0; // @[dcache.scala 30:22]
  reg  valid_69_1; // @[dcache.scala 30:22]
  reg  valid_70_0; // @[dcache.scala 30:22]
  reg  valid_70_1; // @[dcache.scala 30:22]
  reg  valid_71_0; // @[dcache.scala 30:22]
  reg  valid_71_1; // @[dcache.scala 30:22]
  reg  valid_72_0; // @[dcache.scala 30:22]
  reg  valid_72_1; // @[dcache.scala 30:22]
  reg  valid_73_0; // @[dcache.scala 30:22]
  reg  valid_73_1; // @[dcache.scala 30:22]
  reg  valid_74_0; // @[dcache.scala 30:22]
  reg  valid_74_1; // @[dcache.scala 30:22]
  reg  valid_75_0; // @[dcache.scala 30:22]
  reg  valid_75_1; // @[dcache.scala 30:22]
  reg  valid_76_0; // @[dcache.scala 30:22]
  reg  valid_76_1; // @[dcache.scala 30:22]
  reg  valid_77_0; // @[dcache.scala 30:22]
  reg  valid_77_1; // @[dcache.scala 30:22]
  reg  valid_78_0; // @[dcache.scala 30:22]
  reg  valid_78_1; // @[dcache.scala 30:22]
  reg  valid_79_0; // @[dcache.scala 30:22]
  reg  valid_79_1; // @[dcache.scala 30:22]
  reg  valid_80_0; // @[dcache.scala 30:22]
  reg  valid_80_1; // @[dcache.scala 30:22]
  reg  valid_81_0; // @[dcache.scala 30:22]
  reg  valid_81_1; // @[dcache.scala 30:22]
  reg  valid_82_0; // @[dcache.scala 30:22]
  reg  valid_82_1; // @[dcache.scala 30:22]
  reg  valid_83_0; // @[dcache.scala 30:22]
  reg  valid_83_1; // @[dcache.scala 30:22]
  reg  valid_84_0; // @[dcache.scala 30:22]
  reg  valid_84_1; // @[dcache.scala 30:22]
  reg  valid_85_0; // @[dcache.scala 30:22]
  reg  valid_85_1; // @[dcache.scala 30:22]
  reg  valid_86_0; // @[dcache.scala 30:22]
  reg  valid_86_1; // @[dcache.scala 30:22]
  reg  valid_87_0; // @[dcache.scala 30:22]
  reg  valid_87_1; // @[dcache.scala 30:22]
  reg  valid_88_0; // @[dcache.scala 30:22]
  reg  valid_88_1; // @[dcache.scala 30:22]
  reg  valid_89_0; // @[dcache.scala 30:22]
  reg  valid_89_1; // @[dcache.scala 30:22]
  reg  valid_90_0; // @[dcache.scala 30:22]
  reg  valid_90_1; // @[dcache.scala 30:22]
  reg  valid_91_0; // @[dcache.scala 30:22]
  reg  valid_91_1; // @[dcache.scala 30:22]
  reg  valid_92_0; // @[dcache.scala 30:22]
  reg  valid_92_1; // @[dcache.scala 30:22]
  reg  valid_93_0; // @[dcache.scala 30:22]
  reg  valid_93_1; // @[dcache.scala 30:22]
  reg  valid_94_0; // @[dcache.scala 30:22]
  reg  valid_94_1; // @[dcache.scala 30:22]
  reg  valid_95_0; // @[dcache.scala 30:22]
  reg  valid_95_1; // @[dcache.scala 30:22]
  reg  valid_96_0; // @[dcache.scala 30:22]
  reg  valid_96_1; // @[dcache.scala 30:22]
  reg  valid_97_0; // @[dcache.scala 30:22]
  reg  valid_97_1; // @[dcache.scala 30:22]
  reg  valid_98_0; // @[dcache.scala 30:22]
  reg  valid_98_1; // @[dcache.scala 30:22]
  reg  valid_99_0; // @[dcache.scala 30:22]
  reg  valid_99_1; // @[dcache.scala 30:22]
  reg  valid_100_0; // @[dcache.scala 30:22]
  reg  valid_100_1; // @[dcache.scala 30:22]
  reg  valid_101_0; // @[dcache.scala 30:22]
  reg  valid_101_1; // @[dcache.scala 30:22]
  reg  valid_102_0; // @[dcache.scala 30:22]
  reg  valid_102_1; // @[dcache.scala 30:22]
  reg  valid_103_0; // @[dcache.scala 30:22]
  reg  valid_103_1; // @[dcache.scala 30:22]
  reg  valid_104_0; // @[dcache.scala 30:22]
  reg  valid_104_1; // @[dcache.scala 30:22]
  reg  valid_105_0; // @[dcache.scala 30:22]
  reg  valid_105_1; // @[dcache.scala 30:22]
  reg  valid_106_0; // @[dcache.scala 30:22]
  reg  valid_106_1; // @[dcache.scala 30:22]
  reg  valid_107_0; // @[dcache.scala 30:22]
  reg  valid_107_1; // @[dcache.scala 30:22]
  reg  valid_108_0; // @[dcache.scala 30:22]
  reg  valid_108_1; // @[dcache.scala 30:22]
  reg  valid_109_0; // @[dcache.scala 30:22]
  reg  valid_109_1; // @[dcache.scala 30:22]
  reg  valid_110_0; // @[dcache.scala 30:22]
  reg  valid_110_1; // @[dcache.scala 30:22]
  reg  valid_111_0; // @[dcache.scala 30:22]
  reg  valid_111_1; // @[dcache.scala 30:22]
  reg  valid_112_0; // @[dcache.scala 30:22]
  reg  valid_112_1; // @[dcache.scala 30:22]
  reg  valid_113_0; // @[dcache.scala 30:22]
  reg  valid_113_1; // @[dcache.scala 30:22]
  reg  valid_114_0; // @[dcache.scala 30:22]
  reg  valid_114_1; // @[dcache.scala 30:22]
  reg  valid_115_0; // @[dcache.scala 30:22]
  reg  valid_115_1; // @[dcache.scala 30:22]
  reg  valid_116_0; // @[dcache.scala 30:22]
  reg  valid_116_1; // @[dcache.scala 30:22]
  reg  valid_117_0; // @[dcache.scala 30:22]
  reg  valid_117_1; // @[dcache.scala 30:22]
  reg  valid_118_0; // @[dcache.scala 30:22]
  reg  valid_118_1; // @[dcache.scala 30:22]
  reg  valid_119_0; // @[dcache.scala 30:22]
  reg  valid_119_1; // @[dcache.scala 30:22]
  reg  valid_120_0; // @[dcache.scala 30:22]
  reg  valid_120_1; // @[dcache.scala 30:22]
  reg  valid_121_0; // @[dcache.scala 30:22]
  reg  valid_121_1; // @[dcache.scala 30:22]
  reg  valid_122_0; // @[dcache.scala 30:22]
  reg  valid_122_1; // @[dcache.scala 30:22]
  reg  valid_123_0; // @[dcache.scala 30:22]
  reg  valid_123_1; // @[dcache.scala 30:22]
  reg  valid_124_0; // @[dcache.scala 30:22]
  reg  valid_124_1; // @[dcache.scala 30:22]
  reg  valid_125_0; // @[dcache.scala 30:22]
  reg  valid_125_1; // @[dcache.scala 30:22]
  reg  valid_126_0; // @[dcache.scala 30:22]
  reg  valid_126_1; // @[dcache.scala 30:22]
  reg  valid_127_0; // @[dcache.scala 30:22]
  reg  valid_127_1; // @[dcache.scala 30:22]
  reg  dirty_0_0; // @[dcache.scala 31:22]
  reg  dirty_0_1; // @[dcache.scala 31:22]
  reg  dirty_1_0; // @[dcache.scala 31:22]
  reg  dirty_1_1; // @[dcache.scala 31:22]
  reg  dirty_2_0; // @[dcache.scala 31:22]
  reg  dirty_2_1; // @[dcache.scala 31:22]
  reg  dirty_3_0; // @[dcache.scala 31:22]
  reg  dirty_3_1; // @[dcache.scala 31:22]
  reg  dirty_4_0; // @[dcache.scala 31:22]
  reg  dirty_4_1; // @[dcache.scala 31:22]
  reg  dirty_5_0; // @[dcache.scala 31:22]
  reg  dirty_5_1; // @[dcache.scala 31:22]
  reg  dirty_6_0; // @[dcache.scala 31:22]
  reg  dirty_6_1; // @[dcache.scala 31:22]
  reg  dirty_7_0; // @[dcache.scala 31:22]
  reg  dirty_7_1; // @[dcache.scala 31:22]
  reg  dirty_8_0; // @[dcache.scala 31:22]
  reg  dirty_8_1; // @[dcache.scala 31:22]
  reg  dirty_9_0; // @[dcache.scala 31:22]
  reg  dirty_9_1; // @[dcache.scala 31:22]
  reg  dirty_10_0; // @[dcache.scala 31:22]
  reg  dirty_10_1; // @[dcache.scala 31:22]
  reg  dirty_11_0; // @[dcache.scala 31:22]
  reg  dirty_11_1; // @[dcache.scala 31:22]
  reg  dirty_12_0; // @[dcache.scala 31:22]
  reg  dirty_12_1; // @[dcache.scala 31:22]
  reg  dirty_13_0; // @[dcache.scala 31:22]
  reg  dirty_13_1; // @[dcache.scala 31:22]
  reg  dirty_14_0; // @[dcache.scala 31:22]
  reg  dirty_14_1; // @[dcache.scala 31:22]
  reg  dirty_15_0; // @[dcache.scala 31:22]
  reg  dirty_15_1; // @[dcache.scala 31:22]
  reg  dirty_16_0; // @[dcache.scala 31:22]
  reg  dirty_16_1; // @[dcache.scala 31:22]
  reg  dirty_17_0; // @[dcache.scala 31:22]
  reg  dirty_17_1; // @[dcache.scala 31:22]
  reg  dirty_18_0; // @[dcache.scala 31:22]
  reg  dirty_18_1; // @[dcache.scala 31:22]
  reg  dirty_19_0; // @[dcache.scala 31:22]
  reg  dirty_19_1; // @[dcache.scala 31:22]
  reg  dirty_20_0; // @[dcache.scala 31:22]
  reg  dirty_20_1; // @[dcache.scala 31:22]
  reg  dirty_21_0; // @[dcache.scala 31:22]
  reg  dirty_21_1; // @[dcache.scala 31:22]
  reg  dirty_22_0; // @[dcache.scala 31:22]
  reg  dirty_22_1; // @[dcache.scala 31:22]
  reg  dirty_23_0; // @[dcache.scala 31:22]
  reg  dirty_23_1; // @[dcache.scala 31:22]
  reg  dirty_24_0; // @[dcache.scala 31:22]
  reg  dirty_24_1; // @[dcache.scala 31:22]
  reg  dirty_25_0; // @[dcache.scala 31:22]
  reg  dirty_25_1; // @[dcache.scala 31:22]
  reg  dirty_26_0; // @[dcache.scala 31:22]
  reg  dirty_26_1; // @[dcache.scala 31:22]
  reg  dirty_27_0; // @[dcache.scala 31:22]
  reg  dirty_27_1; // @[dcache.scala 31:22]
  reg  dirty_28_0; // @[dcache.scala 31:22]
  reg  dirty_28_1; // @[dcache.scala 31:22]
  reg  dirty_29_0; // @[dcache.scala 31:22]
  reg  dirty_29_1; // @[dcache.scala 31:22]
  reg  dirty_30_0; // @[dcache.scala 31:22]
  reg  dirty_30_1; // @[dcache.scala 31:22]
  reg  dirty_31_0; // @[dcache.scala 31:22]
  reg  dirty_31_1; // @[dcache.scala 31:22]
  reg  dirty_32_0; // @[dcache.scala 31:22]
  reg  dirty_32_1; // @[dcache.scala 31:22]
  reg  dirty_33_0; // @[dcache.scala 31:22]
  reg  dirty_33_1; // @[dcache.scala 31:22]
  reg  dirty_34_0; // @[dcache.scala 31:22]
  reg  dirty_34_1; // @[dcache.scala 31:22]
  reg  dirty_35_0; // @[dcache.scala 31:22]
  reg  dirty_35_1; // @[dcache.scala 31:22]
  reg  dirty_36_0; // @[dcache.scala 31:22]
  reg  dirty_36_1; // @[dcache.scala 31:22]
  reg  dirty_37_0; // @[dcache.scala 31:22]
  reg  dirty_37_1; // @[dcache.scala 31:22]
  reg  dirty_38_0; // @[dcache.scala 31:22]
  reg  dirty_38_1; // @[dcache.scala 31:22]
  reg  dirty_39_0; // @[dcache.scala 31:22]
  reg  dirty_39_1; // @[dcache.scala 31:22]
  reg  dirty_40_0; // @[dcache.scala 31:22]
  reg  dirty_40_1; // @[dcache.scala 31:22]
  reg  dirty_41_0; // @[dcache.scala 31:22]
  reg  dirty_41_1; // @[dcache.scala 31:22]
  reg  dirty_42_0; // @[dcache.scala 31:22]
  reg  dirty_42_1; // @[dcache.scala 31:22]
  reg  dirty_43_0; // @[dcache.scala 31:22]
  reg  dirty_43_1; // @[dcache.scala 31:22]
  reg  dirty_44_0; // @[dcache.scala 31:22]
  reg  dirty_44_1; // @[dcache.scala 31:22]
  reg  dirty_45_0; // @[dcache.scala 31:22]
  reg  dirty_45_1; // @[dcache.scala 31:22]
  reg  dirty_46_0; // @[dcache.scala 31:22]
  reg  dirty_46_1; // @[dcache.scala 31:22]
  reg  dirty_47_0; // @[dcache.scala 31:22]
  reg  dirty_47_1; // @[dcache.scala 31:22]
  reg  dirty_48_0; // @[dcache.scala 31:22]
  reg  dirty_48_1; // @[dcache.scala 31:22]
  reg  dirty_49_0; // @[dcache.scala 31:22]
  reg  dirty_49_1; // @[dcache.scala 31:22]
  reg  dirty_50_0; // @[dcache.scala 31:22]
  reg  dirty_50_1; // @[dcache.scala 31:22]
  reg  dirty_51_0; // @[dcache.scala 31:22]
  reg  dirty_51_1; // @[dcache.scala 31:22]
  reg  dirty_52_0; // @[dcache.scala 31:22]
  reg  dirty_52_1; // @[dcache.scala 31:22]
  reg  dirty_53_0; // @[dcache.scala 31:22]
  reg  dirty_53_1; // @[dcache.scala 31:22]
  reg  dirty_54_0; // @[dcache.scala 31:22]
  reg  dirty_54_1; // @[dcache.scala 31:22]
  reg  dirty_55_0; // @[dcache.scala 31:22]
  reg  dirty_55_1; // @[dcache.scala 31:22]
  reg  dirty_56_0; // @[dcache.scala 31:22]
  reg  dirty_56_1; // @[dcache.scala 31:22]
  reg  dirty_57_0; // @[dcache.scala 31:22]
  reg  dirty_57_1; // @[dcache.scala 31:22]
  reg  dirty_58_0; // @[dcache.scala 31:22]
  reg  dirty_58_1; // @[dcache.scala 31:22]
  reg  dirty_59_0; // @[dcache.scala 31:22]
  reg  dirty_59_1; // @[dcache.scala 31:22]
  reg  dirty_60_0; // @[dcache.scala 31:22]
  reg  dirty_60_1; // @[dcache.scala 31:22]
  reg  dirty_61_0; // @[dcache.scala 31:22]
  reg  dirty_61_1; // @[dcache.scala 31:22]
  reg  dirty_62_0; // @[dcache.scala 31:22]
  reg  dirty_62_1; // @[dcache.scala 31:22]
  reg  dirty_63_0; // @[dcache.scala 31:22]
  reg  dirty_63_1; // @[dcache.scala 31:22]
  reg  dirty_64_0; // @[dcache.scala 31:22]
  reg  dirty_64_1; // @[dcache.scala 31:22]
  reg  dirty_65_0; // @[dcache.scala 31:22]
  reg  dirty_65_1; // @[dcache.scala 31:22]
  reg  dirty_66_0; // @[dcache.scala 31:22]
  reg  dirty_66_1; // @[dcache.scala 31:22]
  reg  dirty_67_0; // @[dcache.scala 31:22]
  reg  dirty_67_1; // @[dcache.scala 31:22]
  reg  dirty_68_0; // @[dcache.scala 31:22]
  reg  dirty_68_1; // @[dcache.scala 31:22]
  reg  dirty_69_0; // @[dcache.scala 31:22]
  reg  dirty_69_1; // @[dcache.scala 31:22]
  reg  dirty_70_0; // @[dcache.scala 31:22]
  reg  dirty_70_1; // @[dcache.scala 31:22]
  reg  dirty_71_0; // @[dcache.scala 31:22]
  reg  dirty_71_1; // @[dcache.scala 31:22]
  reg  dirty_72_0; // @[dcache.scala 31:22]
  reg  dirty_72_1; // @[dcache.scala 31:22]
  reg  dirty_73_0; // @[dcache.scala 31:22]
  reg  dirty_73_1; // @[dcache.scala 31:22]
  reg  dirty_74_0; // @[dcache.scala 31:22]
  reg  dirty_74_1; // @[dcache.scala 31:22]
  reg  dirty_75_0; // @[dcache.scala 31:22]
  reg  dirty_75_1; // @[dcache.scala 31:22]
  reg  dirty_76_0; // @[dcache.scala 31:22]
  reg  dirty_76_1; // @[dcache.scala 31:22]
  reg  dirty_77_0; // @[dcache.scala 31:22]
  reg  dirty_77_1; // @[dcache.scala 31:22]
  reg  dirty_78_0; // @[dcache.scala 31:22]
  reg  dirty_78_1; // @[dcache.scala 31:22]
  reg  dirty_79_0; // @[dcache.scala 31:22]
  reg  dirty_79_1; // @[dcache.scala 31:22]
  reg  dirty_80_0; // @[dcache.scala 31:22]
  reg  dirty_80_1; // @[dcache.scala 31:22]
  reg  dirty_81_0; // @[dcache.scala 31:22]
  reg  dirty_81_1; // @[dcache.scala 31:22]
  reg  dirty_82_0; // @[dcache.scala 31:22]
  reg  dirty_82_1; // @[dcache.scala 31:22]
  reg  dirty_83_0; // @[dcache.scala 31:22]
  reg  dirty_83_1; // @[dcache.scala 31:22]
  reg  dirty_84_0; // @[dcache.scala 31:22]
  reg  dirty_84_1; // @[dcache.scala 31:22]
  reg  dirty_85_0; // @[dcache.scala 31:22]
  reg  dirty_85_1; // @[dcache.scala 31:22]
  reg  dirty_86_0; // @[dcache.scala 31:22]
  reg  dirty_86_1; // @[dcache.scala 31:22]
  reg  dirty_87_0; // @[dcache.scala 31:22]
  reg  dirty_87_1; // @[dcache.scala 31:22]
  reg  dirty_88_0; // @[dcache.scala 31:22]
  reg  dirty_88_1; // @[dcache.scala 31:22]
  reg  dirty_89_0; // @[dcache.scala 31:22]
  reg  dirty_89_1; // @[dcache.scala 31:22]
  reg  dirty_90_0; // @[dcache.scala 31:22]
  reg  dirty_90_1; // @[dcache.scala 31:22]
  reg  dirty_91_0; // @[dcache.scala 31:22]
  reg  dirty_91_1; // @[dcache.scala 31:22]
  reg  dirty_92_0; // @[dcache.scala 31:22]
  reg  dirty_92_1; // @[dcache.scala 31:22]
  reg  dirty_93_0; // @[dcache.scala 31:22]
  reg  dirty_93_1; // @[dcache.scala 31:22]
  reg  dirty_94_0; // @[dcache.scala 31:22]
  reg  dirty_94_1; // @[dcache.scala 31:22]
  reg  dirty_95_0; // @[dcache.scala 31:22]
  reg  dirty_95_1; // @[dcache.scala 31:22]
  reg  dirty_96_0; // @[dcache.scala 31:22]
  reg  dirty_96_1; // @[dcache.scala 31:22]
  reg  dirty_97_0; // @[dcache.scala 31:22]
  reg  dirty_97_1; // @[dcache.scala 31:22]
  reg  dirty_98_0; // @[dcache.scala 31:22]
  reg  dirty_98_1; // @[dcache.scala 31:22]
  reg  dirty_99_0; // @[dcache.scala 31:22]
  reg  dirty_99_1; // @[dcache.scala 31:22]
  reg  dirty_100_0; // @[dcache.scala 31:22]
  reg  dirty_100_1; // @[dcache.scala 31:22]
  reg  dirty_101_0; // @[dcache.scala 31:22]
  reg  dirty_101_1; // @[dcache.scala 31:22]
  reg  dirty_102_0; // @[dcache.scala 31:22]
  reg  dirty_102_1; // @[dcache.scala 31:22]
  reg  dirty_103_0; // @[dcache.scala 31:22]
  reg  dirty_103_1; // @[dcache.scala 31:22]
  reg  dirty_104_0; // @[dcache.scala 31:22]
  reg  dirty_104_1; // @[dcache.scala 31:22]
  reg  dirty_105_0; // @[dcache.scala 31:22]
  reg  dirty_105_1; // @[dcache.scala 31:22]
  reg  dirty_106_0; // @[dcache.scala 31:22]
  reg  dirty_106_1; // @[dcache.scala 31:22]
  reg  dirty_107_0; // @[dcache.scala 31:22]
  reg  dirty_107_1; // @[dcache.scala 31:22]
  reg  dirty_108_0; // @[dcache.scala 31:22]
  reg  dirty_108_1; // @[dcache.scala 31:22]
  reg  dirty_109_0; // @[dcache.scala 31:22]
  reg  dirty_109_1; // @[dcache.scala 31:22]
  reg  dirty_110_0; // @[dcache.scala 31:22]
  reg  dirty_110_1; // @[dcache.scala 31:22]
  reg  dirty_111_0; // @[dcache.scala 31:22]
  reg  dirty_111_1; // @[dcache.scala 31:22]
  reg  dirty_112_0; // @[dcache.scala 31:22]
  reg  dirty_112_1; // @[dcache.scala 31:22]
  reg  dirty_113_0; // @[dcache.scala 31:22]
  reg  dirty_113_1; // @[dcache.scala 31:22]
  reg  dirty_114_0; // @[dcache.scala 31:22]
  reg  dirty_114_1; // @[dcache.scala 31:22]
  reg  dirty_115_0; // @[dcache.scala 31:22]
  reg  dirty_115_1; // @[dcache.scala 31:22]
  reg  dirty_116_0; // @[dcache.scala 31:22]
  reg  dirty_116_1; // @[dcache.scala 31:22]
  reg  dirty_117_0; // @[dcache.scala 31:22]
  reg  dirty_117_1; // @[dcache.scala 31:22]
  reg  dirty_118_0; // @[dcache.scala 31:22]
  reg  dirty_118_1; // @[dcache.scala 31:22]
  reg  dirty_119_0; // @[dcache.scala 31:22]
  reg  dirty_119_1; // @[dcache.scala 31:22]
  reg  dirty_120_0; // @[dcache.scala 31:22]
  reg  dirty_120_1; // @[dcache.scala 31:22]
  reg  dirty_121_0; // @[dcache.scala 31:22]
  reg  dirty_121_1; // @[dcache.scala 31:22]
  reg  dirty_122_0; // @[dcache.scala 31:22]
  reg  dirty_122_1; // @[dcache.scala 31:22]
  reg  dirty_123_0; // @[dcache.scala 31:22]
  reg  dirty_123_1; // @[dcache.scala 31:22]
  reg  dirty_124_0; // @[dcache.scala 31:22]
  reg  dirty_124_1; // @[dcache.scala 31:22]
  reg  dirty_125_0; // @[dcache.scala 31:22]
  reg  dirty_125_1; // @[dcache.scala 31:22]
  reg  dirty_126_0; // @[dcache.scala 31:22]
  reg  dirty_126_1; // @[dcache.scala 31:22]
  reg  dirty_127_0; // @[dcache.scala 31:22]
  reg  dirty_127_1; // @[dcache.scala 31:22]
  reg [127:0] buf_; // @[dcache.scala 32:20]
  reg [2:0] state; // @[dcache.scala 36:22]
  reg [2:0] rstate; // @[dcache.scala 37:23]
  reg [2:0] wstate; // @[dcache.scala 38:23]
  wire  _req_T = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 52:35]
  wire  _req_T_1 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 52:35]
  wire  req = _req_T | _req_T_1; // @[dcache.scala 39:28]
  reg [31:0] addr; // @[dcache.scala 41:21]
  reg [63:0] wdata; // @[dcache.scala 42:22]
  reg [7:0] wstrb; // @[dcache.scala 43:22]
  reg  uncache; // @[dcache.scala 44:24]
  wire [20:0] tag = addr[31:11]; // @[dcache.scala 45:17]
  wire [6:0] offset = {addr[3:0], 3'h0}; // @[dcache.scala 46:42]
  wire [6:0] idx = addr[10:4]; // @[dcache.scala 47:17]
  reg  rmode; // @[dcache.scala 55:22]
  reg  wmode; // @[dcache.scala 56:22]
  wire  _rmode_T = state == 3'h0; // @[dcache.scala 57:23]
  wire  _rmode_T_2 = state == 3'h0 & _req_T; // @[dcache.scala 57:35]
  wire  _rmode_T_4 = state == 3'h0 ? 1'h0 : rmode; // @[dcache.scala 57:58]
  wire  _wmode_T_2 = _rmode_T & _req_T_1; // @[dcache.scala 58:35]
  wire  _wmode_T_4 = _rmode_T ? 1'h0 : wmode; // @[dcache.scala 58:58]
  wire [41:0] _GEN_1 = 7'h1 == idx ? cache_tag_1 : cache_tag_0; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_2 = 7'h2 == idx ? cache_tag_2 : _GEN_1; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_3 = 7'h3 == idx ? cache_tag_3 : _GEN_2; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_4 = 7'h4 == idx ? cache_tag_4 : _GEN_3; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_5 = 7'h5 == idx ? cache_tag_5 : _GEN_4; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_6 = 7'h6 == idx ? cache_tag_6 : _GEN_5; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_7 = 7'h7 == idx ? cache_tag_7 : _GEN_6; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_8 = 7'h8 == idx ? cache_tag_8 : _GEN_7; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_9 = 7'h9 == idx ? cache_tag_9 : _GEN_8; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_10 = 7'ha == idx ? cache_tag_10 : _GEN_9; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_11 = 7'hb == idx ? cache_tag_11 : _GEN_10; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_12 = 7'hc == idx ? cache_tag_12 : _GEN_11; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_13 = 7'hd == idx ? cache_tag_13 : _GEN_12; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_14 = 7'he == idx ? cache_tag_14 : _GEN_13; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_15 = 7'hf == idx ? cache_tag_15 : _GEN_14; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_16 = 7'h10 == idx ? cache_tag_16 : _GEN_15; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_17 = 7'h11 == idx ? cache_tag_17 : _GEN_16; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_18 = 7'h12 == idx ? cache_tag_18 : _GEN_17; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_19 = 7'h13 == idx ? cache_tag_19 : _GEN_18; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_20 = 7'h14 == idx ? cache_tag_20 : _GEN_19; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_21 = 7'h15 == idx ? cache_tag_21 : _GEN_20; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_22 = 7'h16 == idx ? cache_tag_22 : _GEN_21; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_23 = 7'h17 == idx ? cache_tag_23 : _GEN_22; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_24 = 7'h18 == idx ? cache_tag_24 : _GEN_23; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_25 = 7'h19 == idx ? cache_tag_25 : _GEN_24; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_26 = 7'h1a == idx ? cache_tag_26 : _GEN_25; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_27 = 7'h1b == idx ? cache_tag_27 : _GEN_26; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_28 = 7'h1c == idx ? cache_tag_28 : _GEN_27; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_29 = 7'h1d == idx ? cache_tag_29 : _GEN_28; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_30 = 7'h1e == idx ? cache_tag_30 : _GEN_29; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_31 = 7'h1f == idx ? cache_tag_31 : _GEN_30; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_32 = 7'h20 == idx ? cache_tag_32 : _GEN_31; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_33 = 7'h21 == idx ? cache_tag_33 : _GEN_32; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_34 = 7'h22 == idx ? cache_tag_34 : _GEN_33; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_35 = 7'h23 == idx ? cache_tag_35 : _GEN_34; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_36 = 7'h24 == idx ? cache_tag_36 : _GEN_35; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_37 = 7'h25 == idx ? cache_tag_37 : _GEN_36; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_38 = 7'h26 == idx ? cache_tag_38 : _GEN_37; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_39 = 7'h27 == idx ? cache_tag_39 : _GEN_38; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_40 = 7'h28 == idx ? cache_tag_40 : _GEN_39; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_41 = 7'h29 == idx ? cache_tag_41 : _GEN_40; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_42 = 7'h2a == idx ? cache_tag_42 : _GEN_41; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_43 = 7'h2b == idx ? cache_tag_43 : _GEN_42; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_44 = 7'h2c == idx ? cache_tag_44 : _GEN_43; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_45 = 7'h2d == idx ? cache_tag_45 : _GEN_44; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_46 = 7'h2e == idx ? cache_tag_46 : _GEN_45; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_47 = 7'h2f == idx ? cache_tag_47 : _GEN_46; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_48 = 7'h30 == idx ? cache_tag_48 : _GEN_47; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_49 = 7'h31 == idx ? cache_tag_49 : _GEN_48; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_50 = 7'h32 == idx ? cache_tag_50 : _GEN_49; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_51 = 7'h33 == idx ? cache_tag_51 : _GEN_50; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_52 = 7'h34 == idx ? cache_tag_52 : _GEN_51; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_53 = 7'h35 == idx ? cache_tag_53 : _GEN_52; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_54 = 7'h36 == idx ? cache_tag_54 : _GEN_53; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_55 = 7'h37 == idx ? cache_tag_55 : _GEN_54; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_56 = 7'h38 == idx ? cache_tag_56 : _GEN_55; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_57 = 7'h39 == idx ? cache_tag_57 : _GEN_56; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_58 = 7'h3a == idx ? cache_tag_58 : _GEN_57; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_59 = 7'h3b == idx ? cache_tag_59 : _GEN_58; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_60 = 7'h3c == idx ? cache_tag_60 : _GEN_59; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_61 = 7'h3d == idx ? cache_tag_61 : _GEN_60; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_62 = 7'h3e == idx ? cache_tag_62 : _GEN_61; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_63 = 7'h3f == idx ? cache_tag_63 : _GEN_62; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_64 = 7'h40 == idx ? cache_tag_64 : _GEN_63; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_65 = 7'h41 == idx ? cache_tag_65 : _GEN_64; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_66 = 7'h42 == idx ? cache_tag_66 : _GEN_65; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_67 = 7'h43 == idx ? cache_tag_67 : _GEN_66; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_68 = 7'h44 == idx ? cache_tag_68 : _GEN_67; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_69 = 7'h45 == idx ? cache_tag_69 : _GEN_68; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_70 = 7'h46 == idx ? cache_tag_70 : _GEN_69; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_71 = 7'h47 == idx ? cache_tag_71 : _GEN_70; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_72 = 7'h48 == idx ? cache_tag_72 : _GEN_71; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_73 = 7'h49 == idx ? cache_tag_73 : _GEN_72; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_74 = 7'h4a == idx ? cache_tag_74 : _GEN_73; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_75 = 7'h4b == idx ? cache_tag_75 : _GEN_74; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_76 = 7'h4c == idx ? cache_tag_76 : _GEN_75; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_77 = 7'h4d == idx ? cache_tag_77 : _GEN_76; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_78 = 7'h4e == idx ? cache_tag_78 : _GEN_77; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_79 = 7'h4f == idx ? cache_tag_79 : _GEN_78; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_80 = 7'h50 == idx ? cache_tag_80 : _GEN_79; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_81 = 7'h51 == idx ? cache_tag_81 : _GEN_80; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_82 = 7'h52 == idx ? cache_tag_82 : _GEN_81; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_83 = 7'h53 == idx ? cache_tag_83 : _GEN_82; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_84 = 7'h54 == idx ? cache_tag_84 : _GEN_83; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_85 = 7'h55 == idx ? cache_tag_85 : _GEN_84; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_86 = 7'h56 == idx ? cache_tag_86 : _GEN_85; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_87 = 7'h57 == idx ? cache_tag_87 : _GEN_86; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_88 = 7'h58 == idx ? cache_tag_88 : _GEN_87; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_89 = 7'h59 == idx ? cache_tag_89 : _GEN_88; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_90 = 7'h5a == idx ? cache_tag_90 : _GEN_89; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_91 = 7'h5b == idx ? cache_tag_91 : _GEN_90; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_92 = 7'h5c == idx ? cache_tag_92 : _GEN_91; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_93 = 7'h5d == idx ? cache_tag_93 : _GEN_92; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_94 = 7'h5e == idx ? cache_tag_94 : _GEN_93; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_95 = 7'h5f == idx ? cache_tag_95 : _GEN_94; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_96 = 7'h60 == idx ? cache_tag_96 : _GEN_95; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_97 = 7'h61 == idx ? cache_tag_97 : _GEN_96; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_98 = 7'h62 == idx ? cache_tag_98 : _GEN_97; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_99 = 7'h63 == idx ? cache_tag_99 : _GEN_98; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_100 = 7'h64 == idx ? cache_tag_100 : _GEN_99; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_101 = 7'h65 == idx ? cache_tag_101 : _GEN_100; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_102 = 7'h66 == idx ? cache_tag_102 : _GEN_101; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_103 = 7'h67 == idx ? cache_tag_103 : _GEN_102; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_104 = 7'h68 == idx ? cache_tag_104 : _GEN_103; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_105 = 7'h69 == idx ? cache_tag_105 : _GEN_104; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_106 = 7'h6a == idx ? cache_tag_106 : _GEN_105; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_107 = 7'h6b == idx ? cache_tag_107 : _GEN_106; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_108 = 7'h6c == idx ? cache_tag_108 : _GEN_107; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_109 = 7'h6d == idx ? cache_tag_109 : _GEN_108; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_110 = 7'h6e == idx ? cache_tag_110 : _GEN_109; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_111 = 7'h6f == idx ? cache_tag_111 : _GEN_110; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_112 = 7'h70 == idx ? cache_tag_112 : _GEN_111; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_113 = 7'h71 == idx ? cache_tag_113 : _GEN_112; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_114 = 7'h72 == idx ? cache_tag_114 : _GEN_113; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_115 = 7'h73 == idx ? cache_tag_115 : _GEN_114; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_116 = 7'h74 == idx ? cache_tag_116 : _GEN_115; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_117 = 7'h75 == idx ? cache_tag_117 : _GEN_116; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_118 = 7'h76 == idx ? cache_tag_118 : _GEN_117; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_119 = 7'h77 == idx ? cache_tag_119 : _GEN_118; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_120 = 7'h78 == idx ? cache_tag_120 : _GEN_119; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_121 = 7'h79 == idx ? cache_tag_121 : _GEN_120; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_122 = 7'h7a == idx ? cache_tag_122 : _GEN_121; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_123 = 7'h7b == idx ? cache_tag_123 : _GEN_122; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_124 = 7'h7c == idx ? cache_tag_124 : _GEN_123; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_125 = 7'h7d == idx ? cache_tag_125 : _GEN_124; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_126 = 7'h7e == idx ? cache_tag_126 : _GEN_125; // @[dcache.scala 61:{33,33}]
  wire [41:0] _GEN_127 = 7'h7f == idx ? cache_tag_127 : _GEN_126; // @[dcache.scala 61:{33,33}]
  wire  _GEN_129 = 7'h1 == idx ? valid_1_0 : valid_0_0; // @[dcache.scala 61:{70,70}]
  wire  _GEN_130 = 7'h2 == idx ? valid_2_0 : _GEN_129; // @[dcache.scala 61:{70,70}]
  wire  _GEN_131 = 7'h3 == idx ? valid_3_0 : _GEN_130; // @[dcache.scala 61:{70,70}]
  wire  _GEN_132 = 7'h4 == idx ? valid_4_0 : _GEN_131; // @[dcache.scala 61:{70,70}]
  wire  _GEN_133 = 7'h5 == idx ? valid_5_0 : _GEN_132; // @[dcache.scala 61:{70,70}]
  wire  _GEN_134 = 7'h6 == idx ? valid_6_0 : _GEN_133; // @[dcache.scala 61:{70,70}]
  wire  _GEN_135 = 7'h7 == idx ? valid_7_0 : _GEN_134; // @[dcache.scala 61:{70,70}]
  wire  _GEN_136 = 7'h8 == idx ? valid_8_0 : _GEN_135; // @[dcache.scala 61:{70,70}]
  wire  _GEN_137 = 7'h9 == idx ? valid_9_0 : _GEN_136; // @[dcache.scala 61:{70,70}]
  wire  _GEN_138 = 7'ha == idx ? valid_10_0 : _GEN_137; // @[dcache.scala 61:{70,70}]
  wire  _GEN_139 = 7'hb == idx ? valid_11_0 : _GEN_138; // @[dcache.scala 61:{70,70}]
  wire  _GEN_140 = 7'hc == idx ? valid_12_0 : _GEN_139; // @[dcache.scala 61:{70,70}]
  wire  _GEN_141 = 7'hd == idx ? valid_13_0 : _GEN_140; // @[dcache.scala 61:{70,70}]
  wire  _GEN_142 = 7'he == idx ? valid_14_0 : _GEN_141; // @[dcache.scala 61:{70,70}]
  wire  _GEN_143 = 7'hf == idx ? valid_15_0 : _GEN_142; // @[dcache.scala 61:{70,70}]
  wire  _GEN_144 = 7'h10 == idx ? valid_16_0 : _GEN_143; // @[dcache.scala 61:{70,70}]
  wire  _GEN_145 = 7'h11 == idx ? valid_17_0 : _GEN_144; // @[dcache.scala 61:{70,70}]
  wire  _GEN_146 = 7'h12 == idx ? valid_18_0 : _GEN_145; // @[dcache.scala 61:{70,70}]
  wire  _GEN_147 = 7'h13 == idx ? valid_19_0 : _GEN_146; // @[dcache.scala 61:{70,70}]
  wire  _GEN_148 = 7'h14 == idx ? valid_20_0 : _GEN_147; // @[dcache.scala 61:{70,70}]
  wire  _GEN_149 = 7'h15 == idx ? valid_21_0 : _GEN_148; // @[dcache.scala 61:{70,70}]
  wire  _GEN_150 = 7'h16 == idx ? valid_22_0 : _GEN_149; // @[dcache.scala 61:{70,70}]
  wire  _GEN_151 = 7'h17 == idx ? valid_23_0 : _GEN_150; // @[dcache.scala 61:{70,70}]
  wire  _GEN_152 = 7'h18 == idx ? valid_24_0 : _GEN_151; // @[dcache.scala 61:{70,70}]
  wire  _GEN_153 = 7'h19 == idx ? valid_25_0 : _GEN_152; // @[dcache.scala 61:{70,70}]
  wire  _GEN_154 = 7'h1a == idx ? valid_26_0 : _GEN_153; // @[dcache.scala 61:{70,70}]
  wire  _GEN_155 = 7'h1b == idx ? valid_27_0 : _GEN_154; // @[dcache.scala 61:{70,70}]
  wire  _GEN_156 = 7'h1c == idx ? valid_28_0 : _GEN_155; // @[dcache.scala 61:{70,70}]
  wire  _GEN_157 = 7'h1d == idx ? valid_29_0 : _GEN_156; // @[dcache.scala 61:{70,70}]
  wire  _GEN_158 = 7'h1e == idx ? valid_30_0 : _GEN_157; // @[dcache.scala 61:{70,70}]
  wire  _GEN_159 = 7'h1f == idx ? valid_31_0 : _GEN_158; // @[dcache.scala 61:{70,70}]
  wire  _GEN_160 = 7'h20 == idx ? valid_32_0 : _GEN_159; // @[dcache.scala 61:{70,70}]
  wire  _GEN_161 = 7'h21 == idx ? valid_33_0 : _GEN_160; // @[dcache.scala 61:{70,70}]
  wire  _GEN_162 = 7'h22 == idx ? valid_34_0 : _GEN_161; // @[dcache.scala 61:{70,70}]
  wire  _GEN_163 = 7'h23 == idx ? valid_35_0 : _GEN_162; // @[dcache.scala 61:{70,70}]
  wire  _GEN_164 = 7'h24 == idx ? valid_36_0 : _GEN_163; // @[dcache.scala 61:{70,70}]
  wire  _GEN_165 = 7'h25 == idx ? valid_37_0 : _GEN_164; // @[dcache.scala 61:{70,70}]
  wire  _GEN_166 = 7'h26 == idx ? valid_38_0 : _GEN_165; // @[dcache.scala 61:{70,70}]
  wire  _GEN_167 = 7'h27 == idx ? valid_39_0 : _GEN_166; // @[dcache.scala 61:{70,70}]
  wire  _GEN_168 = 7'h28 == idx ? valid_40_0 : _GEN_167; // @[dcache.scala 61:{70,70}]
  wire  _GEN_169 = 7'h29 == idx ? valid_41_0 : _GEN_168; // @[dcache.scala 61:{70,70}]
  wire  _GEN_170 = 7'h2a == idx ? valid_42_0 : _GEN_169; // @[dcache.scala 61:{70,70}]
  wire  _GEN_171 = 7'h2b == idx ? valid_43_0 : _GEN_170; // @[dcache.scala 61:{70,70}]
  wire  _GEN_172 = 7'h2c == idx ? valid_44_0 : _GEN_171; // @[dcache.scala 61:{70,70}]
  wire  _GEN_173 = 7'h2d == idx ? valid_45_0 : _GEN_172; // @[dcache.scala 61:{70,70}]
  wire  _GEN_174 = 7'h2e == idx ? valid_46_0 : _GEN_173; // @[dcache.scala 61:{70,70}]
  wire  _GEN_175 = 7'h2f == idx ? valid_47_0 : _GEN_174; // @[dcache.scala 61:{70,70}]
  wire  _GEN_176 = 7'h30 == idx ? valid_48_0 : _GEN_175; // @[dcache.scala 61:{70,70}]
  wire  _GEN_177 = 7'h31 == idx ? valid_49_0 : _GEN_176; // @[dcache.scala 61:{70,70}]
  wire  _GEN_178 = 7'h32 == idx ? valid_50_0 : _GEN_177; // @[dcache.scala 61:{70,70}]
  wire  _GEN_179 = 7'h33 == idx ? valid_51_0 : _GEN_178; // @[dcache.scala 61:{70,70}]
  wire  _GEN_180 = 7'h34 == idx ? valid_52_0 : _GEN_179; // @[dcache.scala 61:{70,70}]
  wire  _GEN_181 = 7'h35 == idx ? valid_53_0 : _GEN_180; // @[dcache.scala 61:{70,70}]
  wire  _GEN_182 = 7'h36 == idx ? valid_54_0 : _GEN_181; // @[dcache.scala 61:{70,70}]
  wire  _GEN_183 = 7'h37 == idx ? valid_55_0 : _GEN_182; // @[dcache.scala 61:{70,70}]
  wire  _GEN_184 = 7'h38 == idx ? valid_56_0 : _GEN_183; // @[dcache.scala 61:{70,70}]
  wire  _GEN_185 = 7'h39 == idx ? valid_57_0 : _GEN_184; // @[dcache.scala 61:{70,70}]
  wire  _GEN_186 = 7'h3a == idx ? valid_58_0 : _GEN_185; // @[dcache.scala 61:{70,70}]
  wire  _GEN_187 = 7'h3b == idx ? valid_59_0 : _GEN_186; // @[dcache.scala 61:{70,70}]
  wire  _GEN_188 = 7'h3c == idx ? valid_60_0 : _GEN_187; // @[dcache.scala 61:{70,70}]
  wire  _GEN_189 = 7'h3d == idx ? valid_61_0 : _GEN_188; // @[dcache.scala 61:{70,70}]
  wire  _GEN_190 = 7'h3e == idx ? valid_62_0 : _GEN_189; // @[dcache.scala 61:{70,70}]
  wire  _GEN_191 = 7'h3f == idx ? valid_63_0 : _GEN_190; // @[dcache.scala 61:{70,70}]
  wire  _GEN_192 = 7'h40 == idx ? valid_64_0 : _GEN_191; // @[dcache.scala 61:{70,70}]
  wire  _GEN_193 = 7'h41 == idx ? valid_65_0 : _GEN_192; // @[dcache.scala 61:{70,70}]
  wire  _GEN_194 = 7'h42 == idx ? valid_66_0 : _GEN_193; // @[dcache.scala 61:{70,70}]
  wire  _GEN_195 = 7'h43 == idx ? valid_67_0 : _GEN_194; // @[dcache.scala 61:{70,70}]
  wire  _GEN_196 = 7'h44 == idx ? valid_68_0 : _GEN_195; // @[dcache.scala 61:{70,70}]
  wire  _GEN_197 = 7'h45 == idx ? valid_69_0 : _GEN_196; // @[dcache.scala 61:{70,70}]
  wire  _GEN_198 = 7'h46 == idx ? valid_70_0 : _GEN_197; // @[dcache.scala 61:{70,70}]
  wire  _GEN_199 = 7'h47 == idx ? valid_71_0 : _GEN_198; // @[dcache.scala 61:{70,70}]
  wire  _GEN_200 = 7'h48 == idx ? valid_72_0 : _GEN_199; // @[dcache.scala 61:{70,70}]
  wire  _GEN_201 = 7'h49 == idx ? valid_73_0 : _GEN_200; // @[dcache.scala 61:{70,70}]
  wire  _GEN_202 = 7'h4a == idx ? valid_74_0 : _GEN_201; // @[dcache.scala 61:{70,70}]
  wire  _GEN_203 = 7'h4b == idx ? valid_75_0 : _GEN_202; // @[dcache.scala 61:{70,70}]
  wire  _GEN_204 = 7'h4c == idx ? valid_76_0 : _GEN_203; // @[dcache.scala 61:{70,70}]
  wire  _GEN_205 = 7'h4d == idx ? valid_77_0 : _GEN_204; // @[dcache.scala 61:{70,70}]
  wire  _GEN_206 = 7'h4e == idx ? valid_78_0 : _GEN_205; // @[dcache.scala 61:{70,70}]
  wire  _GEN_207 = 7'h4f == idx ? valid_79_0 : _GEN_206; // @[dcache.scala 61:{70,70}]
  wire  _GEN_208 = 7'h50 == idx ? valid_80_0 : _GEN_207; // @[dcache.scala 61:{70,70}]
  wire  _GEN_209 = 7'h51 == idx ? valid_81_0 : _GEN_208; // @[dcache.scala 61:{70,70}]
  wire  _GEN_210 = 7'h52 == idx ? valid_82_0 : _GEN_209; // @[dcache.scala 61:{70,70}]
  wire  _GEN_211 = 7'h53 == idx ? valid_83_0 : _GEN_210; // @[dcache.scala 61:{70,70}]
  wire  _GEN_212 = 7'h54 == idx ? valid_84_0 : _GEN_211; // @[dcache.scala 61:{70,70}]
  wire  _GEN_213 = 7'h55 == idx ? valid_85_0 : _GEN_212; // @[dcache.scala 61:{70,70}]
  wire  _GEN_214 = 7'h56 == idx ? valid_86_0 : _GEN_213; // @[dcache.scala 61:{70,70}]
  wire  _GEN_215 = 7'h57 == idx ? valid_87_0 : _GEN_214; // @[dcache.scala 61:{70,70}]
  wire  _GEN_216 = 7'h58 == idx ? valid_88_0 : _GEN_215; // @[dcache.scala 61:{70,70}]
  wire  _GEN_217 = 7'h59 == idx ? valid_89_0 : _GEN_216; // @[dcache.scala 61:{70,70}]
  wire  _GEN_218 = 7'h5a == idx ? valid_90_0 : _GEN_217; // @[dcache.scala 61:{70,70}]
  wire  _GEN_219 = 7'h5b == idx ? valid_91_0 : _GEN_218; // @[dcache.scala 61:{70,70}]
  wire  _GEN_220 = 7'h5c == idx ? valid_92_0 : _GEN_219; // @[dcache.scala 61:{70,70}]
  wire  _GEN_221 = 7'h5d == idx ? valid_93_0 : _GEN_220; // @[dcache.scala 61:{70,70}]
  wire  _GEN_222 = 7'h5e == idx ? valid_94_0 : _GEN_221; // @[dcache.scala 61:{70,70}]
  wire  _GEN_223 = 7'h5f == idx ? valid_95_0 : _GEN_222; // @[dcache.scala 61:{70,70}]
  wire  _GEN_224 = 7'h60 == idx ? valid_96_0 : _GEN_223; // @[dcache.scala 61:{70,70}]
  wire  _GEN_225 = 7'h61 == idx ? valid_97_0 : _GEN_224; // @[dcache.scala 61:{70,70}]
  wire  _GEN_226 = 7'h62 == idx ? valid_98_0 : _GEN_225; // @[dcache.scala 61:{70,70}]
  wire  _GEN_227 = 7'h63 == idx ? valid_99_0 : _GEN_226; // @[dcache.scala 61:{70,70}]
  wire  _GEN_228 = 7'h64 == idx ? valid_100_0 : _GEN_227; // @[dcache.scala 61:{70,70}]
  wire  _GEN_229 = 7'h65 == idx ? valid_101_0 : _GEN_228; // @[dcache.scala 61:{70,70}]
  wire  _GEN_230 = 7'h66 == idx ? valid_102_0 : _GEN_229; // @[dcache.scala 61:{70,70}]
  wire  _GEN_231 = 7'h67 == idx ? valid_103_0 : _GEN_230; // @[dcache.scala 61:{70,70}]
  wire  _GEN_232 = 7'h68 == idx ? valid_104_0 : _GEN_231; // @[dcache.scala 61:{70,70}]
  wire  _GEN_233 = 7'h69 == idx ? valid_105_0 : _GEN_232; // @[dcache.scala 61:{70,70}]
  wire  _GEN_234 = 7'h6a == idx ? valid_106_0 : _GEN_233; // @[dcache.scala 61:{70,70}]
  wire  _GEN_235 = 7'h6b == idx ? valid_107_0 : _GEN_234; // @[dcache.scala 61:{70,70}]
  wire  _GEN_236 = 7'h6c == idx ? valid_108_0 : _GEN_235; // @[dcache.scala 61:{70,70}]
  wire  _GEN_237 = 7'h6d == idx ? valid_109_0 : _GEN_236; // @[dcache.scala 61:{70,70}]
  wire  _GEN_238 = 7'h6e == idx ? valid_110_0 : _GEN_237; // @[dcache.scala 61:{70,70}]
  wire  _GEN_239 = 7'h6f == idx ? valid_111_0 : _GEN_238; // @[dcache.scala 61:{70,70}]
  wire  _GEN_240 = 7'h70 == idx ? valid_112_0 : _GEN_239; // @[dcache.scala 61:{70,70}]
  wire  _GEN_241 = 7'h71 == idx ? valid_113_0 : _GEN_240; // @[dcache.scala 61:{70,70}]
  wire  _GEN_242 = 7'h72 == idx ? valid_114_0 : _GEN_241; // @[dcache.scala 61:{70,70}]
  wire  _GEN_243 = 7'h73 == idx ? valid_115_0 : _GEN_242; // @[dcache.scala 61:{70,70}]
  wire  _GEN_244 = 7'h74 == idx ? valid_116_0 : _GEN_243; // @[dcache.scala 61:{70,70}]
  wire  _GEN_245 = 7'h75 == idx ? valid_117_0 : _GEN_244; // @[dcache.scala 61:{70,70}]
  wire  _GEN_246 = 7'h76 == idx ? valid_118_0 : _GEN_245; // @[dcache.scala 61:{70,70}]
  wire  _GEN_247 = 7'h77 == idx ? valid_119_0 : _GEN_246; // @[dcache.scala 61:{70,70}]
  wire  _GEN_248 = 7'h78 == idx ? valid_120_0 : _GEN_247; // @[dcache.scala 61:{70,70}]
  wire  _GEN_249 = 7'h79 == idx ? valid_121_0 : _GEN_248; // @[dcache.scala 61:{70,70}]
  wire  _GEN_250 = 7'h7a == idx ? valid_122_0 : _GEN_249; // @[dcache.scala 61:{70,70}]
  wire  _GEN_251 = 7'h7b == idx ? valid_123_0 : _GEN_250; // @[dcache.scala 61:{70,70}]
  wire  _GEN_252 = 7'h7c == idx ? valid_124_0 : _GEN_251; // @[dcache.scala 61:{70,70}]
  wire  _GEN_253 = 7'h7d == idx ? valid_125_0 : _GEN_252; // @[dcache.scala 61:{70,70}]
  wire  _GEN_254 = 7'h7e == idx ? valid_126_0 : _GEN_253; // @[dcache.scala 61:{70,70}]
  wire  _GEN_255 = 7'h7f == idx ? valid_127_0 : _GEN_254; // @[dcache.scala 61:{70,70}]
  wire  _GEN_257 = 7'h1 == idx ? valid_1_1 : valid_0_1; // @[dcache.scala 62:{70,70}]
  wire  _GEN_258 = 7'h2 == idx ? valid_2_1 : _GEN_257; // @[dcache.scala 62:{70,70}]
  wire  _GEN_259 = 7'h3 == idx ? valid_3_1 : _GEN_258; // @[dcache.scala 62:{70,70}]
  wire  _GEN_260 = 7'h4 == idx ? valid_4_1 : _GEN_259; // @[dcache.scala 62:{70,70}]
  wire  _GEN_261 = 7'h5 == idx ? valid_5_1 : _GEN_260; // @[dcache.scala 62:{70,70}]
  wire  _GEN_262 = 7'h6 == idx ? valid_6_1 : _GEN_261; // @[dcache.scala 62:{70,70}]
  wire  _GEN_263 = 7'h7 == idx ? valid_7_1 : _GEN_262; // @[dcache.scala 62:{70,70}]
  wire  _GEN_264 = 7'h8 == idx ? valid_8_1 : _GEN_263; // @[dcache.scala 62:{70,70}]
  wire  _GEN_265 = 7'h9 == idx ? valid_9_1 : _GEN_264; // @[dcache.scala 62:{70,70}]
  wire  _GEN_266 = 7'ha == idx ? valid_10_1 : _GEN_265; // @[dcache.scala 62:{70,70}]
  wire  _GEN_267 = 7'hb == idx ? valid_11_1 : _GEN_266; // @[dcache.scala 62:{70,70}]
  wire  _GEN_268 = 7'hc == idx ? valid_12_1 : _GEN_267; // @[dcache.scala 62:{70,70}]
  wire  _GEN_269 = 7'hd == idx ? valid_13_1 : _GEN_268; // @[dcache.scala 62:{70,70}]
  wire  _GEN_270 = 7'he == idx ? valid_14_1 : _GEN_269; // @[dcache.scala 62:{70,70}]
  wire  _GEN_271 = 7'hf == idx ? valid_15_1 : _GEN_270; // @[dcache.scala 62:{70,70}]
  wire  _GEN_272 = 7'h10 == idx ? valid_16_1 : _GEN_271; // @[dcache.scala 62:{70,70}]
  wire  _GEN_273 = 7'h11 == idx ? valid_17_1 : _GEN_272; // @[dcache.scala 62:{70,70}]
  wire  _GEN_274 = 7'h12 == idx ? valid_18_1 : _GEN_273; // @[dcache.scala 62:{70,70}]
  wire  _GEN_275 = 7'h13 == idx ? valid_19_1 : _GEN_274; // @[dcache.scala 62:{70,70}]
  wire  _GEN_276 = 7'h14 == idx ? valid_20_1 : _GEN_275; // @[dcache.scala 62:{70,70}]
  wire  _GEN_277 = 7'h15 == idx ? valid_21_1 : _GEN_276; // @[dcache.scala 62:{70,70}]
  wire  _GEN_278 = 7'h16 == idx ? valid_22_1 : _GEN_277; // @[dcache.scala 62:{70,70}]
  wire  _GEN_279 = 7'h17 == idx ? valid_23_1 : _GEN_278; // @[dcache.scala 62:{70,70}]
  wire  _GEN_280 = 7'h18 == idx ? valid_24_1 : _GEN_279; // @[dcache.scala 62:{70,70}]
  wire  _GEN_281 = 7'h19 == idx ? valid_25_1 : _GEN_280; // @[dcache.scala 62:{70,70}]
  wire  _GEN_282 = 7'h1a == idx ? valid_26_1 : _GEN_281; // @[dcache.scala 62:{70,70}]
  wire  _GEN_283 = 7'h1b == idx ? valid_27_1 : _GEN_282; // @[dcache.scala 62:{70,70}]
  wire  _GEN_284 = 7'h1c == idx ? valid_28_1 : _GEN_283; // @[dcache.scala 62:{70,70}]
  wire  _GEN_285 = 7'h1d == idx ? valid_29_1 : _GEN_284; // @[dcache.scala 62:{70,70}]
  wire  _GEN_286 = 7'h1e == idx ? valid_30_1 : _GEN_285; // @[dcache.scala 62:{70,70}]
  wire  _GEN_287 = 7'h1f == idx ? valid_31_1 : _GEN_286; // @[dcache.scala 62:{70,70}]
  wire  _GEN_288 = 7'h20 == idx ? valid_32_1 : _GEN_287; // @[dcache.scala 62:{70,70}]
  wire  _GEN_289 = 7'h21 == idx ? valid_33_1 : _GEN_288; // @[dcache.scala 62:{70,70}]
  wire  _GEN_290 = 7'h22 == idx ? valid_34_1 : _GEN_289; // @[dcache.scala 62:{70,70}]
  wire  _GEN_291 = 7'h23 == idx ? valid_35_1 : _GEN_290; // @[dcache.scala 62:{70,70}]
  wire  _GEN_292 = 7'h24 == idx ? valid_36_1 : _GEN_291; // @[dcache.scala 62:{70,70}]
  wire  _GEN_293 = 7'h25 == idx ? valid_37_1 : _GEN_292; // @[dcache.scala 62:{70,70}]
  wire  _GEN_294 = 7'h26 == idx ? valid_38_1 : _GEN_293; // @[dcache.scala 62:{70,70}]
  wire  _GEN_295 = 7'h27 == idx ? valid_39_1 : _GEN_294; // @[dcache.scala 62:{70,70}]
  wire  _GEN_296 = 7'h28 == idx ? valid_40_1 : _GEN_295; // @[dcache.scala 62:{70,70}]
  wire  _GEN_297 = 7'h29 == idx ? valid_41_1 : _GEN_296; // @[dcache.scala 62:{70,70}]
  wire  _GEN_298 = 7'h2a == idx ? valid_42_1 : _GEN_297; // @[dcache.scala 62:{70,70}]
  wire  _GEN_299 = 7'h2b == idx ? valid_43_1 : _GEN_298; // @[dcache.scala 62:{70,70}]
  wire  _GEN_300 = 7'h2c == idx ? valid_44_1 : _GEN_299; // @[dcache.scala 62:{70,70}]
  wire  _GEN_301 = 7'h2d == idx ? valid_45_1 : _GEN_300; // @[dcache.scala 62:{70,70}]
  wire  _GEN_302 = 7'h2e == idx ? valid_46_1 : _GEN_301; // @[dcache.scala 62:{70,70}]
  wire  _GEN_303 = 7'h2f == idx ? valid_47_1 : _GEN_302; // @[dcache.scala 62:{70,70}]
  wire  _GEN_304 = 7'h30 == idx ? valid_48_1 : _GEN_303; // @[dcache.scala 62:{70,70}]
  wire  _GEN_305 = 7'h31 == idx ? valid_49_1 : _GEN_304; // @[dcache.scala 62:{70,70}]
  wire  _GEN_306 = 7'h32 == idx ? valid_50_1 : _GEN_305; // @[dcache.scala 62:{70,70}]
  wire  _GEN_307 = 7'h33 == idx ? valid_51_1 : _GEN_306; // @[dcache.scala 62:{70,70}]
  wire  _GEN_308 = 7'h34 == idx ? valid_52_1 : _GEN_307; // @[dcache.scala 62:{70,70}]
  wire  _GEN_309 = 7'h35 == idx ? valid_53_1 : _GEN_308; // @[dcache.scala 62:{70,70}]
  wire  _GEN_310 = 7'h36 == idx ? valid_54_1 : _GEN_309; // @[dcache.scala 62:{70,70}]
  wire  _GEN_311 = 7'h37 == idx ? valid_55_1 : _GEN_310; // @[dcache.scala 62:{70,70}]
  wire  _GEN_312 = 7'h38 == idx ? valid_56_1 : _GEN_311; // @[dcache.scala 62:{70,70}]
  wire  _GEN_313 = 7'h39 == idx ? valid_57_1 : _GEN_312; // @[dcache.scala 62:{70,70}]
  wire  _GEN_314 = 7'h3a == idx ? valid_58_1 : _GEN_313; // @[dcache.scala 62:{70,70}]
  wire  _GEN_315 = 7'h3b == idx ? valid_59_1 : _GEN_314; // @[dcache.scala 62:{70,70}]
  wire  _GEN_316 = 7'h3c == idx ? valid_60_1 : _GEN_315; // @[dcache.scala 62:{70,70}]
  wire  _GEN_317 = 7'h3d == idx ? valid_61_1 : _GEN_316; // @[dcache.scala 62:{70,70}]
  wire  _GEN_318 = 7'h3e == idx ? valid_62_1 : _GEN_317; // @[dcache.scala 62:{70,70}]
  wire  _GEN_319 = 7'h3f == idx ? valid_63_1 : _GEN_318; // @[dcache.scala 62:{70,70}]
  wire  _GEN_320 = 7'h40 == idx ? valid_64_1 : _GEN_319; // @[dcache.scala 62:{70,70}]
  wire  _GEN_321 = 7'h41 == idx ? valid_65_1 : _GEN_320; // @[dcache.scala 62:{70,70}]
  wire  _GEN_322 = 7'h42 == idx ? valid_66_1 : _GEN_321; // @[dcache.scala 62:{70,70}]
  wire  _GEN_323 = 7'h43 == idx ? valid_67_1 : _GEN_322; // @[dcache.scala 62:{70,70}]
  wire  _GEN_324 = 7'h44 == idx ? valid_68_1 : _GEN_323; // @[dcache.scala 62:{70,70}]
  wire  _GEN_325 = 7'h45 == idx ? valid_69_1 : _GEN_324; // @[dcache.scala 62:{70,70}]
  wire  _GEN_326 = 7'h46 == idx ? valid_70_1 : _GEN_325; // @[dcache.scala 62:{70,70}]
  wire  _GEN_327 = 7'h47 == idx ? valid_71_1 : _GEN_326; // @[dcache.scala 62:{70,70}]
  wire  _GEN_328 = 7'h48 == idx ? valid_72_1 : _GEN_327; // @[dcache.scala 62:{70,70}]
  wire  _GEN_329 = 7'h49 == idx ? valid_73_1 : _GEN_328; // @[dcache.scala 62:{70,70}]
  wire  _GEN_330 = 7'h4a == idx ? valid_74_1 : _GEN_329; // @[dcache.scala 62:{70,70}]
  wire  _GEN_331 = 7'h4b == idx ? valid_75_1 : _GEN_330; // @[dcache.scala 62:{70,70}]
  wire  _GEN_332 = 7'h4c == idx ? valid_76_1 : _GEN_331; // @[dcache.scala 62:{70,70}]
  wire  _GEN_333 = 7'h4d == idx ? valid_77_1 : _GEN_332; // @[dcache.scala 62:{70,70}]
  wire  _GEN_334 = 7'h4e == idx ? valid_78_1 : _GEN_333; // @[dcache.scala 62:{70,70}]
  wire  _GEN_335 = 7'h4f == idx ? valid_79_1 : _GEN_334; // @[dcache.scala 62:{70,70}]
  wire  _GEN_336 = 7'h50 == idx ? valid_80_1 : _GEN_335; // @[dcache.scala 62:{70,70}]
  wire  _GEN_337 = 7'h51 == idx ? valid_81_1 : _GEN_336; // @[dcache.scala 62:{70,70}]
  wire  _GEN_338 = 7'h52 == idx ? valid_82_1 : _GEN_337; // @[dcache.scala 62:{70,70}]
  wire  _GEN_339 = 7'h53 == idx ? valid_83_1 : _GEN_338; // @[dcache.scala 62:{70,70}]
  wire  _GEN_340 = 7'h54 == idx ? valid_84_1 : _GEN_339; // @[dcache.scala 62:{70,70}]
  wire  _GEN_341 = 7'h55 == idx ? valid_85_1 : _GEN_340; // @[dcache.scala 62:{70,70}]
  wire  _GEN_342 = 7'h56 == idx ? valid_86_1 : _GEN_341; // @[dcache.scala 62:{70,70}]
  wire  _GEN_343 = 7'h57 == idx ? valid_87_1 : _GEN_342; // @[dcache.scala 62:{70,70}]
  wire  _GEN_344 = 7'h58 == idx ? valid_88_1 : _GEN_343; // @[dcache.scala 62:{70,70}]
  wire  _GEN_345 = 7'h59 == idx ? valid_89_1 : _GEN_344; // @[dcache.scala 62:{70,70}]
  wire  _GEN_346 = 7'h5a == idx ? valid_90_1 : _GEN_345; // @[dcache.scala 62:{70,70}]
  wire  _GEN_347 = 7'h5b == idx ? valid_91_1 : _GEN_346; // @[dcache.scala 62:{70,70}]
  wire  _GEN_348 = 7'h5c == idx ? valid_92_1 : _GEN_347; // @[dcache.scala 62:{70,70}]
  wire  _GEN_349 = 7'h5d == idx ? valid_93_1 : _GEN_348; // @[dcache.scala 62:{70,70}]
  wire  _GEN_350 = 7'h5e == idx ? valid_94_1 : _GEN_349; // @[dcache.scala 62:{70,70}]
  wire  _GEN_351 = 7'h5f == idx ? valid_95_1 : _GEN_350; // @[dcache.scala 62:{70,70}]
  wire  _GEN_352 = 7'h60 == idx ? valid_96_1 : _GEN_351; // @[dcache.scala 62:{70,70}]
  wire  _GEN_353 = 7'h61 == idx ? valid_97_1 : _GEN_352; // @[dcache.scala 62:{70,70}]
  wire  _GEN_354 = 7'h62 == idx ? valid_98_1 : _GEN_353; // @[dcache.scala 62:{70,70}]
  wire  _GEN_355 = 7'h63 == idx ? valid_99_1 : _GEN_354; // @[dcache.scala 62:{70,70}]
  wire  _GEN_356 = 7'h64 == idx ? valid_100_1 : _GEN_355; // @[dcache.scala 62:{70,70}]
  wire  _GEN_357 = 7'h65 == idx ? valid_101_1 : _GEN_356; // @[dcache.scala 62:{70,70}]
  wire  _GEN_358 = 7'h66 == idx ? valid_102_1 : _GEN_357; // @[dcache.scala 62:{70,70}]
  wire  _GEN_359 = 7'h67 == idx ? valid_103_1 : _GEN_358; // @[dcache.scala 62:{70,70}]
  wire  _GEN_360 = 7'h68 == idx ? valid_104_1 : _GEN_359; // @[dcache.scala 62:{70,70}]
  wire  _GEN_361 = 7'h69 == idx ? valid_105_1 : _GEN_360; // @[dcache.scala 62:{70,70}]
  wire  _GEN_362 = 7'h6a == idx ? valid_106_1 : _GEN_361; // @[dcache.scala 62:{70,70}]
  wire  _GEN_363 = 7'h6b == idx ? valid_107_1 : _GEN_362; // @[dcache.scala 62:{70,70}]
  wire  _GEN_364 = 7'h6c == idx ? valid_108_1 : _GEN_363; // @[dcache.scala 62:{70,70}]
  wire  _GEN_365 = 7'h6d == idx ? valid_109_1 : _GEN_364; // @[dcache.scala 62:{70,70}]
  wire  _GEN_366 = 7'h6e == idx ? valid_110_1 : _GEN_365; // @[dcache.scala 62:{70,70}]
  wire  _GEN_367 = 7'h6f == idx ? valid_111_1 : _GEN_366; // @[dcache.scala 62:{70,70}]
  wire  _GEN_368 = 7'h70 == idx ? valid_112_1 : _GEN_367; // @[dcache.scala 62:{70,70}]
  wire  _GEN_369 = 7'h71 == idx ? valid_113_1 : _GEN_368; // @[dcache.scala 62:{70,70}]
  wire  _GEN_370 = 7'h72 == idx ? valid_114_1 : _GEN_369; // @[dcache.scala 62:{70,70}]
  wire  _GEN_371 = 7'h73 == idx ? valid_115_1 : _GEN_370; // @[dcache.scala 62:{70,70}]
  wire  _GEN_372 = 7'h74 == idx ? valid_116_1 : _GEN_371; // @[dcache.scala 62:{70,70}]
  wire  _GEN_373 = 7'h75 == idx ? valid_117_1 : _GEN_372; // @[dcache.scala 62:{70,70}]
  wire  _GEN_374 = 7'h76 == idx ? valid_118_1 : _GEN_373; // @[dcache.scala 62:{70,70}]
  wire  _GEN_375 = 7'h77 == idx ? valid_119_1 : _GEN_374; // @[dcache.scala 62:{70,70}]
  wire  _GEN_376 = 7'h78 == idx ? valid_120_1 : _GEN_375; // @[dcache.scala 62:{70,70}]
  wire  _GEN_377 = 7'h79 == idx ? valid_121_1 : _GEN_376; // @[dcache.scala 62:{70,70}]
  wire  _GEN_378 = 7'h7a == idx ? valid_122_1 : _GEN_377; // @[dcache.scala 62:{70,70}]
  wire  _GEN_379 = 7'h7b == idx ? valid_123_1 : _GEN_378; // @[dcache.scala 62:{70,70}]
  wire  _GEN_380 = 7'h7c == idx ? valid_124_1 : _GEN_379; // @[dcache.scala 62:{70,70}]
  wire  _GEN_381 = 7'h7d == idx ? valid_125_1 : _GEN_380; // @[dcache.scala 62:{70,70}]
  wire  _GEN_382 = 7'h7e == idx ? valid_126_1 : _GEN_381; // @[dcache.scala 62:{70,70}]
  wire  _GEN_383 = 7'h7f == idx ? valid_127_1 : _GEN_382; // @[dcache.scala 62:{70,70}]
  wire [1:0] _hit_T_8 = _GEN_127[41:21] == tag & _GEN_383 ? 2'h1 : 2'h3; // @[dcache.scala 62:16]
  wire [1:0] hit = _GEN_127[20:0] == tag & _GEN_255 ? 2'h0 : _hit_T_8; // @[dcache.scala 61:16]
  wire  _miss_T_2 = state == 3'h1; // @[dcache.scala 64:39]
  wire  miss = hit[1] & state == 3'h1; // @[dcache.scala 64:29]
  reg  way; // @[Reg.scala 35:20]
  wire  hit_way = hit[1] ? way : hit[0]; // @[dcache.scala 68:21]
  wire  _tag_way_T = ~way; // @[dcache.scala 71:22]
  wire [20:0] tag_way = ~way ? _GEN_127[20:0] : _GEN_127[41:21]; // @[dcache.scala 71:17]
  wire [2:0] _state_T_1 = req ? 3'h1 : 3'h0; // @[dcache.scala 76:49]
  wire [2:0] _state_T_2 = io_flush ? 3'h0 : _state_T_1; // @[dcache.scala 76:22]
  wire [2:0] _state_T_4 = miss ? 3'h2 : 3'h0; // @[dcache.scala 77:68]
  wire [2:0] _state_T_5 = uncache ? 3'h0 : _state_T_4; // @[dcache.scala 77:49]
  wire [2:0] _state_T_6 = io_flush ? 3'h0 : _state_T_5; // @[dcache.scala 77:22]
  wire  _GEN_2561 = 7'h0 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_386 = 7'h0 == idx & way ? dirty_0_1 : dirty_0_0; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2562 = 7'h1 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_387 = 7'h1 == idx & _tag_way_T ? dirty_1_0 : _GEN_386; // @[dcache.scala 78:{90,90}]
  wire  _GEN_388 = 7'h1 == idx & way ? dirty_1_1 : _GEN_387; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2565 = 7'h2 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_389 = 7'h2 == idx & _tag_way_T ? dirty_2_0 : _GEN_388; // @[dcache.scala 78:{90,90}]
  wire  _GEN_390 = 7'h2 == idx & way ? dirty_2_1 : _GEN_389; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2568 = 7'h3 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_391 = 7'h3 == idx & _tag_way_T ? dirty_3_0 : _GEN_390; // @[dcache.scala 78:{90,90}]
  wire  _GEN_392 = 7'h3 == idx & way ? dirty_3_1 : _GEN_391; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2571 = 7'h4 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_393 = 7'h4 == idx & _tag_way_T ? dirty_4_0 : _GEN_392; // @[dcache.scala 78:{90,90}]
  wire  _GEN_394 = 7'h4 == idx & way ? dirty_4_1 : _GEN_393; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2574 = 7'h5 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_395 = 7'h5 == idx & _tag_way_T ? dirty_5_0 : _GEN_394; // @[dcache.scala 78:{90,90}]
  wire  _GEN_396 = 7'h5 == idx & way ? dirty_5_1 : _GEN_395; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2577 = 7'h6 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_397 = 7'h6 == idx & _tag_way_T ? dirty_6_0 : _GEN_396; // @[dcache.scala 78:{90,90}]
  wire  _GEN_398 = 7'h6 == idx & way ? dirty_6_1 : _GEN_397; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2580 = 7'h7 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_399 = 7'h7 == idx & _tag_way_T ? dirty_7_0 : _GEN_398; // @[dcache.scala 78:{90,90}]
  wire  _GEN_400 = 7'h7 == idx & way ? dirty_7_1 : _GEN_399; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2583 = 7'h8 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_401 = 7'h8 == idx & _tag_way_T ? dirty_8_0 : _GEN_400; // @[dcache.scala 78:{90,90}]
  wire  _GEN_402 = 7'h8 == idx & way ? dirty_8_1 : _GEN_401; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2586 = 7'h9 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_403 = 7'h9 == idx & _tag_way_T ? dirty_9_0 : _GEN_402; // @[dcache.scala 78:{90,90}]
  wire  _GEN_404 = 7'h9 == idx & way ? dirty_9_1 : _GEN_403; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2589 = 7'ha == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_405 = 7'ha == idx & _tag_way_T ? dirty_10_0 : _GEN_404; // @[dcache.scala 78:{90,90}]
  wire  _GEN_406 = 7'ha == idx & way ? dirty_10_1 : _GEN_405; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2592 = 7'hb == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_407 = 7'hb == idx & _tag_way_T ? dirty_11_0 : _GEN_406; // @[dcache.scala 78:{90,90}]
  wire  _GEN_408 = 7'hb == idx & way ? dirty_11_1 : _GEN_407; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2595 = 7'hc == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_409 = 7'hc == idx & _tag_way_T ? dirty_12_0 : _GEN_408; // @[dcache.scala 78:{90,90}]
  wire  _GEN_410 = 7'hc == idx & way ? dirty_12_1 : _GEN_409; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2598 = 7'hd == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_411 = 7'hd == idx & _tag_way_T ? dirty_13_0 : _GEN_410; // @[dcache.scala 78:{90,90}]
  wire  _GEN_412 = 7'hd == idx & way ? dirty_13_1 : _GEN_411; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2601 = 7'he == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_413 = 7'he == idx & _tag_way_T ? dirty_14_0 : _GEN_412; // @[dcache.scala 78:{90,90}]
  wire  _GEN_414 = 7'he == idx & way ? dirty_14_1 : _GEN_413; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2604 = 7'hf == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_415 = 7'hf == idx & _tag_way_T ? dirty_15_0 : _GEN_414; // @[dcache.scala 78:{90,90}]
  wire  _GEN_416 = 7'hf == idx & way ? dirty_15_1 : _GEN_415; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2607 = 7'h10 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_417 = 7'h10 == idx & _tag_way_T ? dirty_16_0 : _GEN_416; // @[dcache.scala 78:{90,90}]
  wire  _GEN_418 = 7'h10 == idx & way ? dirty_16_1 : _GEN_417; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2610 = 7'h11 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_419 = 7'h11 == idx & _tag_way_T ? dirty_17_0 : _GEN_418; // @[dcache.scala 78:{90,90}]
  wire  _GEN_420 = 7'h11 == idx & way ? dirty_17_1 : _GEN_419; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2613 = 7'h12 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_421 = 7'h12 == idx & _tag_way_T ? dirty_18_0 : _GEN_420; // @[dcache.scala 78:{90,90}]
  wire  _GEN_422 = 7'h12 == idx & way ? dirty_18_1 : _GEN_421; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2616 = 7'h13 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_423 = 7'h13 == idx & _tag_way_T ? dirty_19_0 : _GEN_422; // @[dcache.scala 78:{90,90}]
  wire  _GEN_424 = 7'h13 == idx & way ? dirty_19_1 : _GEN_423; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2619 = 7'h14 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_425 = 7'h14 == idx & _tag_way_T ? dirty_20_0 : _GEN_424; // @[dcache.scala 78:{90,90}]
  wire  _GEN_426 = 7'h14 == idx & way ? dirty_20_1 : _GEN_425; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2622 = 7'h15 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_427 = 7'h15 == idx & _tag_way_T ? dirty_21_0 : _GEN_426; // @[dcache.scala 78:{90,90}]
  wire  _GEN_428 = 7'h15 == idx & way ? dirty_21_1 : _GEN_427; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2625 = 7'h16 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_429 = 7'h16 == idx & _tag_way_T ? dirty_22_0 : _GEN_428; // @[dcache.scala 78:{90,90}]
  wire  _GEN_430 = 7'h16 == idx & way ? dirty_22_1 : _GEN_429; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2628 = 7'h17 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_431 = 7'h17 == idx & _tag_way_T ? dirty_23_0 : _GEN_430; // @[dcache.scala 78:{90,90}]
  wire  _GEN_432 = 7'h17 == idx & way ? dirty_23_1 : _GEN_431; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2631 = 7'h18 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_433 = 7'h18 == idx & _tag_way_T ? dirty_24_0 : _GEN_432; // @[dcache.scala 78:{90,90}]
  wire  _GEN_434 = 7'h18 == idx & way ? dirty_24_1 : _GEN_433; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2634 = 7'h19 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_435 = 7'h19 == idx & _tag_way_T ? dirty_25_0 : _GEN_434; // @[dcache.scala 78:{90,90}]
  wire  _GEN_436 = 7'h19 == idx & way ? dirty_25_1 : _GEN_435; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2637 = 7'h1a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_437 = 7'h1a == idx & _tag_way_T ? dirty_26_0 : _GEN_436; // @[dcache.scala 78:{90,90}]
  wire  _GEN_438 = 7'h1a == idx & way ? dirty_26_1 : _GEN_437; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2640 = 7'h1b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_439 = 7'h1b == idx & _tag_way_T ? dirty_27_0 : _GEN_438; // @[dcache.scala 78:{90,90}]
  wire  _GEN_440 = 7'h1b == idx & way ? dirty_27_1 : _GEN_439; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2643 = 7'h1c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_441 = 7'h1c == idx & _tag_way_T ? dirty_28_0 : _GEN_440; // @[dcache.scala 78:{90,90}]
  wire  _GEN_442 = 7'h1c == idx & way ? dirty_28_1 : _GEN_441; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2646 = 7'h1d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_443 = 7'h1d == idx & _tag_way_T ? dirty_29_0 : _GEN_442; // @[dcache.scala 78:{90,90}]
  wire  _GEN_444 = 7'h1d == idx & way ? dirty_29_1 : _GEN_443; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2649 = 7'h1e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_445 = 7'h1e == idx & _tag_way_T ? dirty_30_0 : _GEN_444; // @[dcache.scala 78:{90,90}]
  wire  _GEN_446 = 7'h1e == idx & way ? dirty_30_1 : _GEN_445; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2652 = 7'h1f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_447 = 7'h1f == idx & _tag_way_T ? dirty_31_0 : _GEN_446; // @[dcache.scala 78:{90,90}]
  wire  _GEN_448 = 7'h1f == idx & way ? dirty_31_1 : _GEN_447; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2655 = 7'h20 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_449 = 7'h20 == idx & _tag_way_T ? dirty_32_0 : _GEN_448; // @[dcache.scala 78:{90,90}]
  wire  _GEN_450 = 7'h20 == idx & way ? dirty_32_1 : _GEN_449; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2658 = 7'h21 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_451 = 7'h21 == idx & _tag_way_T ? dirty_33_0 : _GEN_450; // @[dcache.scala 78:{90,90}]
  wire  _GEN_452 = 7'h21 == idx & way ? dirty_33_1 : _GEN_451; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2661 = 7'h22 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_453 = 7'h22 == idx & _tag_way_T ? dirty_34_0 : _GEN_452; // @[dcache.scala 78:{90,90}]
  wire  _GEN_454 = 7'h22 == idx & way ? dirty_34_1 : _GEN_453; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2664 = 7'h23 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_455 = 7'h23 == idx & _tag_way_T ? dirty_35_0 : _GEN_454; // @[dcache.scala 78:{90,90}]
  wire  _GEN_456 = 7'h23 == idx & way ? dirty_35_1 : _GEN_455; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2667 = 7'h24 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_457 = 7'h24 == idx & _tag_way_T ? dirty_36_0 : _GEN_456; // @[dcache.scala 78:{90,90}]
  wire  _GEN_458 = 7'h24 == idx & way ? dirty_36_1 : _GEN_457; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2670 = 7'h25 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_459 = 7'h25 == idx & _tag_way_T ? dirty_37_0 : _GEN_458; // @[dcache.scala 78:{90,90}]
  wire  _GEN_460 = 7'h25 == idx & way ? dirty_37_1 : _GEN_459; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2673 = 7'h26 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_461 = 7'h26 == idx & _tag_way_T ? dirty_38_0 : _GEN_460; // @[dcache.scala 78:{90,90}]
  wire  _GEN_462 = 7'h26 == idx & way ? dirty_38_1 : _GEN_461; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2676 = 7'h27 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_463 = 7'h27 == idx & _tag_way_T ? dirty_39_0 : _GEN_462; // @[dcache.scala 78:{90,90}]
  wire  _GEN_464 = 7'h27 == idx & way ? dirty_39_1 : _GEN_463; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2679 = 7'h28 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_465 = 7'h28 == idx & _tag_way_T ? dirty_40_0 : _GEN_464; // @[dcache.scala 78:{90,90}]
  wire  _GEN_466 = 7'h28 == idx & way ? dirty_40_1 : _GEN_465; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2682 = 7'h29 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_467 = 7'h29 == idx & _tag_way_T ? dirty_41_0 : _GEN_466; // @[dcache.scala 78:{90,90}]
  wire  _GEN_468 = 7'h29 == idx & way ? dirty_41_1 : _GEN_467; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2685 = 7'h2a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_469 = 7'h2a == idx & _tag_way_T ? dirty_42_0 : _GEN_468; // @[dcache.scala 78:{90,90}]
  wire  _GEN_470 = 7'h2a == idx & way ? dirty_42_1 : _GEN_469; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2688 = 7'h2b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_471 = 7'h2b == idx & _tag_way_T ? dirty_43_0 : _GEN_470; // @[dcache.scala 78:{90,90}]
  wire  _GEN_472 = 7'h2b == idx & way ? dirty_43_1 : _GEN_471; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2691 = 7'h2c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_473 = 7'h2c == idx & _tag_way_T ? dirty_44_0 : _GEN_472; // @[dcache.scala 78:{90,90}]
  wire  _GEN_474 = 7'h2c == idx & way ? dirty_44_1 : _GEN_473; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2694 = 7'h2d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_475 = 7'h2d == idx & _tag_way_T ? dirty_45_0 : _GEN_474; // @[dcache.scala 78:{90,90}]
  wire  _GEN_476 = 7'h2d == idx & way ? dirty_45_1 : _GEN_475; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2697 = 7'h2e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_477 = 7'h2e == idx & _tag_way_T ? dirty_46_0 : _GEN_476; // @[dcache.scala 78:{90,90}]
  wire  _GEN_478 = 7'h2e == idx & way ? dirty_46_1 : _GEN_477; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2700 = 7'h2f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_479 = 7'h2f == idx & _tag_way_T ? dirty_47_0 : _GEN_478; // @[dcache.scala 78:{90,90}]
  wire  _GEN_480 = 7'h2f == idx & way ? dirty_47_1 : _GEN_479; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2703 = 7'h30 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_481 = 7'h30 == idx & _tag_way_T ? dirty_48_0 : _GEN_480; // @[dcache.scala 78:{90,90}]
  wire  _GEN_482 = 7'h30 == idx & way ? dirty_48_1 : _GEN_481; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2706 = 7'h31 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_483 = 7'h31 == idx & _tag_way_T ? dirty_49_0 : _GEN_482; // @[dcache.scala 78:{90,90}]
  wire  _GEN_484 = 7'h31 == idx & way ? dirty_49_1 : _GEN_483; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2709 = 7'h32 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_485 = 7'h32 == idx & _tag_way_T ? dirty_50_0 : _GEN_484; // @[dcache.scala 78:{90,90}]
  wire  _GEN_486 = 7'h32 == idx & way ? dirty_50_1 : _GEN_485; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2712 = 7'h33 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_487 = 7'h33 == idx & _tag_way_T ? dirty_51_0 : _GEN_486; // @[dcache.scala 78:{90,90}]
  wire  _GEN_488 = 7'h33 == idx & way ? dirty_51_1 : _GEN_487; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2715 = 7'h34 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_489 = 7'h34 == idx & _tag_way_T ? dirty_52_0 : _GEN_488; // @[dcache.scala 78:{90,90}]
  wire  _GEN_490 = 7'h34 == idx & way ? dirty_52_1 : _GEN_489; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2718 = 7'h35 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_491 = 7'h35 == idx & _tag_way_T ? dirty_53_0 : _GEN_490; // @[dcache.scala 78:{90,90}]
  wire  _GEN_492 = 7'h35 == idx & way ? dirty_53_1 : _GEN_491; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2721 = 7'h36 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_493 = 7'h36 == idx & _tag_way_T ? dirty_54_0 : _GEN_492; // @[dcache.scala 78:{90,90}]
  wire  _GEN_494 = 7'h36 == idx & way ? dirty_54_1 : _GEN_493; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2724 = 7'h37 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_495 = 7'h37 == idx & _tag_way_T ? dirty_55_0 : _GEN_494; // @[dcache.scala 78:{90,90}]
  wire  _GEN_496 = 7'h37 == idx & way ? dirty_55_1 : _GEN_495; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2727 = 7'h38 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_497 = 7'h38 == idx & _tag_way_T ? dirty_56_0 : _GEN_496; // @[dcache.scala 78:{90,90}]
  wire  _GEN_498 = 7'h38 == idx & way ? dirty_56_1 : _GEN_497; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2730 = 7'h39 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_499 = 7'h39 == idx & _tag_way_T ? dirty_57_0 : _GEN_498; // @[dcache.scala 78:{90,90}]
  wire  _GEN_500 = 7'h39 == idx & way ? dirty_57_1 : _GEN_499; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2733 = 7'h3a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_501 = 7'h3a == idx & _tag_way_T ? dirty_58_0 : _GEN_500; // @[dcache.scala 78:{90,90}]
  wire  _GEN_502 = 7'h3a == idx & way ? dirty_58_1 : _GEN_501; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2736 = 7'h3b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_503 = 7'h3b == idx & _tag_way_T ? dirty_59_0 : _GEN_502; // @[dcache.scala 78:{90,90}]
  wire  _GEN_504 = 7'h3b == idx & way ? dirty_59_1 : _GEN_503; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2739 = 7'h3c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_505 = 7'h3c == idx & _tag_way_T ? dirty_60_0 : _GEN_504; // @[dcache.scala 78:{90,90}]
  wire  _GEN_506 = 7'h3c == idx & way ? dirty_60_1 : _GEN_505; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2742 = 7'h3d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_507 = 7'h3d == idx & _tag_way_T ? dirty_61_0 : _GEN_506; // @[dcache.scala 78:{90,90}]
  wire  _GEN_508 = 7'h3d == idx & way ? dirty_61_1 : _GEN_507; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2745 = 7'h3e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_509 = 7'h3e == idx & _tag_way_T ? dirty_62_0 : _GEN_508; // @[dcache.scala 78:{90,90}]
  wire  _GEN_510 = 7'h3e == idx & way ? dirty_62_1 : _GEN_509; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2748 = 7'h3f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_511 = 7'h3f == idx & _tag_way_T ? dirty_63_0 : _GEN_510; // @[dcache.scala 78:{90,90}]
  wire  _GEN_512 = 7'h3f == idx & way ? dirty_63_1 : _GEN_511; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2751 = 7'h40 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_513 = 7'h40 == idx & _tag_way_T ? dirty_64_0 : _GEN_512; // @[dcache.scala 78:{90,90}]
  wire  _GEN_514 = 7'h40 == idx & way ? dirty_64_1 : _GEN_513; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2754 = 7'h41 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_515 = 7'h41 == idx & _tag_way_T ? dirty_65_0 : _GEN_514; // @[dcache.scala 78:{90,90}]
  wire  _GEN_516 = 7'h41 == idx & way ? dirty_65_1 : _GEN_515; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2757 = 7'h42 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_517 = 7'h42 == idx & _tag_way_T ? dirty_66_0 : _GEN_516; // @[dcache.scala 78:{90,90}]
  wire  _GEN_518 = 7'h42 == idx & way ? dirty_66_1 : _GEN_517; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2760 = 7'h43 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_519 = 7'h43 == idx & _tag_way_T ? dirty_67_0 : _GEN_518; // @[dcache.scala 78:{90,90}]
  wire  _GEN_520 = 7'h43 == idx & way ? dirty_67_1 : _GEN_519; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2763 = 7'h44 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_521 = 7'h44 == idx & _tag_way_T ? dirty_68_0 : _GEN_520; // @[dcache.scala 78:{90,90}]
  wire  _GEN_522 = 7'h44 == idx & way ? dirty_68_1 : _GEN_521; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2766 = 7'h45 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_523 = 7'h45 == idx & _tag_way_T ? dirty_69_0 : _GEN_522; // @[dcache.scala 78:{90,90}]
  wire  _GEN_524 = 7'h45 == idx & way ? dirty_69_1 : _GEN_523; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2769 = 7'h46 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_525 = 7'h46 == idx & _tag_way_T ? dirty_70_0 : _GEN_524; // @[dcache.scala 78:{90,90}]
  wire  _GEN_526 = 7'h46 == idx & way ? dirty_70_1 : _GEN_525; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2772 = 7'h47 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_527 = 7'h47 == idx & _tag_way_T ? dirty_71_0 : _GEN_526; // @[dcache.scala 78:{90,90}]
  wire  _GEN_528 = 7'h47 == idx & way ? dirty_71_1 : _GEN_527; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2775 = 7'h48 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_529 = 7'h48 == idx & _tag_way_T ? dirty_72_0 : _GEN_528; // @[dcache.scala 78:{90,90}]
  wire  _GEN_530 = 7'h48 == idx & way ? dirty_72_1 : _GEN_529; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2778 = 7'h49 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_531 = 7'h49 == idx & _tag_way_T ? dirty_73_0 : _GEN_530; // @[dcache.scala 78:{90,90}]
  wire  _GEN_532 = 7'h49 == idx & way ? dirty_73_1 : _GEN_531; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2781 = 7'h4a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_533 = 7'h4a == idx & _tag_way_T ? dirty_74_0 : _GEN_532; // @[dcache.scala 78:{90,90}]
  wire  _GEN_534 = 7'h4a == idx & way ? dirty_74_1 : _GEN_533; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2784 = 7'h4b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_535 = 7'h4b == idx & _tag_way_T ? dirty_75_0 : _GEN_534; // @[dcache.scala 78:{90,90}]
  wire  _GEN_536 = 7'h4b == idx & way ? dirty_75_1 : _GEN_535; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2787 = 7'h4c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_537 = 7'h4c == idx & _tag_way_T ? dirty_76_0 : _GEN_536; // @[dcache.scala 78:{90,90}]
  wire  _GEN_538 = 7'h4c == idx & way ? dirty_76_1 : _GEN_537; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2790 = 7'h4d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_539 = 7'h4d == idx & _tag_way_T ? dirty_77_0 : _GEN_538; // @[dcache.scala 78:{90,90}]
  wire  _GEN_540 = 7'h4d == idx & way ? dirty_77_1 : _GEN_539; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2793 = 7'h4e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_541 = 7'h4e == idx & _tag_way_T ? dirty_78_0 : _GEN_540; // @[dcache.scala 78:{90,90}]
  wire  _GEN_542 = 7'h4e == idx & way ? dirty_78_1 : _GEN_541; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2796 = 7'h4f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_543 = 7'h4f == idx & _tag_way_T ? dirty_79_0 : _GEN_542; // @[dcache.scala 78:{90,90}]
  wire  _GEN_544 = 7'h4f == idx & way ? dirty_79_1 : _GEN_543; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2799 = 7'h50 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_545 = 7'h50 == idx & _tag_way_T ? dirty_80_0 : _GEN_544; // @[dcache.scala 78:{90,90}]
  wire  _GEN_546 = 7'h50 == idx & way ? dirty_80_1 : _GEN_545; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2802 = 7'h51 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_547 = 7'h51 == idx & _tag_way_T ? dirty_81_0 : _GEN_546; // @[dcache.scala 78:{90,90}]
  wire  _GEN_548 = 7'h51 == idx & way ? dirty_81_1 : _GEN_547; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2805 = 7'h52 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_549 = 7'h52 == idx & _tag_way_T ? dirty_82_0 : _GEN_548; // @[dcache.scala 78:{90,90}]
  wire  _GEN_550 = 7'h52 == idx & way ? dirty_82_1 : _GEN_549; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2808 = 7'h53 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_551 = 7'h53 == idx & _tag_way_T ? dirty_83_0 : _GEN_550; // @[dcache.scala 78:{90,90}]
  wire  _GEN_552 = 7'h53 == idx & way ? dirty_83_1 : _GEN_551; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2811 = 7'h54 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_553 = 7'h54 == idx & _tag_way_T ? dirty_84_0 : _GEN_552; // @[dcache.scala 78:{90,90}]
  wire  _GEN_554 = 7'h54 == idx & way ? dirty_84_1 : _GEN_553; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2814 = 7'h55 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_555 = 7'h55 == idx & _tag_way_T ? dirty_85_0 : _GEN_554; // @[dcache.scala 78:{90,90}]
  wire  _GEN_556 = 7'h55 == idx & way ? dirty_85_1 : _GEN_555; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2817 = 7'h56 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_557 = 7'h56 == idx & _tag_way_T ? dirty_86_0 : _GEN_556; // @[dcache.scala 78:{90,90}]
  wire  _GEN_558 = 7'h56 == idx & way ? dirty_86_1 : _GEN_557; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2820 = 7'h57 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_559 = 7'h57 == idx & _tag_way_T ? dirty_87_0 : _GEN_558; // @[dcache.scala 78:{90,90}]
  wire  _GEN_560 = 7'h57 == idx & way ? dirty_87_1 : _GEN_559; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2823 = 7'h58 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_561 = 7'h58 == idx & _tag_way_T ? dirty_88_0 : _GEN_560; // @[dcache.scala 78:{90,90}]
  wire  _GEN_562 = 7'h58 == idx & way ? dirty_88_1 : _GEN_561; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2826 = 7'h59 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_563 = 7'h59 == idx & _tag_way_T ? dirty_89_0 : _GEN_562; // @[dcache.scala 78:{90,90}]
  wire  _GEN_564 = 7'h59 == idx & way ? dirty_89_1 : _GEN_563; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2829 = 7'h5a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_565 = 7'h5a == idx & _tag_way_T ? dirty_90_0 : _GEN_564; // @[dcache.scala 78:{90,90}]
  wire  _GEN_566 = 7'h5a == idx & way ? dirty_90_1 : _GEN_565; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2832 = 7'h5b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_567 = 7'h5b == idx & _tag_way_T ? dirty_91_0 : _GEN_566; // @[dcache.scala 78:{90,90}]
  wire  _GEN_568 = 7'h5b == idx & way ? dirty_91_1 : _GEN_567; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2835 = 7'h5c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_569 = 7'h5c == idx & _tag_way_T ? dirty_92_0 : _GEN_568; // @[dcache.scala 78:{90,90}]
  wire  _GEN_570 = 7'h5c == idx & way ? dirty_92_1 : _GEN_569; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2838 = 7'h5d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_571 = 7'h5d == idx & _tag_way_T ? dirty_93_0 : _GEN_570; // @[dcache.scala 78:{90,90}]
  wire  _GEN_572 = 7'h5d == idx & way ? dirty_93_1 : _GEN_571; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2841 = 7'h5e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_573 = 7'h5e == idx & _tag_way_T ? dirty_94_0 : _GEN_572; // @[dcache.scala 78:{90,90}]
  wire  _GEN_574 = 7'h5e == idx & way ? dirty_94_1 : _GEN_573; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2844 = 7'h5f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_575 = 7'h5f == idx & _tag_way_T ? dirty_95_0 : _GEN_574; // @[dcache.scala 78:{90,90}]
  wire  _GEN_576 = 7'h5f == idx & way ? dirty_95_1 : _GEN_575; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2847 = 7'h60 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_577 = 7'h60 == idx & _tag_way_T ? dirty_96_0 : _GEN_576; // @[dcache.scala 78:{90,90}]
  wire  _GEN_578 = 7'h60 == idx & way ? dirty_96_1 : _GEN_577; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2850 = 7'h61 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_579 = 7'h61 == idx & _tag_way_T ? dirty_97_0 : _GEN_578; // @[dcache.scala 78:{90,90}]
  wire  _GEN_580 = 7'h61 == idx & way ? dirty_97_1 : _GEN_579; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2853 = 7'h62 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_581 = 7'h62 == idx & _tag_way_T ? dirty_98_0 : _GEN_580; // @[dcache.scala 78:{90,90}]
  wire  _GEN_582 = 7'h62 == idx & way ? dirty_98_1 : _GEN_581; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2856 = 7'h63 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_583 = 7'h63 == idx & _tag_way_T ? dirty_99_0 : _GEN_582; // @[dcache.scala 78:{90,90}]
  wire  _GEN_584 = 7'h63 == idx & way ? dirty_99_1 : _GEN_583; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2859 = 7'h64 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_585 = 7'h64 == idx & _tag_way_T ? dirty_100_0 : _GEN_584; // @[dcache.scala 78:{90,90}]
  wire  _GEN_586 = 7'h64 == idx & way ? dirty_100_1 : _GEN_585; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2862 = 7'h65 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_587 = 7'h65 == idx & _tag_way_T ? dirty_101_0 : _GEN_586; // @[dcache.scala 78:{90,90}]
  wire  _GEN_588 = 7'h65 == idx & way ? dirty_101_1 : _GEN_587; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2865 = 7'h66 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_589 = 7'h66 == idx & _tag_way_T ? dirty_102_0 : _GEN_588; // @[dcache.scala 78:{90,90}]
  wire  _GEN_590 = 7'h66 == idx & way ? dirty_102_1 : _GEN_589; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2868 = 7'h67 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_591 = 7'h67 == idx & _tag_way_T ? dirty_103_0 : _GEN_590; // @[dcache.scala 78:{90,90}]
  wire  _GEN_592 = 7'h67 == idx & way ? dirty_103_1 : _GEN_591; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2871 = 7'h68 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_593 = 7'h68 == idx & _tag_way_T ? dirty_104_0 : _GEN_592; // @[dcache.scala 78:{90,90}]
  wire  _GEN_594 = 7'h68 == idx & way ? dirty_104_1 : _GEN_593; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2874 = 7'h69 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_595 = 7'h69 == idx & _tag_way_T ? dirty_105_0 : _GEN_594; // @[dcache.scala 78:{90,90}]
  wire  _GEN_596 = 7'h69 == idx & way ? dirty_105_1 : _GEN_595; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2877 = 7'h6a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_597 = 7'h6a == idx & _tag_way_T ? dirty_106_0 : _GEN_596; // @[dcache.scala 78:{90,90}]
  wire  _GEN_598 = 7'h6a == idx & way ? dirty_106_1 : _GEN_597; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2880 = 7'h6b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_599 = 7'h6b == idx & _tag_way_T ? dirty_107_0 : _GEN_598; // @[dcache.scala 78:{90,90}]
  wire  _GEN_600 = 7'h6b == idx & way ? dirty_107_1 : _GEN_599; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2883 = 7'h6c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_601 = 7'h6c == idx & _tag_way_T ? dirty_108_0 : _GEN_600; // @[dcache.scala 78:{90,90}]
  wire  _GEN_602 = 7'h6c == idx & way ? dirty_108_1 : _GEN_601; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2886 = 7'h6d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_603 = 7'h6d == idx & _tag_way_T ? dirty_109_0 : _GEN_602; // @[dcache.scala 78:{90,90}]
  wire  _GEN_604 = 7'h6d == idx & way ? dirty_109_1 : _GEN_603; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2889 = 7'h6e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_605 = 7'h6e == idx & _tag_way_T ? dirty_110_0 : _GEN_604; // @[dcache.scala 78:{90,90}]
  wire  _GEN_606 = 7'h6e == idx & way ? dirty_110_1 : _GEN_605; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2892 = 7'h6f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_607 = 7'h6f == idx & _tag_way_T ? dirty_111_0 : _GEN_606; // @[dcache.scala 78:{90,90}]
  wire  _GEN_608 = 7'h6f == idx & way ? dirty_111_1 : _GEN_607; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2895 = 7'h70 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_609 = 7'h70 == idx & _tag_way_T ? dirty_112_0 : _GEN_608; // @[dcache.scala 78:{90,90}]
  wire  _GEN_610 = 7'h70 == idx & way ? dirty_112_1 : _GEN_609; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2898 = 7'h71 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_611 = 7'h71 == idx & _tag_way_T ? dirty_113_0 : _GEN_610; // @[dcache.scala 78:{90,90}]
  wire  _GEN_612 = 7'h71 == idx & way ? dirty_113_1 : _GEN_611; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2901 = 7'h72 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_613 = 7'h72 == idx & _tag_way_T ? dirty_114_0 : _GEN_612; // @[dcache.scala 78:{90,90}]
  wire  _GEN_614 = 7'h72 == idx & way ? dirty_114_1 : _GEN_613; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2904 = 7'h73 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_615 = 7'h73 == idx & _tag_way_T ? dirty_115_0 : _GEN_614; // @[dcache.scala 78:{90,90}]
  wire  _GEN_616 = 7'h73 == idx & way ? dirty_115_1 : _GEN_615; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2907 = 7'h74 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_617 = 7'h74 == idx & _tag_way_T ? dirty_116_0 : _GEN_616; // @[dcache.scala 78:{90,90}]
  wire  _GEN_618 = 7'h74 == idx & way ? dirty_116_1 : _GEN_617; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2910 = 7'h75 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_619 = 7'h75 == idx & _tag_way_T ? dirty_117_0 : _GEN_618; // @[dcache.scala 78:{90,90}]
  wire  _GEN_620 = 7'h75 == idx & way ? dirty_117_1 : _GEN_619; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2913 = 7'h76 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_621 = 7'h76 == idx & _tag_way_T ? dirty_118_0 : _GEN_620; // @[dcache.scala 78:{90,90}]
  wire  _GEN_622 = 7'h76 == idx & way ? dirty_118_1 : _GEN_621; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2916 = 7'h77 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_623 = 7'h77 == idx & _tag_way_T ? dirty_119_0 : _GEN_622; // @[dcache.scala 78:{90,90}]
  wire  _GEN_624 = 7'h77 == idx & way ? dirty_119_1 : _GEN_623; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2919 = 7'h78 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_625 = 7'h78 == idx & _tag_way_T ? dirty_120_0 : _GEN_624; // @[dcache.scala 78:{90,90}]
  wire  _GEN_626 = 7'h78 == idx & way ? dirty_120_1 : _GEN_625; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2922 = 7'h79 == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_627 = 7'h79 == idx & _tag_way_T ? dirty_121_0 : _GEN_626; // @[dcache.scala 78:{90,90}]
  wire  _GEN_628 = 7'h79 == idx & way ? dirty_121_1 : _GEN_627; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2925 = 7'h7a == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_629 = 7'h7a == idx & _tag_way_T ? dirty_122_0 : _GEN_628; // @[dcache.scala 78:{90,90}]
  wire  _GEN_630 = 7'h7a == idx & way ? dirty_122_1 : _GEN_629; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2928 = 7'h7b == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_631 = 7'h7b == idx & _tag_way_T ? dirty_123_0 : _GEN_630; // @[dcache.scala 78:{90,90}]
  wire  _GEN_632 = 7'h7b == idx & way ? dirty_123_1 : _GEN_631; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2931 = 7'h7c == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_633 = 7'h7c == idx & _tag_way_T ? dirty_124_0 : _GEN_632; // @[dcache.scala 78:{90,90}]
  wire  _GEN_634 = 7'h7c == idx & way ? dirty_124_1 : _GEN_633; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2934 = 7'h7d == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_635 = 7'h7d == idx & _tag_way_T ? dirty_125_0 : _GEN_634; // @[dcache.scala 78:{90,90}]
  wire  _GEN_636 = 7'h7d == idx & way ? dirty_125_1 : _GEN_635; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2937 = 7'h7e == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_637 = 7'h7e == idx & _tag_way_T ? dirty_126_0 : _GEN_636; // @[dcache.scala 78:{90,90}]
  wire  _GEN_638 = 7'h7e == idx & way ? dirty_126_1 : _GEN_637; // @[dcache.scala 78:{90,90}]
  wire  _GEN_2940 = 7'h7f == idx; // @[dcache.scala 78:{90,90}]
  wire  _GEN_639 = 7'h7f == idx & _tag_way_T ? dirty_127_0 : _GEN_638; // @[dcache.scala 78:{90,90}]
  wire  _GEN_640 = 7'h7f == idx & way ? dirty_127_1 : _GEN_639; // @[dcache.scala 78:{90,90}]
  wire [2:0] _state_T_19 = rstate == 3'h6 & (_GEN_640 & wstate == 3'h6 | ~_GEN_640) ? 3'h3 : 3'h2; // @[dcache.scala 78:49]
  wire [2:0] _state_T_22 = 3'h0 == state ? _state_T_2 : 3'h0; // @[Mux.scala 81:58]
  wire  _rstate_T_1 = state == 3'h2; // @[dcache.scala 83:53]
  wire  _rstate_T_2 = io_mem_ar_ready & io_mem_ar_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _rstate_T_4 = state == 3'h2 & _rstate_T_2 ? 3'h4 : 3'h0; // @[dcache.scala 83:46]
  wire [2:0] _rstate_T_5 = io_flush ? 3'h0 : _rstate_T_4; // @[dcache.scala 83:19]
  wire  _rstate_T_7 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _rstate_T_8 = _rstate_T_7 ? 3'h5 : 3'h4; // @[dcache.scala 84:46]
  wire [2:0] _rstate_T_9 = io_flush ? 3'h0 : _rstate_T_8; // @[dcache.scala 84:19]
  wire [2:0] _rstate_T_12 = _rstate_T_7 ? 3'h6 : 3'h5; // @[dcache.scala 85:46]
  wire [2:0] _rstate_T_19 = 3'h0 == rstate ? _rstate_T_5 : 3'h0; // @[Mux.scala 81:58]
  wire  _wstate_T_2 = io_mem_aw_ready & io_mem_aw_valid; // @[Decoupled.scala 52:35]
  wire  _wstate_T_4 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _wstate_T_6 = _rstate_T_1 & _wstate_T_2 & _wstate_T_4 ? 3'h4 : 3'h0; // @[dcache.scala 90:46]
  wire [2:0] _wstate_T_7 = io_flush ? 3'h0 : _wstate_T_6; // @[dcache.scala 90:19]
  wire [2:0] _wstate_T_10 = _wstate_T_4 ? 3'h5 : 3'h4; // @[dcache.scala 91:46]
  wire [2:0] _wstate_T_11 = io_flush ? 3'h0 : _wstate_T_10; // @[dcache.scala 91:19]
  wire  _wstate_T_13 = io_mem_b_ready & io_mem_b_valid; // @[Decoupled.scala 52:35]
  wire [2:0] _wstate_T_14 = _wstate_T_13 ? 3'h6 : 3'h5; // @[dcache.scala 92:46]
  wire [2:0] _wstate_T_21 = 3'h0 == wstate ? _wstate_T_7 : 3'h0; // @[Mux.scala 81:58]
  wire  _valid_T_1 = ~uncache; // @[dcache.scala 98:46]
  wire  _valid_T_2 = _rstate_T_1 & ~uncache; // @[dcache.scala 98:43]
  wire  _GEN_898 = _GEN_2561 & way ? valid_0_1 : valid_0_0; // @[dcache.scala 98:{25,25}]
  wire  _GEN_899 = _GEN_2562 & _tag_way_T ? valid_1_0 : _GEN_898; // @[dcache.scala 98:{25,25}]
  wire  _GEN_900 = _GEN_2562 & way ? valid_1_1 : _GEN_899; // @[dcache.scala 98:{25,25}]
  wire  _GEN_901 = _GEN_2565 & _tag_way_T ? valid_2_0 : _GEN_900; // @[dcache.scala 98:{25,25}]
  wire  _GEN_902 = _GEN_2565 & way ? valid_2_1 : _GEN_901; // @[dcache.scala 98:{25,25}]
  wire  _GEN_903 = _GEN_2568 & _tag_way_T ? valid_3_0 : _GEN_902; // @[dcache.scala 98:{25,25}]
  wire  _GEN_904 = _GEN_2568 & way ? valid_3_1 : _GEN_903; // @[dcache.scala 98:{25,25}]
  wire  _GEN_905 = _GEN_2571 & _tag_way_T ? valid_4_0 : _GEN_904; // @[dcache.scala 98:{25,25}]
  wire  _GEN_906 = _GEN_2571 & way ? valid_4_1 : _GEN_905; // @[dcache.scala 98:{25,25}]
  wire  _GEN_907 = _GEN_2574 & _tag_way_T ? valid_5_0 : _GEN_906; // @[dcache.scala 98:{25,25}]
  wire  _GEN_908 = _GEN_2574 & way ? valid_5_1 : _GEN_907; // @[dcache.scala 98:{25,25}]
  wire  _GEN_909 = _GEN_2577 & _tag_way_T ? valid_6_0 : _GEN_908; // @[dcache.scala 98:{25,25}]
  wire  _GEN_910 = _GEN_2577 & way ? valid_6_1 : _GEN_909; // @[dcache.scala 98:{25,25}]
  wire  _GEN_911 = _GEN_2580 & _tag_way_T ? valid_7_0 : _GEN_910; // @[dcache.scala 98:{25,25}]
  wire  _GEN_912 = _GEN_2580 & way ? valid_7_1 : _GEN_911; // @[dcache.scala 98:{25,25}]
  wire  _GEN_913 = _GEN_2583 & _tag_way_T ? valid_8_0 : _GEN_912; // @[dcache.scala 98:{25,25}]
  wire  _GEN_914 = _GEN_2583 & way ? valid_8_1 : _GEN_913; // @[dcache.scala 98:{25,25}]
  wire  _GEN_915 = _GEN_2586 & _tag_way_T ? valid_9_0 : _GEN_914; // @[dcache.scala 98:{25,25}]
  wire  _GEN_916 = _GEN_2586 & way ? valid_9_1 : _GEN_915; // @[dcache.scala 98:{25,25}]
  wire  _GEN_917 = _GEN_2589 & _tag_way_T ? valid_10_0 : _GEN_916; // @[dcache.scala 98:{25,25}]
  wire  _GEN_918 = _GEN_2589 & way ? valid_10_1 : _GEN_917; // @[dcache.scala 98:{25,25}]
  wire  _GEN_919 = _GEN_2592 & _tag_way_T ? valid_11_0 : _GEN_918; // @[dcache.scala 98:{25,25}]
  wire  _GEN_920 = _GEN_2592 & way ? valid_11_1 : _GEN_919; // @[dcache.scala 98:{25,25}]
  wire  _GEN_921 = _GEN_2595 & _tag_way_T ? valid_12_0 : _GEN_920; // @[dcache.scala 98:{25,25}]
  wire  _GEN_922 = _GEN_2595 & way ? valid_12_1 : _GEN_921; // @[dcache.scala 98:{25,25}]
  wire  _GEN_923 = _GEN_2598 & _tag_way_T ? valid_13_0 : _GEN_922; // @[dcache.scala 98:{25,25}]
  wire  _GEN_924 = _GEN_2598 & way ? valid_13_1 : _GEN_923; // @[dcache.scala 98:{25,25}]
  wire  _GEN_925 = _GEN_2601 & _tag_way_T ? valid_14_0 : _GEN_924; // @[dcache.scala 98:{25,25}]
  wire  _GEN_926 = _GEN_2601 & way ? valid_14_1 : _GEN_925; // @[dcache.scala 98:{25,25}]
  wire  _GEN_927 = _GEN_2604 & _tag_way_T ? valid_15_0 : _GEN_926; // @[dcache.scala 98:{25,25}]
  wire  _GEN_928 = _GEN_2604 & way ? valid_15_1 : _GEN_927; // @[dcache.scala 98:{25,25}]
  wire  _GEN_929 = _GEN_2607 & _tag_way_T ? valid_16_0 : _GEN_928; // @[dcache.scala 98:{25,25}]
  wire  _GEN_930 = _GEN_2607 & way ? valid_16_1 : _GEN_929; // @[dcache.scala 98:{25,25}]
  wire  _GEN_931 = _GEN_2610 & _tag_way_T ? valid_17_0 : _GEN_930; // @[dcache.scala 98:{25,25}]
  wire  _GEN_932 = _GEN_2610 & way ? valid_17_1 : _GEN_931; // @[dcache.scala 98:{25,25}]
  wire  _GEN_933 = _GEN_2613 & _tag_way_T ? valid_18_0 : _GEN_932; // @[dcache.scala 98:{25,25}]
  wire  _GEN_934 = _GEN_2613 & way ? valid_18_1 : _GEN_933; // @[dcache.scala 98:{25,25}]
  wire  _GEN_935 = _GEN_2616 & _tag_way_T ? valid_19_0 : _GEN_934; // @[dcache.scala 98:{25,25}]
  wire  _GEN_936 = _GEN_2616 & way ? valid_19_1 : _GEN_935; // @[dcache.scala 98:{25,25}]
  wire  _GEN_937 = _GEN_2619 & _tag_way_T ? valid_20_0 : _GEN_936; // @[dcache.scala 98:{25,25}]
  wire  _GEN_938 = _GEN_2619 & way ? valid_20_1 : _GEN_937; // @[dcache.scala 98:{25,25}]
  wire  _GEN_939 = _GEN_2622 & _tag_way_T ? valid_21_0 : _GEN_938; // @[dcache.scala 98:{25,25}]
  wire  _GEN_940 = _GEN_2622 & way ? valid_21_1 : _GEN_939; // @[dcache.scala 98:{25,25}]
  wire  _GEN_941 = _GEN_2625 & _tag_way_T ? valid_22_0 : _GEN_940; // @[dcache.scala 98:{25,25}]
  wire  _GEN_942 = _GEN_2625 & way ? valid_22_1 : _GEN_941; // @[dcache.scala 98:{25,25}]
  wire  _GEN_943 = _GEN_2628 & _tag_way_T ? valid_23_0 : _GEN_942; // @[dcache.scala 98:{25,25}]
  wire  _GEN_944 = _GEN_2628 & way ? valid_23_1 : _GEN_943; // @[dcache.scala 98:{25,25}]
  wire  _GEN_945 = _GEN_2631 & _tag_way_T ? valid_24_0 : _GEN_944; // @[dcache.scala 98:{25,25}]
  wire  _GEN_946 = _GEN_2631 & way ? valid_24_1 : _GEN_945; // @[dcache.scala 98:{25,25}]
  wire  _GEN_947 = _GEN_2634 & _tag_way_T ? valid_25_0 : _GEN_946; // @[dcache.scala 98:{25,25}]
  wire  _GEN_948 = _GEN_2634 & way ? valid_25_1 : _GEN_947; // @[dcache.scala 98:{25,25}]
  wire  _GEN_949 = _GEN_2637 & _tag_way_T ? valid_26_0 : _GEN_948; // @[dcache.scala 98:{25,25}]
  wire  _GEN_950 = _GEN_2637 & way ? valid_26_1 : _GEN_949; // @[dcache.scala 98:{25,25}]
  wire  _GEN_951 = _GEN_2640 & _tag_way_T ? valid_27_0 : _GEN_950; // @[dcache.scala 98:{25,25}]
  wire  _GEN_952 = _GEN_2640 & way ? valid_27_1 : _GEN_951; // @[dcache.scala 98:{25,25}]
  wire  _GEN_953 = _GEN_2643 & _tag_way_T ? valid_28_0 : _GEN_952; // @[dcache.scala 98:{25,25}]
  wire  _GEN_954 = _GEN_2643 & way ? valid_28_1 : _GEN_953; // @[dcache.scala 98:{25,25}]
  wire  _GEN_955 = _GEN_2646 & _tag_way_T ? valid_29_0 : _GEN_954; // @[dcache.scala 98:{25,25}]
  wire  _GEN_956 = _GEN_2646 & way ? valid_29_1 : _GEN_955; // @[dcache.scala 98:{25,25}]
  wire  _GEN_957 = _GEN_2649 & _tag_way_T ? valid_30_0 : _GEN_956; // @[dcache.scala 98:{25,25}]
  wire  _GEN_958 = _GEN_2649 & way ? valid_30_1 : _GEN_957; // @[dcache.scala 98:{25,25}]
  wire  _GEN_959 = _GEN_2652 & _tag_way_T ? valid_31_0 : _GEN_958; // @[dcache.scala 98:{25,25}]
  wire  _GEN_960 = _GEN_2652 & way ? valid_31_1 : _GEN_959; // @[dcache.scala 98:{25,25}]
  wire  _GEN_961 = _GEN_2655 & _tag_way_T ? valid_32_0 : _GEN_960; // @[dcache.scala 98:{25,25}]
  wire  _GEN_962 = _GEN_2655 & way ? valid_32_1 : _GEN_961; // @[dcache.scala 98:{25,25}]
  wire  _GEN_963 = _GEN_2658 & _tag_way_T ? valid_33_0 : _GEN_962; // @[dcache.scala 98:{25,25}]
  wire  _GEN_964 = _GEN_2658 & way ? valid_33_1 : _GEN_963; // @[dcache.scala 98:{25,25}]
  wire  _GEN_965 = _GEN_2661 & _tag_way_T ? valid_34_0 : _GEN_964; // @[dcache.scala 98:{25,25}]
  wire  _GEN_966 = _GEN_2661 & way ? valid_34_1 : _GEN_965; // @[dcache.scala 98:{25,25}]
  wire  _GEN_967 = _GEN_2664 & _tag_way_T ? valid_35_0 : _GEN_966; // @[dcache.scala 98:{25,25}]
  wire  _GEN_968 = _GEN_2664 & way ? valid_35_1 : _GEN_967; // @[dcache.scala 98:{25,25}]
  wire  _GEN_969 = _GEN_2667 & _tag_way_T ? valid_36_0 : _GEN_968; // @[dcache.scala 98:{25,25}]
  wire  _GEN_970 = _GEN_2667 & way ? valid_36_1 : _GEN_969; // @[dcache.scala 98:{25,25}]
  wire  _GEN_971 = _GEN_2670 & _tag_way_T ? valid_37_0 : _GEN_970; // @[dcache.scala 98:{25,25}]
  wire  _GEN_972 = _GEN_2670 & way ? valid_37_1 : _GEN_971; // @[dcache.scala 98:{25,25}]
  wire  _GEN_973 = _GEN_2673 & _tag_way_T ? valid_38_0 : _GEN_972; // @[dcache.scala 98:{25,25}]
  wire  _GEN_974 = _GEN_2673 & way ? valid_38_1 : _GEN_973; // @[dcache.scala 98:{25,25}]
  wire  _GEN_975 = _GEN_2676 & _tag_way_T ? valid_39_0 : _GEN_974; // @[dcache.scala 98:{25,25}]
  wire  _GEN_976 = _GEN_2676 & way ? valid_39_1 : _GEN_975; // @[dcache.scala 98:{25,25}]
  wire  _GEN_977 = _GEN_2679 & _tag_way_T ? valid_40_0 : _GEN_976; // @[dcache.scala 98:{25,25}]
  wire  _GEN_978 = _GEN_2679 & way ? valid_40_1 : _GEN_977; // @[dcache.scala 98:{25,25}]
  wire  _GEN_979 = _GEN_2682 & _tag_way_T ? valid_41_0 : _GEN_978; // @[dcache.scala 98:{25,25}]
  wire  _GEN_980 = _GEN_2682 & way ? valid_41_1 : _GEN_979; // @[dcache.scala 98:{25,25}]
  wire  _GEN_981 = _GEN_2685 & _tag_way_T ? valid_42_0 : _GEN_980; // @[dcache.scala 98:{25,25}]
  wire  _GEN_982 = _GEN_2685 & way ? valid_42_1 : _GEN_981; // @[dcache.scala 98:{25,25}]
  wire  _GEN_983 = _GEN_2688 & _tag_way_T ? valid_43_0 : _GEN_982; // @[dcache.scala 98:{25,25}]
  wire  _GEN_984 = _GEN_2688 & way ? valid_43_1 : _GEN_983; // @[dcache.scala 98:{25,25}]
  wire  _GEN_985 = _GEN_2691 & _tag_way_T ? valid_44_0 : _GEN_984; // @[dcache.scala 98:{25,25}]
  wire  _GEN_986 = _GEN_2691 & way ? valid_44_1 : _GEN_985; // @[dcache.scala 98:{25,25}]
  wire  _GEN_987 = _GEN_2694 & _tag_way_T ? valid_45_0 : _GEN_986; // @[dcache.scala 98:{25,25}]
  wire  _GEN_988 = _GEN_2694 & way ? valid_45_1 : _GEN_987; // @[dcache.scala 98:{25,25}]
  wire  _GEN_989 = _GEN_2697 & _tag_way_T ? valid_46_0 : _GEN_988; // @[dcache.scala 98:{25,25}]
  wire  _GEN_990 = _GEN_2697 & way ? valid_46_1 : _GEN_989; // @[dcache.scala 98:{25,25}]
  wire  _GEN_991 = _GEN_2700 & _tag_way_T ? valid_47_0 : _GEN_990; // @[dcache.scala 98:{25,25}]
  wire  _GEN_992 = _GEN_2700 & way ? valid_47_1 : _GEN_991; // @[dcache.scala 98:{25,25}]
  wire  _GEN_993 = _GEN_2703 & _tag_way_T ? valid_48_0 : _GEN_992; // @[dcache.scala 98:{25,25}]
  wire  _GEN_994 = _GEN_2703 & way ? valid_48_1 : _GEN_993; // @[dcache.scala 98:{25,25}]
  wire  _GEN_995 = _GEN_2706 & _tag_way_T ? valid_49_0 : _GEN_994; // @[dcache.scala 98:{25,25}]
  wire  _GEN_996 = _GEN_2706 & way ? valid_49_1 : _GEN_995; // @[dcache.scala 98:{25,25}]
  wire  _GEN_997 = _GEN_2709 & _tag_way_T ? valid_50_0 : _GEN_996; // @[dcache.scala 98:{25,25}]
  wire  _GEN_998 = _GEN_2709 & way ? valid_50_1 : _GEN_997; // @[dcache.scala 98:{25,25}]
  wire  _GEN_999 = _GEN_2712 & _tag_way_T ? valid_51_0 : _GEN_998; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1000 = _GEN_2712 & way ? valid_51_1 : _GEN_999; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1001 = _GEN_2715 & _tag_way_T ? valid_52_0 : _GEN_1000; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1002 = _GEN_2715 & way ? valid_52_1 : _GEN_1001; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1003 = _GEN_2718 & _tag_way_T ? valid_53_0 : _GEN_1002; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1004 = _GEN_2718 & way ? valid_53_1 : _GEN_1003; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1005 = _GEN_2721 & _tag_way_T ? valid_54_0 : _GEN_1004; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1006 = _GEN_2721 & way ? valid_54_1 : _GEN_1005; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1007 = _GEN_2724 & _tag_way_T ? valid_55_0 : _GEN_1006; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1008 = _GEN_2724 & way ? valid_55_1 : _GEN_1007; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1009 = _GEN_2727 & _tag_way_T ? valid_56_0 : _GEN_1008; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1010 = _GEN_2727 & way ? valid_56_1 : _GEN_1009; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1011 = _GEN_2730 & _tag_way_T ? valid_57_0 : _GEN_1010; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1012 = _GEN_2730 & way ? valid_57_1 : _GEN_1011; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1013 = _GEN_2733 & _tag_way_T ? valid_58_0 : _GEN_1012; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1014 = _GEN_2733 & way ? valid_58_1 : _GEN_1013; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1015 = _GEN_2736 & _tag_way_T ? valid_59_0 : _GEN_1014; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1016 = _GEN_2736 & way ? valid_59_1 : _GEN_1015; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1017 = _GEN_2739 & _tag_way_T ? valid_60_0 : _GEN_1016; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1018 = _GEN_2739 & way ? valid_60_1 : _GEN_1017; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1019 = _GEN_2742 & _tag_way_T ? valid_61_0 : _GEN_1018; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1020 = _GEN_2742 & way ? valid_61_1 : _GEN_1019; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1021 = _GEN_2745 & _tag_way_T ? valid_62_0 : _GEN_1020; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1022 = _GEN_2745 & way ? valid_62_1 : _GEN_1021; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1023 = _GEN_2748 & _tag_way_T ? valid_63_0 : _GEN_1022; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1024 = _GEN_2748 & way ? valid_63_1 : _GEN_1023; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1025 = _GEN_2751 & _tag_way_T ? valid_64_0 : _GEN_1024; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1026 = _GEN_2751 & way ? valid_64_1 : _GEN_1025; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1027 = _GEN_2754 & _tag_way_T ? valid_65_0 : _GEN_1026; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1028 = _GEN_2754 & way ? valid_65_1 : _GEN_1027; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1029 = _GEN_2757 & _tag_way_T ? valid_66_0 : _GEN_1028; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1030 = _GEN_2757 & way ? valid_66_1 : _GEN_1029; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1031 = _GEN_2760 & _tag_way_T ? valid_67_0 : _GEN_1030; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1032 = _GEN_2760 & way ? valid_67_1 : _GEN_1031; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1033 = _GEN_2763 & _tag_way_T ? valid_68_0 : _GEN_1032; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1034 = _GEN_2763 & way ? valid_68_1 : _GEN_1033; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1035 = _GEN_2766 & _tag_way_T ? valid_69_0 : _GEN_1034; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1036 = _GEN_2766 & way ? valid_69_1 : _GEN_1035; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1037 = _GEN_2769 & _tag_way_T ? valid_70_0 : _GEN_1036; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1038 = _GEN_2769 & way ? valid_70_1 : _GEN_1037; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1039 = _GEN_2772 & _tag_way_T ? valid_71_0 : _GEN_1038; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1040 = _GEN_2772 & way ? valid_71_1 : _GEN_1039; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1041 = _GEN_2775 & _tag_way_T ? valid_72_0 : _GEN_1040; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1042 = _GEN_2775 & way ? valid_72_1 : _GEN_1041; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1043 = _GEN_2778 & _tag_way_T ? valid_73_0 : _GEN_1042; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1044 = _GEN_2778 & way ? valid_73_1 : _GEN_1043; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1045 = _GEN_2781 & _tag_way_T ? valid_74_0 : _GEN_1044; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1046 = _GEN_2781 & way ? valid_74_1 : _GEN_1045; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1047 = _GEN_2784 & _tag_way_T ? valid_75_0 : _GEN_1046; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1048 = _GEN_2784 & way ? valid_75_1 : _GEN_1047; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1049 = _GEN_2787 & _tag_way_T ? valid_76_0 : _GEN_1048; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1050 = _GEN_2787 & way ? valid_76_1 : _GEN_1049; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1051 = _GEN_2790 & _tag_way_T ? valid_77_0 : _GEN_1050; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1052 = _GEN_2790 & way ? valid_77_1 : _GEN_1051; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1053 = _GEN_2793 & _tag_way_T ? valid_78_0 : _GEN_1052; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1054 = _GEN_2793 & way ? valid_78_1 : _GEN_1053; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1055 = _GEN_2796 & _tag_way_T ? valid_79_0 : _GEN_1054; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1056 = _GEN_2796 & way ? valid_79_1 : _GEN_1055; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1057 = _GEN_2799 & _tag_way_T ? valid_80_0 : _GEN_1056; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1058 = _GEN_2799 & way ? valid_80_1 : _GEN_1057; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1059 = _GEN_2802 & _tag_way_T ? valid_81_0 : _GEN_1058; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1060 = _GEN_2802 & way ? valid_81_1 : _GEN_1059; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1061 = _GEN_2805 & _tag_way_T ? valid_82_0 : _GEN_1060; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1062 = _GEN_2805 & way ? valid_82_1 : _GEN_1061; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1063 = _GEN_2808 & _tag_way_T ? valid_83_0 : _GEN_1062; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1064 = _GEN_2808 & way ? valid_83_1 : _GEN_1063; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1065 = _GEN_2811 & _tag_way_T ? valid_84_0 : _GEN_1064; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1066 = _GEN_2811 & way ? valid_84_1 : _GEN_1065; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1067 = _GEN_2814 & _tag_way_T ? valid_85_0 : _GEN_1066; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1068 = _GEN_2814 & way ? valid_85_1 : _GEN_1067; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1069 = _GEN_2817 & _tag_way_T ? valid_86_0 : _GEN_1068; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1070 = _GEN_2817 & way ? valid_86_1 : _GEN_1069; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1071 = _GEN_2820 & _tag_way_T ? valid_87_0 : _GEN_1070; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1072 = _GEN_2820 & way ? valid_87_1 : _GEN_1071; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1073 = _GEN_2823 & _tag_way_T ? valid_88_0 : _GEN_1072; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1074 = _GEN_2823 & way ? valid_88_1 : _GEN_1073; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1075 = _GEN_2826 & _tag_way_T ? valid_89_0 : _GEN_1074; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1076 = _GEN_2826 & way ? valid_89_1 : _GEN_1075; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1077 = _GEN_2829 & _tag_way_T ? valid_90_0 : _GEN_1076; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1078 = _GEN_2829 & way ? valid_90_1 : _GEN_1077; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1079 = _GEN_2832 & _tag_way_T ? valid_91_0 : _GEN_1078; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1080 = _GEN_2832 & way ? valid_91_1 : _GEN_1079; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1081 = _GEN_2835 & _tag_way_T ? valid_92_0 : _GEN_1080; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1082 = _GEN_2835 & way ? valid_92_1 : _GEN_1081; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1083 = _GEN_2838 & _tag_way_T ? valid_93_0 : _GEN_1082; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1084 = _GEN_2838 & way ? valid_93_1 : _GEN_1083; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1085 = _GEN_2841 & _tag_way_T ? valid_94_0 : _GEN_1084; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1086 = _GEN_2841 & way ? valid_94_1 : _GEN_1085; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1087 = _GEN_2844 & _tag_way_T ? valid_95_0 : _GEN_1086; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1088 = _GEN_2844 & way ? valid_95_1 : _GEN_1087; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1089 = _GEN_2847 & _tag_way_T ? valid_96_0 : _GEN_1088; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1090 = _GEN_2847 & way ? valid_96_1 : _GEN_1089; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1091 = _GEN_2850 & _tag_way_T ? valid_97_0 : _GEN_1090; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1092 = _GEN_2850 & way ? valid_97_1 : _GEN_1091; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1093 = _GEN_2853 & _tag_way_T ? valid_98_0 : _GEN_1092; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1094 = _GEN_2853 & way ? valid_98_1 : _GEN_1093; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1095 = _GEN_2856 & _tag_way_T ? valid_99_0 : _GEN_1094; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1096 = _GEN_2856 & way ? valid_99_1 : _GEN_1095; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1097 = _GEN_2859 & _tag_way_T ? valid_100_0 : _GEN_1096; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1098 = _GEN_2859 & way ? valid_100_1 : _GEN_1097; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1099 = _GEN_2862 & _tag_way_T ? valid_101_0 : _GEN_1098; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1100 = _GEN_2862 & way ? valid_101_1 : _GEN_1099; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1101 = _GEN_2865 & _tag_way_T ? valid_102_0 : _GEN_1100; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1102 = _GEN_2865 & way ? valid_102_1 : _GEN_1101; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1103 = _GEN_2868 & _tag_way_T ? valid_103_0 : _GEN_1102; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1104 = _GEN_2868 & way ? valid_103_1 : _GEN_1103; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1105 = _GEN_2871 & _tag_way_T ? valid_104_0 : _GEN_1104; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1106 = _GEN_2871 & way ? valid_104_1 : _GEN_1105; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1107 = _GEN_2874 & _tag_way_T ? valid_105_0 : _GEN_1106; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1108 = _GEN_2874 & way ? valid_105_1 : _GEN_1107; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1109 = _GEN_2877 & _tag_way_T ? valid_106_0 : _GEN_1108; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1110 = _GEN_2877 & way ? valid_106_1 : _GEN_1109; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1111 = _GEN_2880 & _tag_way_T ? valid_107_0 : _GEN_1110; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1112 = _GEN_2880 & way ? valid_107_1 : _GEN_1111; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1113 = _GEN_2883 & _tag_way_T ? valid_108_0 : _GEN_1112; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1114 = _GEN_2883 & way ? valid_108_1 : _GEN_1113; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1115 = _GEN_2886 & _tag_way_T ? valid_109_0 : _GEN_1114; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1116 = _GEN_2886 & way ? valid_109_1 : _GEN_1115; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1117 = _GEN_2889 & _tag_way_T ? valid_110_0 : _GEN_1116; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1118 = _GEN_2889 & way ? valid_110_1 : _GEN_1117; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1119 = _GEN_2892 & _tag_way_T ? valid_111_0 : _GEN_1118; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1120 = _GEN_2892 & way ? valid_111_1 : _GEN_1119; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1121 = _GEN_2895 & _tag_way_T ? valid_112_0 : _GEN_1120; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1122 = _GEN_2895 & way ? valid_112_1 : _GEN_1121; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1123 = _GEN_2898 & _tag_way_T ? valid_113_0 : _GEN_1122; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1124 = _GEN_2898 & way ? valid_113_1 : _GEN_1123; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1125 = _GEN_2901 & _tag_way_T ? valid_114_0 : _GEN_1124; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1126 = _GEN_2901 & way ? valid_114_1 : _GEN_1125; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1127 = _GEN_2904 & _tag_way_T ? valid_115_0 : _GEN_1126; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1128 = _GEN_2904 & way ? valid_115_1 : _GEN_1127; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1129 = _GEN_2907 & _tag_way_T ? valid_116_0 : _GEN_1128; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1130 = _GEN_2907 & way ? valid_116_1 : _GEN_1129; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1131 = _GEN_2910 & _tag_way_T ? valid_117_0 : _GEN_1130; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1132 = _GEN_2910 & way ? valid_117_1 : _GEN_1131; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1133 = _GEN_2913 & _tag_way_T ? valid_118_0 : _GEN_1132; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1134 = _GEN_2913 & way ? valid_118_1 : _GEN_1133; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1135 = _GEN_2916 & _tag_way_T ? valid_119_0 : _GEN_1134; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1136 = _GEN_2916 & way ? valid_119_1 : _GEN_1135; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1137 = _GEN_2919 & _tag_way_T ? valid_120_0 : _GEN_1136; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1138 = _GEN_2919 & way ? valid_120_1 : _GEN_1137; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1139 = _GEN_2922 & _tag_way_T ? valid_121_0 : _GEN_1138; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1140 = _GEN_2922 & way ? valid_121_1 : _GEN_1139; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1141 = _GEN_2925 & _tag_way_T ? valid_122_0 : _GEN_1140; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1142 = _GEN_2925 & way ? valid_122_1 : _GEN_1141; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1143 = _GEN_2928 & _tag_way_T ? valid_123_0 : _GEN_1142; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1144 = _GEN_2928 & way ? valid_123_1 : _GEN_1143; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1145 = _GEN_2931 & _tag_way_T ? valid_124_0 : _GEN_1144; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1146 = _GEN_2931 & way ? valid_124_1 : _GEN_1145; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1147 = _GEN_2934 & _tag_way_T ? valid_125_0 : _GEN_1146; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1148 = _GEN_2934 & way ? valid_125_1 : _GEN_1147; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1149 = _GEN_2937 & _tag_way_T ? valid_126_0 : _GEN_1148; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1150 = _GEN_2937 & way ? valid_126_1 : _GEN_1149; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1151 = _GEN_2940 & _tag_way_T ? valid_127_0 : _GEN_1150; // @[dcache.scala 98:{25,25}]
  wire  _GEN_1152 = _GEN_2940 & way ? valid_127_1 : _GEN_1151; // @[dcache.scala 98:{25,25}]
  wire [41:0] _cache_tag_T_5 = {_GEN_127[41:21],tag}; // @[Cat.scala 33:92]
  wire [41:0] _cache_tag_T_7 = {tag,_GEN_127[20:0]}; // @[Cat.scala 33:92]
  wire  _dirty_T_2 = _miss_T_2 & wmode; // @[dcache.scala 102:52]
  wire  _dirty_T_3 = ~miss; // @[dcache.scala 102:73]
  wire  _dirty_T_4 = _miss_T_2 & wmode & ~miss; // @[dcache.scala 102:69]
  wire  _dirty_T_11 = state == 3'h3; // @[dcache.scala 103:33]
  wire  _GEN_1538 = _GEN_2561 & hit_way ? dirty_0_1 : dirty_0_0; // @[dcache.scala 103:{26,26}]
  wire  _GEN_4093 = ~hit_way; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1539 = _GEN_2562 & ~hit_way ? dirty_1_0 : _GEN_1538; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1540 = _GEN_2562 & hit_way ? dirty_1_1 : _GEN_1539; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1541 = _GEN_2565 & ~hit_way ? dirty_2_0 : _GEN_1540; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1542 = _GEN_2565 & hit_way ? dirty_2_1 : _GEN_1541; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1543 = _GEN_2568 & ~hit_way ? dirty_3_0 : _GEN_1542; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1544 = _GEN_2568 & hit_way ? dirty_3_1 : _GEN_1543; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1545 = _GEN_2571 & ~hit_way ? dirty_4_0 : _GEN_1544; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1546 = _GEN_2571 & hit_way ? dirty_4_1 : _GEN_1545; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1547 = _GEN_2574 & ~hit_way ? dirty_5_0 : _GEN_1546; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1548 = _GEN_2574 & hit_way ? dirty_5_1 : _GEN_1547; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1549 = _GEN_2577 & ~hit_way ? dirty_6_0 : _GEN_1548; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1550 = _GEN_2577 & hit_way ? dirty_6_1 : _GEN_1549; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1551 = _GEN_2580 & ~hit_way ? dirty_7_0 : _GEN_1550; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1552 = _GEN_2580 & hit_way ? dirty_7_1 : _GEN_1551; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1553 = _GEN_2583 & ~hit_way ? dirty_8_0 : _GEN_1552; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1554 = _GEN_2583 & hit_way ? dirty_8_1 : _GEN_1553; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1555 = _GEN_2586 & ~hit_way ? dirty_9_0 : _GEN_1554; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1556 = _GEN_2586 & hit_way ? dirty_9_1 : _GEN_1555; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1557 = _GEN_2589 & ~hit_way ? dirty_10_0 : _GEN_1556; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1558 = _GEN_2589 & hit_way ? dirty_10_1 : _GEN_1557; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1559 = _GEN_2592 & ~hit_way ? dirty_11_0 : _GEN_1558; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1560 = _GEN_2592 & hit_way ? dirty_11_1 : _GEN_1559; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1561 = _GEN_2595 & ~hit_way ? dirty_12_0 : _GEN_1560; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1562 = _GEN_2595 & hit_way ? dirty_12_1 : _GEN_1561; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1563 = _GEN_2598 & ~hit_way ? dirty_13_0 : _GEN_1562; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1564 = _GEN_2598 & hit_way ? dirty_13_1 : _GEN_1563; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1565 = _GEN_2601 & ~hit_way ? dirty_14_0 : _GEN_1564; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1566 = _GEN_2601 & hit_way ? dirty_14_1 : _GEN_1565; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1567 = _GEN_2604 & ~hit_way ? dirty_15_0 : _GEN_1566; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1568 = _GEN_2604 & hit_way ? dirty_15_1 : _GEN_1567; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1569 = _GEN_2607 & ~hit_way ? dirty_16_0 : _GEN_1568; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1570 = _GEN_2607 & hit_way ? dirty_16_1 : _GEN_1569; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1571 = _GEN_2610 & ~hit_way ? dirty_17_0 : _GEN_1570; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1572 = _GEN_2610 & hit_way ? dirty_17_1 : _GEN_1571; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1573 = _GEN_2613 & ~hit_way ? dirty_18_0 : _GEN_1572; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1574 = _GEN_2613 & hit_way ? dirty_18_1 : _GEN_1573; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1575 = _GEN_2616 & ~hit_way ? dirty_19_0 : _GEN_1574; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1576 = _GEN_2616 & hit_way ? dirty_19_1 : _GEN_1575; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1577 = _GEN_2619 & ~hit_way ? dirty_20_0 : _GEN_1576; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1578 = _GEN_2619 & hit_way ? dirty_20_1 : _GEN_1577; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1579 = _GEN_2622 & ~hit_way ? dirty_21_0 : _GEN_1578; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1580 = _GEN_2622 & hit_way ? dirty_21_1 : _GEN_1579; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1581 = _GEN_2625 & ~hit_way ? dirty_22_0 : _GEN_1580; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1582 = _GEN_2625 & hit_way ? dirty_22_1 : _GEN_1581; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1583 = _GEN_2628 & ~hit_way ? dirty_23_0 : _GEN_1582; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1584 = _GEN_2628 & hit_way ? dirty_23_1 : _GEN_1583; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1585 = _GEN_2631 & ~hit_way ? dirty_24_0 : _GEN_1584; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1586 = _GEN_2631 & hit_way ? dirty_24_1 : _GEN_1585; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1587 = _GEN_2634 & ~hit_way ? dirty_25_0 : _GEN_1586; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1588 = _GEN_2634 & hit_way ? dirty_25_1 : _GEN_1587; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1589 = _GEN_2637 & ~hit_way ? dirty_26_0 : _GEN_1588; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1590 = _GEN_2637 & hit_way ? dirty_26_1 : _GEN_1589; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1591 = _GEN_2640 & ~hit_way ? dirty_27_0 : _GEN_1590; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1592 = _GEN_2640 & hit_way ? dirty_27_1 : _GEN_1591; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1593 = _GEN_2643 & ~hit_way ? dirty_28_0 : _GEN_1592; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1594 = _GEN_2643 & hit_way ? dirty_28_1 : _GEN_1593; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1595 = _GEN_2646 & ~hit_way ? dirty_29_0 : _GEN_1594; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1596 = _GEN_2646 & hit_way ? dirty_29_1 : _GEN_1595; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1597 = _GEN_2649 & ~hit_way ? dirty_30_0 : _GEN_1596; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1598 = _GEN_2649 & hit_way ? dirty_30_1 : _GEN_1597; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1599 = _GEN_2652 & ~hit_way ? dirty_31_0 : _GEN_1598; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1600 = _GEN_2652 & hit_way ? dirty_31_1 : _GEN_1599; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1601 = _GEN_2655 & ~hit_way ? dirty_32_0 : _GEN_1600; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1602 = _GEN_2655 & hit_way ? dirty_32_1 : _GEN_1601; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1603 = _GEN_2658 & ~hit_way ? dirty_33_0 : _GEN_1602; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1604 = _GEN_2658 & hit_way ? dirty_33_1 : _GEN_1603; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1605 = _GEN_2661 & ~hit_way ? dirty_34_0 : _GEN_1604; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1606 = _GEN_2661 & hit_way ? dirty_34_1 : _GEN_1605; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1607 = _GEN_2664 & ~hit_way ? dirty_35_0 : _GEN_1606; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1608 = _GEN_2664 & hit_way ? dirty_35_1 : _GEN_1607; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1609 = _GEN_2667 & ~hit_way ? dirty_36_0 : _GEN_1608; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1610 = _GEN_2667 & hit_way ? dirty_36_1 : _GEN_1609; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1611 = _GEN_2670 & ~hit_way ? dirty_37_0 : _GEN_1610; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1612 = _GEN_2670 & hit_way ? dirty_37_1 : _GEN_1611; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1613 = _GEN_2673 & ~hit_way ? dirty_38_0 : _GEN_1612; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1614 = _GEN_2673 & hit_way ? dirty_38_1 : _GEN_1613; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1615 = _GEN_2676 & ~hit_way ? dirty_39_0 : _GEN_1614; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1616 = _GEN_2676 & hit_way ? dirty_39_1 : _GEN_1615; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1617 = _GEN_2679 & ~hit_way ? dirty_40_0 : _GEN_1616; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1618 = _GEN_2679 & hit_way ? dirty_40_1 : _GEN_1617; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1619 = _GEN_2682 & ~hit_way ? dirty_41_0 : _GEN_1618; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1620 = _GEN_2682 & hit_way ? dirty_41_1 : _GEN_1619; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1621 = _GEN_2685 & ~hit_way ? dirty_42_0 : _GEN_1620; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1622 = _GEN_2685 & hit_way ? dirty_42_1 : _GEN_1621; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1623 = _GEN_2688 & ~hit_way ? dirty_43_0 : _GEN_1622; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1624 = _GEN_2688 & hit_way ? dirty_43_1 : _GEN_1623; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1625 = _GEN_2691 & ~hit_way ? dirty_44_0 : _GEN_1624; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1626 = _GEN_2691 & hit_way ? dirty_44_1 : _GEN_1625; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1627 = _GEN_2694 & ~hit_way ? dirty_45_0 : _GEN_1626; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1628 = _GEN_2694 & hit_way ? dirty_45_1 : _GEN_1627; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1629 = _GEN_2697 & ~hit_way ? dirty_46_0 : _GEN_1628; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1630 = _GEN_2697 & hit_way ? dirty_46_1 : _GEN_1629; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1631 = _GEN_2700 & ~hit_way ? dirty_47_0 : _GEN_1630; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1632 = _GEN_2700 & hit_way ? dirty_47_1 : _GEN_1631; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1633 = _GEN_2703 & ~hit_way ? dirty_48_0 : _GEN_1632; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1634 = _GEN_2703 & hit_way ? dirty_48_1 : _GEN_1633; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1635 = _GEN_2706 & ~hit_way ? dirty_49_0 : _GEN_1634; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1636 = _GEN_2706 & hit_way ? dirty_49_1 : _GEN_1635; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1637 = _GEN_2709 & ~hit_way ? dirty_50_0 : _GEN_1636; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1638 = _GEN_2709 & hit_way ? dirty_50_1 : _GEN_1637; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1639 = _GEN_2712 & ~hit_way ? dirty_51_0 : _GEN_1638; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1640 = _GEN_2712 & hit_way ? dirty_51_1 : _GEN_1639; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1641 = _GEN_2715 & ~hit_way ? dirty_52_0 : _GEN_1640; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1642 = _GEN_2715 & hit_way ? dirty_52_1 : _GEN_1641; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1643 = _GEN_2718 & ~hit_way ? dirty_53_0 : _GEN_1642; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1644 = _GEN_2718 & hit_way ? dirty_53_1 : _GEN_1643; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1645 = _GEN_2721 & ~hit_way ? dirty_54_0 : _GEN_1644; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1646 = _GEN_2721 & hit_way ? dirty_54_1 : _GEN_1645; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1647 = _GEN_2724 & ~hit_way ? dirty_55_0 : _GEN_1646; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1648 = _GEN_2724 & hit_way ? dirty_55_1 : _GEN_1647; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1649 = _GEN_2727 & ~hit_way ? dirty_56_0 : _GEN_1648; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1650 = _GEN_2727 & hit_way ? dirty_56_1 : _GEN_1649; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1651 = _GEN_2730 & ~hit_way ? dirty_57_0 : _GEN_1650; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1652 = _GEN_2730 & hit_way ? dirty_57_1 : _GEN_1651; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1653 = _GEN_2733 & ~hit_way ? dirty_58_0 : _GEN_1652; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1654 = _GEN_2733 & hit_way ? dirty_58_1 : _GEN_1653; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1655 = _GEN_2736 & ~hit_way ? dirty_59_0 : _GEN_1654; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1656 = _GEN_2736 & hit_way ? dirty_59_1 : _GEN_1655; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1657 = _GEN_2739 & ~hit_way ? dirty_60_0 : _GEN_1656; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1658 = _GEN_2739 & hit_way ? dirty_60_1 : _GEN_1657; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1659 = _GEN_2742 & ~hit_way ? dirty_61_0 : _GEN_1658; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1660 = _GEN_2742 & hit_way ? dirty_61_1 : _GEN_1659; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1661 = _GEN_2745 & ~hit_way ? dirty_62_0 : _GEN_1660; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1662 = _GEN_2745 & hit_way ? dirty_62_1 : _GEN_1661; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1663 = _GEN_2748 & ~hit_way ? dirty_63_0 : _GEN_1662; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1664 = _GEN_2748 & hit_way ? dirty_63_1 : _GEN_1663; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1665 = _GEN_2751 & ~hit_way ? dirty_64_0 : _GEN_1664; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1666 = _GEN_2751 & hit_way ? dirty_64_1 : _GEN_1665; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1667 = _GEN_2754 & ~hit_way ? dirty_65_0 : _GEN_1666; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1668 = _GEN_2754 & hit_way ? dirty_65_1 : _GEN_1667; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1669 = _GEN_2757 & ~hit_way ? dirty_66_0 : _GEN_1668; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1670 = _GEN_2757 & hit_way ? dirty_66_1 : _GEN_1669; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1671 = _GEN_2760 & ~hit_way ? dirty_67_0 : _GEN_1670; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1672 = _GEN_2760 & hit_way ? dirty_67_1 : _GEN_1671; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1673 = _GEN_2763 & ~hit_way ? dirty_68_0 : _GEN_1672; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1674 = _GEN_2763 & hit_way ? dirty_68_1 : _GEN_1673; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1675 = _GEN_2766 & ~hit_way ? dirty_69_0 : _GEN_1674; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1676 = _GEN_2766 & hit_way ? dirty_69_1 : _GEN_1675; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1677 = _GEN_2769 & ~hit_way ? dirty_70_0 : _GEN_1676; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1678 = _GEN_2769 & hit_way ? dirty_70_1 : _GEN_1677; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1679 = _GEN_2772 & ~hit_way ? dirty_71_0 : _GEN_1678; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1680 = _GEN_2772 & hit_way ? dirty_71_1 : _GEN_1679; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1681 = _GEN_2775 & ~hit_way ? dirty_72_0 : _GEN_1680; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1682 = _GEN_2775 & hit_way ? dirty_72_1 : _GEN_1681; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1683 = _GEN_2778 & ~hit_way ? dirty_73_0 : _GEN_1682; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1684 = _GEN_2778 & hit_way ? dirty_73_1 : _GEN_1683; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1685 = _GEN_2781 & ~hit_way ? dirty_74_0 : _GEN_1684; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1686 = _GEN_2781 & hit_way ? dirty_74_1 : _GEN_1685; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1687 = _GEN_2784 & ~hit_way ? dirty_75_0 : _GEN_1686; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1688 = _GEN_2784 & hit_way ? dirty_75_1 : _GEN_1687; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1689 = _GEN_2787 & ~hit_way ? dirty_76_0 : _GEN_1688; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1690 = _GEN_2787 & hit_way ? dirty_76_1 : _GEN_1689; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1691 = _GEN_2790 & ~hit_way ? dirty_77_0 : _GEN_1690; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1692 = _GEN_2790 & hit_way ? dirty_77_1 : _GEN_1691; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1693 = _GEN_2793 & ~hit_way ? dirty_78_0 : _GEN_1692; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1694 = _GEN_2793 & hit_way ? dirty_78_1 : _GEN_1693; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1695 = _GEN_2796 & ~hit_way ? dirty_79_0 : _GEN_1694; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1696 = _GEN_2796 & hit_way ? dirty_79_1 : _GEN_1695; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1697 = _GEN_2799 & ~hit_way ? dirty_80_0 : _GEN_1696; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1698 = _GEN_2799 & hit_way ? dirty_80_1 : _GEN_1697; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1699 = _GEN_2802 & ~hit_way ? dirty_81_0 : _GEN_1698; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1700 = _GEN_2802 & hit_way ? dirty_81_1 : _GEN_1699; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1701 = _GEN_2805 & ~hit_way ? dirty_82_0 : _GEN_1700; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1702 = _GEN_2805 & hit_way ? dirty_82_1 : _GEN_1701; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1703 = _GEN_2808 & ~hit_way ? dirty_83_0 : _GEN_1702; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1704 = _GEN_2808 & hit_way ? dirty_83_1 : _GEN_1703; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1705 = _GEN_2811 & ~hit_way ? dirty_84_0 : _GEN_1704; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1706 = _GEN_2811 & hit_way ? dirty_84_1 : _GEN_1705; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1707 = _GEN_2814 & ~hit_way ? dirty_85_0 : _GEN_1706; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1708 = _GEN_2814 & hit_way ? dirty_85_1 : _GEN_1707; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1709 = _GEN_2817 & ~hit_way ? dirty_86_0 : _GEN_1708; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1710 = _GEN_2817 & hit_way ? dirty_86_1 : _GEN_1709; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1711 = _GEN_2820 & ~hit_way ? dirty_87_0 : _GEN_1710; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1712 = _GEN_2820 & hit_way ? dirty_87_1 : _GEN_1711; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1713 = _GEN_2823 & ~hit_way ? dirty_88_0 : _GEN_1712; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1714 = _GEN_2823 & hit_way ? dirty_88_1 : _GEN_1713; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1715 = _GEN_2826 & ~hit_way ? dirty_89_0 : _GEN_1714; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1716 = _GEN_2826 & hit_way ? dirty_89_1 : _GEN_1715; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1717 = _GEN_2829 & ~hit_way ? dirty_90_0 : _GEN_1716; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1718 = _GEN_2829 & hit_way ? dirty_90_1 : _GEN_1717; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1719 = _GEN_2832 & ~hit_way ? dirty_91_0 : _GEN_1718; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1720 = _GEN_2832 & hit_way ? dirty_91_1 : _GEN_1719; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1721 = _GEN_2835 & ~hit_way ? dirty_92_0 : _GEN_1720; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1722 = _GEN_2835 & hit_way ? dirty_92_1 : _GEN_1721; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1723 = _GEN_2838 & ~hit_way ? dirty_93_0 : _GEN_1722; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1724 = _GEN_2838 & hit_way ? dirty_93_1 : _GEN_1723; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1725 = _GEN_2841 & ~hit_way ? dirty_94_0 : _GEN_1724; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1726 = _GEN_2841 & hit_way ? dirty_94_1 : _GEN_1725; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1727 = _GEN_2844 & ~hit_way ? dirty_95_0 : _GEN_1726; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1728 = _GEN_2844 & hit_way ? dirty_95_1 : _GEN_1727; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1729 = _GEN_2847 & ~hit_way ? dirty_96_0 : _GEN_1728; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1730 = _GEN_2847 & hit_way ? dirty_96_1 : _GEN_1729; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1731 = _GEN_2850 & ~hit_way ? dirty_97_0 : _GEN_1730; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1732 = _GEN_2850 & hit_way ? dirty_97_1 : _GEN_1731; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1733 = _GEN_2853 & ~hit_way ? dirty_98_0 : _GEN_1732; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1734 = _GEN_2853 & hit_way ? dirty_98_1 : _GEN_1733; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1735 = _GEN_2856 & ~hit_way ? dirty_99_0 : _GEN_1734; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1736 = _GEN_2856 & hit_way ? dirty_99_1 : _GEN_1735; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1737 = _GEN_2859 & ~hit_way ? dirty_100_0 : _GEN_1736; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1738 = _GEN_2859 & hit_way ? dirty_100_1 : _GEN_1737; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1739 = _GEN_2862 & ~hit_way ? dirty_101_0 : _GEN_1738; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1740 = _GEN_2862 & hit_way ? dirty_101_1 : _GEN_1739; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1741 = _GEN_2865 & ~hit_way ? dirty_102_0 : _GEN_1740; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1742 = _GEN_2865 & hit_way ? dirty_102_1 : _GEN_1741; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1743 = _GEN_2868 & ~hit_way ? dirty_103_0 : _GEN_1742; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1744 = _GEN_2868 & hit_way ? dirty_103_1 : _GEN_1743; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1745 = _GEN_2871 & ~hit_way ? dirty_104_0 : _GEN_1744; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1746 = _GEN_2871 & hit_way ? dirty_104_1 : _GEN_1745; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1747 = _GEN_2874 & ~hit_way ? dirty_105_0 : _GEN_1746; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1748 = _GEN_2874 & hit_way ? dirty_105_1 : _GEN_1747; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1749 = _GEN_2877 & ~hit_way ? dirty_106_0 : _GEN_1748; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1750 = _GEN_2877 & hit_way ? dirty_106_1 : _GEN_1749; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1751 = _GEN_2880 & ~hit_way ? dirty_107_0 : _GEN_1750; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1752 = _GEN_2880 & hit_way ? dirty_107_1 : _GEN_1751; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1753 = _GEN_2883 & ~hit_way ? dirty_108_0 : _GEN_1752; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1754 = _GEN_2883 & hit_way ? dirty_108_1 : _GEN_1753; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1755 = _GEN_2886 & ~hit_way ? dirty_109_0 : _GEN_1754; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1756 = _GEN_2886 & hit_way ? dirty_109_1 : _GEN_1755; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1757 = _GEN_2889 & ~hit_way ? dirty_110_0 : _GEN_1756; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1758 = _GEN_2889 & hit_way ? dirty_110_1 : _GEN_1757; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1759 = _GEN_2892 & ~hit_way ? dirty_111_0 : _GEN_1758; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1760 = _GEN_2892 & hit_way ? dirty_111_1 : _GEN_1759; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1761 = _GEN_2895 & ~hit_way ? dirty_112_0 : _GEN_1760; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1762 = _GEN_2895 & hit_way ? dirty_112_1 : _GEN_1761; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1763 = _GEN_2898 & ~hit_way ? dirty_113_0 : _GEN_1762; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1764 = _GEN_2898 & hit_way ? dirty_113_1 : _GEN_1763; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1765 = _GEN_2901 & ~hit_way ? dirty_114_0 : _GEN_1764; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1766 = _GEN_2901 & hit_way ? dirty_114_1 : _GEN_1765; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1767 = _GEN_2904 & ~hit_way ? dirty_115_0 : _GEN_1766; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1768 = _GEN_2904 & hit_way ? dirty_115_1 : _GEN_1767; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1769 = _GEN_2907 & ~hit_way ? dirty_116_0 : _GEN_1768; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1770 = _GEN_2907 & hit_way ? dirty_116_1 : _GEN_1769; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1771 = _GEN_2910 & ~hit_way ? dirty_117_0 : _GEN_1770; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1772 = _GEN_2910 & hit_way ? dirty_117_1 : _GEN_1771; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1773 = _GEN_2913 & ~hit_way ? dirty_118_0 : _GEN_1772; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1774 = _GEN_2913 & hit_way ? dirty_118_1 : _GEN_1773; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1775 = _GEN_2916 & ~hit_way ? dirty_119_0 : _GEN_1774; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1776 = _GEN_2916 & hit_way ? dirty_119_1 : _GEN_1775; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1777 = _GEN_2919 & ~hit_way ? dirty_120_0 : _GEN_1776; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1778 = _GEN_2919 & hit_way ? dirty_120_1 : _GEN_1777; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1779 = _GEN_2922 & ~hit_way ? dirty_121_0 : _GEN_1778; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1780 = _GEN_2922 & hit_way ? dirty_121_1 : _GEN_1779; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1781 = _GEN_2925 & ~hit_way ? dirty_122_0 : _GEN_1780; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1782 = _GEN_2925 & hit_way ? dirty_122_1 : _GEN_1781; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1783 = _GEN_2928 & ~hit_way ? dirty_123_0 : _GEN_1782; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1784 = _GEN_2928 & hit_way ? dirty_123_1 : _GEN_1783; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1785 = _GEN_2931 & ~hit_way ? dirty_124_0 : _GEN_1784; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1786 = _GEN_2931 & hit_way ? dirty_124_1 : _GEN_1785; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1787 = _GEN_2934 & ~hit_way ? dirty_125_0 : _GEN_1786; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1788 = _GEN_2934 & hit_way ? dirty_125_1 : _GEN_1787; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1789 = _GEN_2937 & ~hit_way ? dirty_126_0 : _GEN_1788; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1790 = _GEN_2937 & hit_way ? dirty_126_1 : _GEN_1789; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1791 = _GEN_2940 & ~hit_way ? dirty_127_0 : _GEN_1790; // @[dcache.scala 103:{26,26}]
  wire  _GEN_1792 = _GEN_2940 & hit_way ? dirty_127_1 : _GEN_1791; // @[dcache.scala 103:{26,26}]
  wire  _dirty_T_12 = state == 3'h3 ? 1'h0 : _GEN_1792; // @[dcache.scala 103:26]
  wire  _addr_T_3 = ~io_uncache; // @[dcache.scala 105:52]
  wire  _wdata_T_1 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 52:35]
  wire  _wdata_T_2 = _rmode_T & _wdata_T_1; // @[dcache.scala 110:33]
  wire [63:0] _wstrb_map_T_8 = wstrb == 8'hff ? 64'hffffffffffffffff : 64'h0; // @[dcache.scala 123:20]
  wire [63:0] _wstrb_map_T_9 = wstrb == 8'hf ? 64'hffffffff : _wstrb_map_T_8; // @[dcache.scala 122:20]
  wire [63:0] _wstrb_map_T_10 = wstrb == 8'h3 ? 64'hffff : _wstrb_map_T_9; // @[dcache.scala 121:20]
  wire [63:0] _wstrb_map_T_11 = wstrb == 8'h1 ? 64'hff : _wstrb_map_T_10; // @[dcache.scala 120:19]
  wire [190:0] _GEN_0 = {{127'd0}, _wstrb_map_T_11}; // @[dcache.scala 123:68]
  wire [190:0] _wstrb_map_T_12 = _GEN_0 << offset; // @[dcache.scala 123:68]
  wire [190:0] _GEN_128 = {{127'd0}, wdata}; // @[dcache.scala 126:22]
  wire [190:0] _wdata_map_T = _GEN_128 << offset; // @[dcache.scala 126:22]
  wire  en_w = (_dirty_T_11 | _dirty_T_4) & _valid_T_1; // @[dcache.scala 128:92]
  wire  _io_ram_bits_BWEN_T_4 = _dirty_T_2 & _valid_T_1; // @[dcache.scala 131:66]
  wire [127:0] wstrb_map = _wstrb_map_T_12[127:0]; // @[dcache.scala 119:23 120:13]
  wire [127:0] _io_ram_bits_BWEN_T_5 = ~wstrb_map; // @[dcache.scala 131:81]
  wire [127:0] _io_ram_bits_D_T_7 = buf_ & _io_ram_bits_BWEN_T_5; // @[dcache.scala 135:41]
  wire [127:0] wdata_map = _wdata_map_T[127:0]; // @[dcache.scala 125:23 126:13]
  wire [127:0] _io_ram_bits_D_T_8 = wdata_map & wstrb_map; // @[dcache.scala 135:66]
  wire [127:0] _io_ram_bits_D_T_9 = _io_ram_bits_D_T_7 | _io_ram_bits_D_T_8; // @[dcache.scala 135:55]
  wire [127:0] _io_ram_bits_D_T_10 = wmode ? _io_ram_bits_D_T_9 : buf_; // @[dcache.scala 135:22]
  reg  rcnt; // @[dcache.scala 139:21]
  wire  _rcnt_T = rstate == 3'h0; // @[dcache.scala 140:22]
  wire [127:0] _buf_T_7 = {buf_[127:64],io_mem_r_bits_data}; // @[Cat.scala 33:92]
  wire [127:0] _buf_T_9 = {io_mem_r_bits_data,buf_[63:0]}; // @[Cat.scala 33:92]
  wire  _io_mem_ar_bits_addr_T_1 = io_uncache & _req_T; // @[dcache.scala 148:42]
  wire [34:0] _GEN_4857 = {{3'd0}, addr}; // @[dcache.scala 148:84]
  wire [34:0] _io_mem_ar_bits_addr_T_4 = _GEN_4857 & 35'h7fffffff8; // @[dcache.scala 148:84]
  wire [34:0] _io_mem_ar_bits_addr_T_5 = io_uncache & _req_T ? {{3'd0}, io_in_ar_bits_addr} : _io_mem_ar_bits_addr_T_4; // @[dcache.scala 148:29]
  wire  _io_mem_ar_bits_len_T = io_uncache ? 1'h0 : 1'h1; // @[dcache.scala 150:28]
  wire [27:0] _io_mem_aw_bits_addr_T = {tag_way, 7'h0}; // @[dcache.scala 158:70]
  wire [27:0] _GEN_4858 = {{21'd0}, idx}; // @[dcache.scala 158:85]
  wire [27:0] _io_mem_aw_bits_addr_T_1 = _io_mem_aw_bits_addr_T | _GEN_4858; // @[dcache.scala 158:85]
  wire [31:0] _io_mem_aw_bits_addr_T_2 = {_io_mem_aw_bits_addr_T_1, 4'h0}; // @[dcache.scala 158:92]
  wire  _io_mem_aw_valid_T_1 = _rmode_T & io_uncache; // @[dcache.scala 161:45]
  wire  _io_mem_aw_valid_T_5 = wstate == 3'h0; // @[dcache.scala 161:108]
  wire  _io_mem_w_bits_data_T = wstate == 3'h4; // @[dcache.scala 167:37]
  wire [63:0] _io_mem_w_bits_data_T_5 = way ? io_ram_bits_Q1[127:64] : io_ram_bits_Q0[127:64]; // @[dcache.scala 167:53]
  wire [63:0] _io_mem_w_bits_data_T_10 = way ? io_ram_bits_Q1[63:0] : io_ram_bits_Q0[63:0]; // @[dcache.scala 168:28]
  wire [63:0] _io_mem_w_bits_data_T_11 = wstate == 3'h4 ? _io_mem_w_bits_data_T_5 : _io_mem_w_bits_data_T_10; // @[dcache.scala 167:28]
  wire  _io_in_r_bits_data_T_2 = _miss_T_2 & _dirty_T_3; // @[dcache.scala 175:50]
  wire [127:0] _io_in_r_bits_data_T_3 = io_ram_bits_Q1 >> offset; // @[dcache.scala 176:54]
  wire [127:0] _io_in_r_bits_data_T_5 = io_ram_bits_Q0 >> offset; // @[dcache.scala 176:86]
  wire [63:0] _io_in_r_bits_data_T_7 = hit_way ? _io_in_r_bits_data_T_3[63:0] : _io_in_r_bits_data_T_5[63:0]; // @[dcache.scala 176:30]
  wire [127:0] _io_in_r_bits_data_T_9 = buf_ >> offset; // @[dcache.scala 177:57]
  wire [127:0] _io_in_r_bits_data_T_10 = _dirty_T_11 ? _io_in_r_bits_data_T_9 : 128'h0; // @[dcache.scala 177:30]
  wire [127:0] _io_in_r_bits_data_T_11 = _miss_T_2 & _dirty_T_3 ? {{64'd0}, _io_in_r_bits_data_T_7} :
    _io_in_r_bits_data_T_10; // @[dcache.scala 175:28]
  wire [127:0] _io_in_r_bits_data_T_12 = uncache ? {{64'd0}, io_mem_r_bits_data} : _io_in_r_bits_data_T_11; // @[dcache.scala 174:28]
  wire  _io_in_r_valid_T_4 = _io_in_r_bits_data_T_2 | _dirty_T_11; // @[dcache.scala 179:55]
  reg [31:0] hit_num; // @[dcache.scala 186:22]
  reg [31:0] inst_num; // @[dcache.scala 187:23]
  wire [31:0] _hit_num_T_4 = hit_num + 32'h1; // @[dcache.scala 189:58]
  wire [31:0] _inst_num_T_4 = inst_num + 32'h1; // @[dcache.scala 190:59]
  LFSR_8 lfsr8 ( // @[dcache.scala 65:21]
    .clock(lfsr8_clock),
    .reset(lfsr8_reset),
    .io_en(lfsr8_io_en),
    .io_out(lfsr8_io_out)
  );
  assign io_in_ar_ready = state == 3'h0; // @[dcache.scala 178:28]
  assign io_in_r_valid = (_io_in_r_bits_data_T_2 | _dirty_T_11 | _rstate_T_7 & uncache) & rmode; // @[dcache.scala 179:110]
  assign io_in_r_bits_data = _io_in_r_bits_data_T_12[63:0]; // @[dcache.scala 174:21]
  assign io_in_aw_ready = state == 3'h0; // @[dcache.scala 183:28]
  assign io_in_w_ready = state == 3'h0; // @[dcache.scala 184:27]
  assign io_in_b_valid = (_io_in_r_valid_T_4 | _wstate_T_13 & uncache) & wmode; // @[dcache.scala 182:111]
  assign io_mem_ar_valid = _io_mem_ar_bits_addr_T_1 | _rstate_T_1 & _rcnt_T; // @[dcache.scala 149:26]
  assign io_mem_ar_bits_addr = _io_mem_ar_bits_addr_T_5[31:0]; // @[dcache.scala 148:23]
  assign io_mem_ar_bits_len = {{7'd0}, _io_mem_ar_bits_len_T}; // @[dcache.scala 150:22]
  assign io_mem_r_ready = 1'h1; // @[dcache.scala 155:18]
  assign io_mem_aw_valid = _rmode_T & io_uncache & _req_T_1 | _rstate_T_1 & wstate == 3'h0 & _GEN_640; // @[dcache.scala 161:25]
  assign io_mem_aw_bits_addr = io_uncache ? io_in_aw_bits_addr : _io_mem_aw_bits_addr_T_2; // @[dcache.scala 158:30]
  assign io_mem_w_valid = _io_mem_aw_valid_T_1 & _wdata_T_1 | _rstate_T_1 & (_io_mem_aw_valid_T_5 |
    _io_mem_w_bits_data_T) & _GEN_640; // @[dcache.scala 171:24]
  assign io_mem_w_bits_data = io_uncache ? io_in_w_bits_data : _io_mem_w_bits_data_T_11; // @[dcache.scala 166:28]
  assign io_mem_w_bits_strb = io_uncache ? io_in_w_bits_strb : 8'hff; // @[dcache.scala 169:29]
  assign io_mem_w_bits_last = io_uncache & _wdata_T_1 | _io_mem_w_bits_data_T; // @[dcache.scala 170:29]
  assign io_mem_b_ready = 1'h1; // @[dcache.scala 172:18]
  assign io_ram_bits_WEN = ~en_w; // @[dcache.scala 130:21]
  assign io_ram_bits_BWEN = _dirty_T_2 & _valid_T_1 ? _io_ram_bits_BWEN_T_5 : 128'h0; // @[dcache.scala 131:25]
  assign io_ram_bits_A = _rmode_T ? io_in_ar_bits_addr[10:4] : idx; // @[dcache.scala 133:22]
  assign io_ram_bits_D = _io_ram_bits_BWEN_T_4 ? wdata_map : _io_ram_bits_D_T_10; // @[dcache.scala 134:22]
  assign io_ram_bits_WAY = hit[1] ? way : hit[0]; // @[dcache.scala 68:21]
  assign io_hitrate = {inst_num,hit_num}; // @[Cat.scala 33:92]
  assign lfsr8_clock = clock;
  assign lfsr8_reset = reset;
  assign lfsr8_io_en = hit[1] & state == 3'h1; // @[dcache.scala 64:29]
  always @(posedge clock) begin
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_0 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h0 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_0 <= _cache_tag_T_5;
        end else begin
          cache_tag_0 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_0 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_0 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_1 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_1 <= _cache_tag_T_5;
        end else begin
          cache_tag_1 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_1 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_1 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_2 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_2 <= _cache_tag_T_5;
        end else begin
          cache_tag_2 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_2 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_2 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_3 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_3 <= _cache_tag_T_5;
        end else begin
          cache_tag_3 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_3 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_3 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_4 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_4 <= _cache_tag_T_5;
        end else begin
          cache_tag_4 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_4 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_4 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_5 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_5 <= _cache_tag_T_5;
        end else begin
          cache_tag_5 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_5 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_5 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_6 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_6 <= _cache_tag_T_5;
        end else begin
          cache_tag_6 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_6 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_6 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_7 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_7 <= _cache_tag_T_5;
        end else begin
          cache_tag_7 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_7 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_7 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_8 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h8 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_8 <= _cache_tag_T_5;
        end else begin
          cache_tag_8 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_8 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_8 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_9 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h9 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_9 <= _cache_tag_T_5;
        end else begin
          cache_tag_9 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_9 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_9 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_10 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'ha == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_10 <= _cache_tag_T_5;
        end else begin
          cache_tag_10 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_10 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_10 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_11 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'hb == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_11 <= _cache_tag_T_5;
        end else begin
          cache_tag_11 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_11 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_11 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_12 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'hc == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_12 <= _cache_tag_T_5;
        end else begin
          cache_tag_12 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_12 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_12 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_13 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'hd == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_13 <= _cache_tag_T_5;
        end else begin
          cache_tag_13 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_13 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_13 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_14 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'he == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_14 <= _cache_tag_T_5;
        end else begin
          cache_tag_14 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_14 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_14 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_15 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'hf == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_15 <= _cache_tag_T_5;
        end else begin
          cache_tag_15 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_15 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_15 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_16 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h10 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_16 <= _cache_tag_T_5;
        end else begin
          cache_tag_16 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_16 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_16 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_17 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h11 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_17 <= _cache_tag_T_5;
        end else begin
          cache_tag_17 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_17 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_17 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_18 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h12 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_18 <= _cache_tag_T_5;
        end else begin
          cache_tag_18 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_18 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_18 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_19 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h13 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_19 <= _cache_tag_T_5;
        end else begin
          cache_tag_19 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_19 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_19 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_20 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h14 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_20 <= _cache_tag_T_5;
        end else begin
          cache_tag_20 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_20 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_20 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_21 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h15 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_21 <= _cache_tag_T_5;
        end else begin
          cache_tag_21 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_21 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_21 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_22 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h16 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_22 <= _cache_tag_T_5;
        end else begin
          cache_tag_22 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_22 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_22 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_23 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h17 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_23 <= _cache_tag_T_5;
        end else begin
          cache_tag_23 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_23 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_23 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_24 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h18 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_24 <= _cache_tag_T_5;
        end else begin
          cache_tag_24 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_24 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_24 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_25 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h19 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_25 <= _cache_tag_T_5;
        end else begin
          cache_tag_25 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_25 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_25 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_26 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_26 <= _cache_tag_T_5;
        end else begin
          cache_tag_26 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_26 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_26 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_27 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_27 <= _cache_tag_T_5;
        end else begin
          cache_tag_27 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_27 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_27 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_28 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_28 <= _cache_tag_T_5;
        end else begin
          cache_tag_28 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_28 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_28 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_29 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_29 <= _cache_tag_T_5;
        end else begin
          cache_tag_29 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_29 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_29 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_30 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_30 <= _cache_tag_T_5;
        end else begin
          cache_tag_30 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_30 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_30 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_31 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h1f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_31 <= _cache_tag_T_5;
        end else begin
          cache_tag_31 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_31 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_31 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_32 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h20 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_32 <= _cache_tag_T_5;
        end else begin
          cache_tag_32 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_32 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_32 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_33 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h21 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_33 <= _cache_tag_T_5;
        end else begin
          cache_tag_33 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_33 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_33 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_34 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h22 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_34 <= _cache_tag_T_5;
        end else begin
          cache_tag_34 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_34 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_34 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_35 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h23 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_35 <= _cache_tag_T_5;
        end else begin
          cache_tag_35 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_35 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_35 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_36 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h24 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_36 <= _cache_tag_T_5;
        end else begin
          cache_tag_36 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_36 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_36 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_37 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h25 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_37 <= _cache_tag_T_5;
        end else begin
          cache_tag_37 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_37 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_37 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_38 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h26 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_38 <= _cache_tag_T_5;
        end else begin
          cache_tag_38 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_38 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_38 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_39 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h27 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_39 <= _cache_tag_T_5;
        end else begin
          cache_tag_39 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_39 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_39 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_40 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h28 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_40 <= _cache_tag_T_5;
        end else begin
          cache_tag_40 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_40 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_40 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_41 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h29 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_41 <= _cache_tag_T_5;
        end else begin
          cache_tag_41 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_41 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_41 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_42 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_42 <= _cache_tag_T_5;
        end else begin
          cache_tag_42 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_42 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_42 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_43 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_43 <= _cache_tag_T_5;
        end else begin
          cache_tag_43 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_43 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_43 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_44 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_44 <= _cache_tag_T_5;
        end else begin
          cache_tag_44 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_44 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_44 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_45 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_45 <= _cache_tag_T_5;
        end else begin
          cache_tag_45 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_45 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_45 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_46 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_46 <= _cache_tag_T_5;
        end else begin
          cache_tag_46 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_46 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_46 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_47 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h2f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_47 <= _cache_tag_T_5;
        end else begin
          cache_tag_47 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_47 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_47 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_48 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h30 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_48 <= _cache_tag_T_5;
        end else begin
          cache_tag_48 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_48 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_48 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_49 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h31 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_49 <= _cache_tag_T_5;
        end else begin
          cache_tag_49 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_49 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_49 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_50 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h32 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_50 <= _cache_tag_T_5;
        end else begin
          cache_tag_50 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_50 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_50 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_51 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h33 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_51 <= _cache_tag_T_5;
        end else begin
          cache_tag_51 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_51 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_51 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_52 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h34 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_52 <= _cache_tag_T_5;
        end else begin
          cache_tag_52 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_52 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_52 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_53 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h35 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_53 <= _cache_tag_T_5;
        end else begin
          cache_tag_53 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_53 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_53 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_54 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h36 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_54 <= _cache_tag_T_5;
        end else begin
          cache_tag_54 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_54 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_54 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_55 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h37 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_55 <= _cache_tag_T_5;
        end else begin
          cache_tag_55 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_55 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_55 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_56 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h38 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_56 <= _cache_tag_T_5;
        end else begin
          cache_tag_56 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_56 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_56 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_57 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h39 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_57 <= _cache_tag_T_5;
        end else begin
          cache_tag_57 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_57 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_57 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_58 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_58 <= _cache_tag_T_5;
        end else begin
          cache_tag_58 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_58 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_58 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_59 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_59 <= _cache_tag_T_5;
        end else begin
          cache_tag_59 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_59 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_59 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_60 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_60 <= _cache_tag_T_5;
        end else begin
          cache_tag_60 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_60 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_60 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_61 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_61 <= _cache_tag_T_5;
        end else begin
          cache_tag_61 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_61 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_61 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_62 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_62 <= _cache_tag_T_5;
        end else begin
          cache_tag_62 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_62 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_62 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_63 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h3f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_63 <= _cache_tag_T_5;
        end else begin
          cache_tag_63 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_63 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_63 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_64 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h40 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_64 <= _cache_tag_T_5;
        end else begin
          cache_tag_64 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_64 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_64 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_65 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h41 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_65 <= _cache_tag_T_5;
        end else begin
          cache_tag_65 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_65 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_65 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_66 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h42 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_66 <= _cache_tag_T_5;
        end else begin
          cache_tag_66 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_66 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_66 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_67 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h43 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_67 <= _cache_tag_T_5;
        end else begin
          cache_tag_67 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_67 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_67 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_68 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h44 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_68 <= _cache_tag_T_5;
        end else begin
          cache_tag_68 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_68 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_68 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_69 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h45 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_69 <= _cache_tag_T_5;
        end else begin
          cache_tag_69 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_69 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_69 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_70 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h46 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_70 <= _cache_tag_T_5;
        end else begin
          cache_tag_70 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_70 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_70 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_71 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h47 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_71 <= _cache_tag_T_5;
        end else begin
          cache_tag_71 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_71 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_71 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_72 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h48 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_72 <= _cache_tag_T_5;
        end else begin
          cache_tag_72 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_72 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_72 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_73 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h49 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_73 <= _cache_tag_T_5;
        end else begin
          cache_tag_73 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_73 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_73 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_74 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_74 <= _cache_tag_T_5;
        end else begin
          cache_tag_74 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_74 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_74 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_75 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_75 <= _cache_tag_T_5;
        end else begin
          cache_tag_75 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_75 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_75 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_76 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_76 <= _cache_tag_T_5;
        end else begin
          cache_tag_76 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_76 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_76 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_77 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_77 <= _cache_tag_T_5;
        end else begin
          cache_tag_77 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_77 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_77 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_78 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_78 <= _cache_tag_T_5;
        end else begin
          cache_tag_78 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_78 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_78 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_79 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h4f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_79 <= _cache_tag_T_5;
        end else begin
          cache_tag_79 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_79 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_79 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_80 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h50 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_80 <= _cache_tag_T_5;
        end else begin
          cache_tag_80 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_80 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_80 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_81 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h51 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_81 <= _cache_tag_T_5;
        end else begin
          cache_tag_81 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_81 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_81 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_82 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h52 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_82 <= _cache_tag_T_5;
        end else begin
          cache_tag_82 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_82 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_82 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_83 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h53 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_83 <= _cache_tag_T_5;
        end else begin
          cache_tag_83 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_83 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_83 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_84 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h54 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_84 <= _cache_tag_T_5;
        end else begin
          cache_tag_84 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_84 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_84 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_85 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h55 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_85 <= _cache_tag_T_5;
        end else begin
          cache_tag_85 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_85 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_85 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_86 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h56 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_86 <= _cache_tag_T_5;
        end else begin
          cache_tag_86 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_86 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_86 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_87 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h57 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_87 <= _cache_tag_T_5;
        end else begin
          cache_tag_87 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_87 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_87 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_88 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h58 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_88 <= _cache_tag_T_5;
        end else begin
          cache_tag_88 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_88 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_88 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_89 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h59 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_89 <= _cache_tag_T_5;
        end else begin
          cache_tag_89 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_89 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_89 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_90 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_90 <= _cache_tag_T_5;
        end else begin
          cache_tag_90 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_90 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_90 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_91 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_91 <= _cache_tag_T_5;
        end else begin
          cache_tag_91 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_91 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_91 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_92 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_92 <= _cache_tag_T_5;
        end else begin
          cache_tag_92 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_92 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_92 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_93 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_93 <= _cache_tag_T_5;
        end else begin
          cache_tag_93 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_93 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_93 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_94 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_94 <= _cache_tag_T_5;
        end else begin
          cache_tag_94 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_94 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_94 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_95 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h5f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_95 <= _cache_tag_T_5;
        end else begin
          cache_tag_95 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_95 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_95 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_96 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h60 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_96 <= _cache_tag_T_5;
        end else begin
          cache_tag_96 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_96 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_96 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_97 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h61 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_97 <= _cache_tag_T_5;
        end else begin
          cache_tag_97 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_97 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_97 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_98 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h62 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_98 <= _cache_tag_T_5;
        end else begin
          cache_tag_98 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_98 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_98 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_99 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h63 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_99 <= _cache_tag_T_5;
        end else begin
          cache_tag_99 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_99 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_99 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_100 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h64 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_100 <= _cache_tag_T_5;
        end else begin
          cache_tag_100 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_100 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_100 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_101 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h65 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_101 <= _cache_tag_T_5;
        end else begin
          cache_tag_101 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_101 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_101 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_102 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h66 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_102 <= _cache_tag_T_5;
        end else begin
          cache_tag_102 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_102 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_102 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_103 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h67 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_103 <= _cache_tag_T_5;
        end else begin
          cache_tag_103 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_103 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_103 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_104 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h68 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_104 <= _cache_tag_T_5;
        end else begin
          cache_tag_104 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_104 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_104 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_105 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h69 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_105 <= _cache_tag_T_5;
        end else begin
          cache_tag_105 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_105 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_105 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_106 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_106 <= _cache_tag_T_5;
        end else begin
          cache_tag_106 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_106 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_106 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_107 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_107 <= _cache_tag_T_5;
        end else begin
          cache_tag_107 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_107 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_107 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_108 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_108 <= _cache_tag_T_5;
        end else begin
          cache_tag_108 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_108 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_108 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_109 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_109 <= _cache_tag_T_5;
        end else begin
          cache_tag_109 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_109 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_109 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_110 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_110 <= _cache_tag_T_5;
        end else begin
          cache_tag_110 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_110 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_110 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_111 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h6f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_111 <= _cache_tag_T_5;
        end else begin
          cache_tag_111 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_111 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_111 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_112 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h70 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_112 <= _cache_tag_T_5;
        end else begin
          cache_tag_112 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_112 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_112 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_113 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h71 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_113 <= _cache_tag_T_5;
        end else begin
          cache_tag_113 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_113 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_113 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_114 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h72 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_114 <= _cache_tag_T_5;
        end else begin
          cache_tag_114 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_114 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_114 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_115 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h73 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_115 <= _cache_tag_T_5;
        end else begin
          cache_tag_115 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_115 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_115 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_116 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h74 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_116 <= _cache_tag_T_5;
        end else begin
          cache_tag_116 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_116 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_116 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_117 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h75 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_117 <= _cache_tag_T_5;
        end else begin
          cache_tag_117 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_117 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_117 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_118 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h76 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_118 <= _cache_tag_T_5;
        end else begin
          cache_tag_118 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_118 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_118 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_119 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h77 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_119 <= _cache_tag_T_5;
        end else begin
          cache_tag_119 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_119 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_119 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_120 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h78 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_120 <= _cache_tag_T_5;
        end else begin
          cache_tag_120 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_120 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_120 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_121 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h79 == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_121 <= _cache_tag_T_5;
        end else begin
          cache_tag_121 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_121 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_121 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_122 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7a == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_122 <= _cache_tag_T_5;
        end else begin
          cache_tag_122 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_122 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_122 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_123 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7b == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_123 <= _cache_tag_T_5;
        end else begin
          cache_tag_123 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_123 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_123 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_124 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7c == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_124 <= _cache_tag_T_5;
        end else begin
          cache_tag_124 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_124 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_124 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_125 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7d == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_125 <= _cache_tag_T_5;
        end else begin
          cache_tag_125 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_125 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_125 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_126 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7e == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_126 <= _cache_tag_T_5;
        end else begin
          cache_tag_126 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[dcache.scala 61:33]
        cache_tag_126 <= cache_tag_127; // @[dcache.scala 61:33]
      end else begin
        cache_tag_126 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 29:26]
      cache_tag_127 <= 42'h0; // @[dcache.scala 29:26]
    end else if (7'h7f == idx) begin // @[dcache.scala 99:18]
      if (_valid_T_2) begin // @[dcache.scala 99:24]
        if (_tag_way_T) begin // @[dcache.scala 100:26]
          cache_tag_127 <= _cache_tag_T_5;
        end else begin
          cache_tag_127 <= _cache_tag_T_7;
        end
      end else if (!(7'h7f == idx)) begin // @[dcache.scala 61:33]
        cache_tag_127 <= _GEN_126;
      end
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_0_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2561 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_0_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_0_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2561 & way) begin // @[dcache.scala 98:19]
      valid_0_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_1_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2562 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_1_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_1_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2562 & way) begin // @[dcache.scala 98:19]
      valid_1_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_2_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2565 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_2_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_2_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2565 & way) begin // @[dcache.scala 98:19]
      valid_2_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_3_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2568 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_3_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_3_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2568 & way) begin // @[dcache.scala 98:19]
      valid_3_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_4_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2571 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_4_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_4_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2571 & way) begin // @[dcache.scala 98:19]
      valid_4_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_5_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2574 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_5_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_5_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2574 & way) begin // @[dcache.scala 98:19]
      valid_5_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_6_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2577 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_6_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_6_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2577 & way) begin // @[dcache.scala 98:19]
      valid_6_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_7_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2580 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_7_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_7_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2580 & way) begin // @[dcache.scala 98:19]
      valid_7_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_8_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2583 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_8_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_8_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2583 & way) begin // @[dcache.scala 98:19]
      valid_8_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_9_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2586 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_9_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_9_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2586 & way) begin // @[dcache.scala 98:19]
      valid_9_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_10_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2589 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_10_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_10_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2589 & way) begin // @[dcache.scala 98:19]
      valid_10_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_11_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2592 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_11_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_11_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2592 & way) begin // @[dcache.scala 98:19]
      valid_11_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_12_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2595 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_12_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_12_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2595 & way) begin // @[dcache.scala 98:19]
      valid_12_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_13_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2598 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_13_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_13_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2598 & way) begin // @[dcache.scala 98:19]
      valid_13_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_14_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2601 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_14_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_14_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2601 & way) begin // @[dcache.scala 98:19]
      valid_14_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_15_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2604 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_15_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_15_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2604 & way) begin // @[dcache.scala 98:19]
      valid_15_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_16_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2607 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_16_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_16_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2607 & way) begin // @[dcache.scala 98:19]
      valid_16_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_17_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2610 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_17_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_17_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2610 & way) begin // @[dcache.scala 98:19]
      valid_17_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_18_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2613 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_18_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_18_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2613 & way) begin // @[dcache.scala 98:19]
      valid_18_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_19_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2616 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_19_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_19_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2616 & way) begin // @[dcache.scala 98:19]
      valid_19_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_20_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2619 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_20_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_20_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2619 & way) begin // @[dcache.scala 98:19]
      valid_20_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_21_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2622 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_21_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_21_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2622 & way) begin // @[dcache.scala 98:19]
      valid_21_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_22_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2625 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_22_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_22_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2625 & way) begin // @[dcache.scala 98:19]
      valid_22_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_23_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2628 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_23_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_23_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2628 & way) begin // @[dcache.scala 98:19]
      valid_23_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_24_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2631 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_24_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_24_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2631 & way) begin // @[dcache.scala 98:19]
      valid_24_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_25_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2634 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_25_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_25_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2634 & way) begin // @[dcache.scala 98:19]
      valid_25_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_26_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2637 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_26_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_26_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2637 & way) begin // @[dcache.scala 98:19]
      valid_26_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_27_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2640 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_27_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_27_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2640 & way) begin // @[dcache.scala 98:19]
      valid_27_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_28_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2643 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_28_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_28_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2643 & way) begin // @[dcache.scala 98:19]
      valid_28_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_29_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2646 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_29_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_29_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2646 & way) begin // @[dcache.scala 98:19]
      valid_29_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_30_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2649 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_30_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_30_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2649 & way) begin // @[dcache.scala 98:19]
      valid_30_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_31_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2652 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_31_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_31_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2652 & way) begin // @[dcache.scala 98:19]
      valid_31_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_32_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2655 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_32_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_32_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2655 & way) begin // @[dcache.scala 98:19]
      valid_32_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_33_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2658 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_33_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_33_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2658 & way) begin // @[dcache.scala 98:19]
      valid_33_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_34_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2661 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_34_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_34_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2661 & way) begin // @[dcache.scala 98:19]
      valid_34_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_35_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2664 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_35_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_35_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2664 & way) begin // @[dcache.scala 98:19]
      valid_35_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_36_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2667 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_36_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_36_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2667 & way) begin // @[dcache.scala 98:19]
      valid_36_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_37_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2670 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_37_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_37_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2670 & way) begin // @[dcache.scala 98:19]
      valid_37_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_38_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2673 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_38_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_38_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2673 & way) begin // @[dcache.scala 98:19]
      valid_38_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_39_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2676 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_39_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_39_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2676 & way) begin // @[dcache.scala 98:19]
      valid_39_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_40_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2679 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_40_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_40_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2679 & way) begin // @[dcache.scala 98:19]
      valid_40_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_41_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2682 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_41_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_41_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2682 & way) begin // @[dcache.scala 98:19]
      valid_41_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_42_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2685 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_42_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_42_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2685 & way) begin // @[dcache.scala 98:19]
      valid_42_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_43_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2688 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_43_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_43_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2688 & way) begin // @[dcache.scala 98:19]
      valid_43_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_44_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2691 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_44_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_44_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2691 & way) begin // @[dcache.scala 98:19]
      valid_44_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_45_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2694 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_45_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_45_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2694 & way) begin // @[dcache.scala 98:19]
      valid_45_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_46_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2697 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_46_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_46_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2697 & way) begin // @[dcache.scala 98:19]
      valid_46_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_47_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2700 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_47_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_47_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2700 & way) begin // @[dcache.scala 98:19]
      valid_47_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_48_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2703 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_48_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_48_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2703 & way) begin // @[dcache.scala 98:19]
      valid_48_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_49_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2706 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_49_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_49_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2706 & way) begin // @[dcache.scala 98:19]
      valid_49_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_50_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2709 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_50_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_50_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2709 & way) begin // @[dcache.scala 98:19]
      valid_50_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_51_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2712 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_51_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_51_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2712 & way) begin // @[dcache.scala 98:19]
      valid_51_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_52_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2715 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_52_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_52_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2715 & way) begin // @[dcache.scala 98:19]
      valid_52_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_53_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2718 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_53_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_53_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2718 & way) begin // @[dcache.scala 98:19]
      valid_53_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_54_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2721 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_54_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_54_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2721 & way) begin // @[dcache.scala 98:19]
      valid_54_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_55_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2724 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_55_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_55_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2724 & way) begin // @[dcache.scala 98:19]
      valid_55_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_56_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2727 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_56_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_56_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2727 & way) begin // @[dcache.scala 98:19]
      valid_56_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_57_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2730 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_57_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_57_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2730 & way) begin // @[dcache.scala 98:19]
      valid_57_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_58_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2733 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_58_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_58_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2733 & way) begin // @[dcache.scala 98:19]
      valid_58_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_59_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2736 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_59_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_59_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2736 & way) begin // @[dcache.scala 98:19]
      valid_59_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_60_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2739 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_60_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_60_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2739 & way) begin // @[dcache.scala 98:19]
      valid_60_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_61_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2742 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_61_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_61_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2742 & way) begin // @[dcache.scala 98:19]
      valid_61_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_62_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2745 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_62_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_62_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2745 & way) begin // @[dcache.scala 98:19]
      valid_62_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_63_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2748 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_63_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_63_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2748 & way) begin // @[dcache.scala 98:19]
      valid_63_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_64_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2751 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_64_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_64_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2751 & way) begin // @[dcache.scala 98:19]
      valid_64_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_65_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2754 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_65_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_65_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2754 & way) begin // @[dcache.scala 98:19]
      valid_65_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_66_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2757 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_66_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_66_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2757 & way) begin // @[dcache.scala 98:19]
      valid_66_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_67_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2760 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_67_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_67_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2760 & way) begin // @[dcache.scala 98:19]
      valid_67_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_68_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2763 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_68_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_68_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2763 & way) begin // @[dcache.scala 98:19]
      valid_68_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_69_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2766 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_69_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_69_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2766 & way) begin // @[dcache.scala 98:19]
      valid_69_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_70_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2769 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_70_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_70_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2769 & way) begin // @[dcache.scala 98:19]
      valid_70_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_71_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2772 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_71_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_71_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2772 & way) begin // @[dcache.scala 98:19]
      valid_71_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_72_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2775 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_72_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_72_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2775 & way) begin // @[dcache.scala 98:19]
      valid_72_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_73_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2778 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_73_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_73_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2778 & way) begin // @[dcache.scala 98:19]
      valid_73_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_74_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2781 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_74_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_74_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2781 & way) begin // @[dcache.scala 98:19]
      valid_74_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_75_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2784 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_75_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_75_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2784 & way) begin // @[dcache.scala 98:19]
      valid_75_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_76_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2787 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_76_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_76_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2787 & way) begin // @[dcache.scala 98:19]
      valid_76_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_77_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2790 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_77_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_77_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2790 & way) begin // @[dcache.scala 98:19]
      valid_77_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_78_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2793 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_78_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_78_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2793 & way) begin // @[dcache.scala 98:19]
      valid_78_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_79_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2796 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_79_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_79_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2796 & way) begin // @[dcache.scala 98:19]
      valid_79_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_80_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2799 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_80_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_80_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2799 & way) begin // @[dcache.scala 98:19]
      valid_80_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_81_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2802 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_81_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_81_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2802 & way) begin // @[dcache.scala 98:19]
      valid_81_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_82_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2805 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_82_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_82_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2805 & way) begin // @[dcache.scala 98:19]
      valid_82_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_83_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2808 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_83_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_83_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2808 & way) begin // @[dcache.scala 98:19]
      valid_83_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_84_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2811 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_84_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_84_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2811 & way) begin // @[dcache.scala 98:19]
      valid_84_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_85_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2814 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_85_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_85_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2814 & way) begin // @[dcache.scala 98:19]
      valid_85_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_86_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2817 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_86_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_86_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2817 & way) begin // @[dcache.scala 98:19]
      valid_86_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_87_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2820 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_87_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_87_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2820 & way) begin // @[dcache.scala 98:19]
      valid_87_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_88_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2823 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_88_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_88_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2823 & way) begin // @[dcache.scala 98:19]
      valid_88_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_89_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2826 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_89_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_89_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2826 & way) begin // @[dcache.scala 98:19]
      valid_89_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_90_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2829 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_90_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_90_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2829 & way) begin // @[dcache.scala 98:19]
      valid_90_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_91_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2832 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_91_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_91_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2832 & way) begin // @[dcache.scala 98:19]
      valid_91_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_92_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2835 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_92_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_92_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2835 & way) begin // @[dcache.scala 98:19]
      valid_92_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_93_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2838 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_93_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_93_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2838 & way) begin // @[dcache.scala 98:19]
      valid_93_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_94_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2841 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_94_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_94_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2841 & way) begin // @[dcache.scala 98:19]
      valid_94_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_95_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2844 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_95_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_95_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2844 & way) begin // @[dcache.scala 98:19]
      valid_95_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_96_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2847 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_96_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_96_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2847 & way) begin // @[dcache.scala 98:19]
      valid_96_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_97_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2850 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_97_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_97_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2850 & way) begin // @[dcache.scala 98:19]
      valid_97_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_98_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2853 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_98_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_98_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2853 & way) begin // @[dcache.scala 98:19]
      valid_98_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_99_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2856 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_99_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_99_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2856 & way) begin // @[dcache.scala 98:19]
      valid_99_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_100_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2859 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_100_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_100_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2859 & way) begin // @[dcache.scala 98:19]
      valid_100_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_101_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2862 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_101_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_101_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2862 & way) begin // @[dcache.scala 98:19]
      valid_101_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_102_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2865 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_102_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_102_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2865 & way) begin // @[dcache.scala 98:19]
      valid_102_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_103_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2868 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_103_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_103_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2868 & way) begin // @[dcache.scala 98:19]
      valid_103_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_104_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2871 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_104_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_104_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2871 & way) begin // @[dcache.scala 98:19]
      valid_104_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_105_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2874 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_105_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_105_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2874 & way) begin // @[dcache.scala 98:19]
      valid_105_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_106_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2877 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_106_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_106_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2877 & way) begin // @[dcache.scala 98:19]
      valid_106_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_107_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2880 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_107_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_107_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2880 & way) begin // @[dcache.scala 98:19]
      valid_107_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_108_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2883 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_108_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_108_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2883 & way) begin // @[dcache.scala 98:19]
      valid_108_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_109_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2886 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_109_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_109_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2886 & way) begin // @[dcache.scala 98:19]
      valid_109_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_110_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2889 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_110_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_110_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2889 & way) begin // @[dcache.scala 98:19]
      valid_110_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_111_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2892 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_111_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_111_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2892 & way) begin // @[dcache.scala 98:19]
      valid_111_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_112_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2895 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_112_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_112_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2895 & way) begin // @[dcache.scala 98:19]
      valid_112_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_113_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2898 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_113_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_113_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2898 & way) begin // @[dcache.scala 98:19]
      valid_113_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_114_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2901 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_114_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_114_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2901 & way) begin // @[dcache.scala 98:19]
      valid_114_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_115_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2904 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_115_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_115_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2904 & way) begin // @[dcache.scala 98:19]
      valid_115_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_116_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2907 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_116_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_116_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2907 & way) begin // @[dcache.scala 98:19]
      valid_116_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_117_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2910 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_117_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_117_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2910 & way) begin // @[dcache.scala 98:19]
      valid_117_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_118_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2913 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_118_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_118_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2913 & way) begin // @[dcache.scala 98:19]
      valid_118_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_119_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2916 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_119_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_119_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2916 & way) begin // @[dcache.scala 98:19]
      valid_119_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_120_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2919 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_120_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_120_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2919 & way) begin // @[dcache.scala 98:19]
      valid_120_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_121_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2922 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_121_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_121_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2922 & way) begin // @[dcache.scala 98:19]
      valid_121_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_122_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2925 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_122_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_122_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2925 & way) begin // @[dcache.scala 98:19]
      valid_122_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_123_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2928 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_123_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_123_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2928 & way) begin // @[dcache.scala 98:19]
      valid_123_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_124_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2931 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_124_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_124_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2931 & way) begin // @[dcache.scala 98:19]
      valid_124_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_125_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2934 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_125_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_125_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2934 & way) begin // @[dcache.scala 98:19]
      valid_125_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_126_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2937 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_126_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_126_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2937 & way) begin // @[dcache.scala 98:19]
      valid_126_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_127_0 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2940 & _tag_way_T) begin // @[dcache.scala 98:19]
      valid_127_0 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 30:22]
      valid_127_1 <= 1'h0; // @[dcache.scala 30:22]
    end else if (_GEN_2940 & way) begin // @[dcache.scala 98:19]
      valid_127_1 <= _rstate_T_1 & ~uncache | _GEN_1152; // @[dcache.scala 98:19]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_0_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2561 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_0_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_0_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2561 & hit_way) begin // @[dcache.scala 102:23]
      dirty_0_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_1_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2562 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_1_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_1_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2562 & hit_way) begin // @[dcache.scala 102:23]
      dirty_1_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_2_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2565 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_2_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_2_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2565 & hit_way) begin // @[dcache.scala 102:23]
      dirty_2_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_3_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2568 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_3_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_3_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2568 & hit_way) begin // @[dcache.scala 102:23]
      dirty_3_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_4_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2571 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_4_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_4_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2571 & hit_way) begin // @[dcache.scala 102:23]
      dirty_4_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_5_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2574 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_5_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_5_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2574 & hit_way) begin // @[dcache.scala 102:23]
      dirty_5_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_6_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2577 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_6_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_6_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2577 & hit_way) begin // @[dcache.scala 102:23]
      dirty_6_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_7_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2580 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_7_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_7_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2580 & hit_way) begin // @[dcache.scala 102:23]
      dirty_7_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_8_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2583 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_8_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_8_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2583 & hit_way) begin // @[dcache.scala 102:23]
      dirty_8_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_9_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2586 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_9_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_9_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2586 & hit_way) begin // @[dcache.scala 102:23]
      dirty_9_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_10_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2589 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_10_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_10_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2589 & hit_way) begin // @[dcache.scala 102:23]
      dirty_10_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_11_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2592 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_11_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_11_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2592 & hit_way) begin // @[dcache.scala 102:23]
      dirty_11_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_12_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2595 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_12_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_12_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2595 & hit_way) begin // @[dcache.scala 102:23]
      dirty_12_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_13_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2598 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_13_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_13_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2598 & hit_way) begin // @[dcache.scala 102:23]
      dirty_13_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_14_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2601 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_14_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_14_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2601 & hit_way) begin // @[dcache.scala 102:23]
      dirty_14_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_15_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2604 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_15_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_15_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2604 & hit_way) begin // @[dcache.scala 102:23]
      dirty_15_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_16_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2607 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_16_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_16_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2607 & hit_way) begin // @[dcache.scala 102:23]
      dirty_16_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_17_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2610 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_17_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_17_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2610 & hit_way) begin // @[dcache.scala 102:23]
      dirty_17_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_18_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2613 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_18_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_18_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2613 & hit_way) begin // @[dcache.scala 102:23]
      dirty_18_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_19_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2616 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_19_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_19_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2616 & hit_way) begin // @[dcache.scala 102:23]
      dirty_19_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_20_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2619 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_20_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_20_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2619 & hit_way) begin // @[dcache.scala 102:23]
      dirty_20_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_21_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2622 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_21_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_21_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2622 & hit_way) begin // @[dcache.scala 102:23]
      dirty_21_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_22_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2625 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_22_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_22_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2625 & hit_way) begin // @[dcache.scala 102:23]
      dirty_22_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_23_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2628 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_23_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_23_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2628 & hit_way) begin // @[dcache.scala 102:23]
      dirty_23_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_24_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2631 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_24_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_24_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2631 & hit_way) begin // @[dcache.scala 102:23]
      dirty_24_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_25_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2634 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_25_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_25_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2634 & hit_way) begin // @[dcache.scala 102:23]
      dirty_25_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_26_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2637 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_26_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_26_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2637 & hit_way) begin // @[dcache.scala 102:23]
      dirty_26_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_27_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2640 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_27_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_27_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2640 & hit_way) begin // @[dcache.scala 102:23]
      dirty_27_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_28_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2643 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_28_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_28_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2643 & hit_way) begin // @[dcache.scala 102:23]
      dirty_28_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_29_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2646 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_29_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_29_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2646 & hit_way) begin // @[dcache.scala 102:23]
      dirty_29_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_30_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2649 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_30_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_30_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2649 & hit_way) begin // @[dcache.scala 102:23]
      dirty_30_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_31_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2652 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_31_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_31_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2652 & hit_way) begin // @[dcache.scala 102:23]
      dirty_31_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_32_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2655 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_32_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_32_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2655 & hit_way) begin // @[dcache.scala 102:23]
      dirty_32_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_33_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2658 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_33_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_33_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2658 & hit_way) begin // @[dcache.scala 102:23]
      dirty_33_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_34_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2661 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_34_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_34_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2661 & hit_way) begin // @[dcache.scala 102:23]
      dirty_34_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_35_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2664 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_35_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_35_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2664 & hit_way) begin // @[dcache.scala 102:23]
      dirty_35_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_36_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2667 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_36_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_36_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2667 & hit_way) begin // @[dcache.scala 102:23]
      dirty_36_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_37_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2670 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_37_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_37_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2670 & hit_way) begin // @[dcache.scala 102:23]
      dirty_37_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_38_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2673 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_38_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_38_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2673 & hit_way) begin // @[dcache.scala 102:23]
      dirty_38_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_39_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2676 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_39_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_39_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2676 & hit_way) begin // @[dcache.scala 102:23]
      dirty_39_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_40_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2679 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_40_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_40_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2679 & hit_way) begin // @[dcache.scala 102:23]
      dirty_40_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_41_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2682 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_41_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_41_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2682 & hit_way) begin // @[dcache.scala 102:23]
      dirty_41_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_42_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2685 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_42_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_42_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2685 & hit_way) begin // @[dcache.scala 102:23]
      dirty_42_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_43_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2688 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_43_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_43_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2688 & hit_way) begin // @[dcache.scala 102:23]
      dirty_43_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_44_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2691 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_44_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_44_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2691 & hit_way) begin // @[dcache.scala 102:23]
      dirty_44_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_45_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2694 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_45_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_45_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2694 & hit_way) begin // @[dcache.scala 102:23]
      dirty_45_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_46_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2697 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_46_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_46_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2697 & hit_way) begin // @[dcache.scala 102:23]
      dirty_46_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_47_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2700 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_47_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_47_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2700 & hit_way) begin // @[dcache.scala 102:23]
      dirty_47_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_48_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2703 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_48_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_48_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2703 & hit_way) begin // @[dcache.scala 102:23]
      dirty_48_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_49_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2706 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_49_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_49_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2706 & hit_way) begin // @[dcache.scala 102:23]
      dirty_49_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_50_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2709 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_50_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_50_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2709 & hit_way) begin // @[dcache.scala 102:23]
      dirty_50_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_51_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2712 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_51_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_51_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2712 & hit_way) begin // @[dcache.scala 102:23]
      dirty_51_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_52_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2715 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_52_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_52_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2715 & hit_way) begin // @[dcache.scala 102:23]
      dirty_52_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_53_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2718 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_53_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_53_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2718 & hit_way) begin // @[dcache.scala 102:23]
      dirty_53_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_54_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2721 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_54_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_54_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2721 & hit_way) begin // @[dcache.scala 102:23]
      dirty_54_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_55_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2724 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_55_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_55_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2724 & hit_way) begin // @[dcache.scala 102:23]
      dirty_55_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_56_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2727 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_56_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_56_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2727 & hit_way) begin // @[dcache.scala 102:23]
      dirty_56_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_57_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2730 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_57_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_57_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2730 & hit_way) begin // @[dcache.scala 102:23]
      dirty_57_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_58_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2733 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_58_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_58_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2733 & hit_way) begin // @[dcache.scala 102:23]
      dirty_58_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_59_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2736 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_59_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_59_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2736 & hit_way) begin // @[dcache.scala 102:23]
      dirty_59_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_60_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2739 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_60_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_60_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2739 & hit_way) begin // @[dcache.scala 102:23]
      dirty_60_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_61_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2742 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_61_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_61_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2742 & hit_way) begin // @[dcache.scala 102:23]
      dirty_61_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_62_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2745 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_62_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_62_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2745 & hit_way) begin // @[dcache.scala 102:23]
      dirty_62_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_63_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2748 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_63_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_63_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2748 & hit_way) begin // @[dcache.scala 102:23]
      dirty_63_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_64_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2751 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_64_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_64_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2751 & hit_way) begin // @[dcache.scala 102:23]
      dirty_64_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_65_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2754 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_65_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_65_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2754 & hit_way) begin // @[dcache.scala 102:23]
      dirty_65_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_66_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2757 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_66_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_66_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2757 & hit_way) begin // @[dcache.scala 102:23]
      dirty_66_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_67_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2760 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_67_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_67_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2760 & hit_way) begin // @[dcache.scala 102:23]
      dirty_67_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_68_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2763 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_68_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_68_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2763 & hit_way) begin // @[dcache.scala 102:23]
      dirty_68_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_69_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2766 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_69_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_69_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2766 & hit_way) begin // @[dcache.scala 102:23]
      dirty_69_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_70_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2769 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_70_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_70_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2769 & hit_way) begin // @[dcache.scala 102:23]
      dirty_70_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_71_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2772 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_71_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_71_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2772 & hit_way) begin // @[dcache.scala 102:23]
      dirty_71_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_72_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2775 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_72_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_72_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2775 & hit_way) begin // @[dcache.scala 102:23]
      dirty_72_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_73_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2778 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_73_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_73_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2778 & hit_way) begin // @[dcache.scala 102:23]
      dirty_73_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_74_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2781 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_74_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_74_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2781 & hit_way) begin // @[dcache.scala 102:23]
      dirty_74_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_75_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2784 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_75_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_75_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2784 & hit_way) begin // @[dcache.scala 102:23]
      dirty_75_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_76_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2787 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_76_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_76_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2787 & hit_way) begin // @[dcache.scala 102:23]
      dirty_76_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_77_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2790 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_77_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_77_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2790 & hit_way) begin // @[dcache.scala 102:23]
      dirty_77_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_78_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2793 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_78_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_78_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2793 & hit_way) begin // @[dcache.scala 102:23]
      dirty_78_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_79_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2796 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_79_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_79_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2796 & hit_way) begin // @[dcache.scala 102:23]
      dirty_79_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_80_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2799 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_80_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_80_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2799 & hit_way) begin // @[dcache.scala 102:23]
      dirty_80_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_81_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2802 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_81_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_81_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2802 & hit_way) begin // @[dcache.scala 102:23]
      dirty_81_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_82_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2805 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_82_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_82_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2805 & hit_way) begin // @[dcache.scala 102:23]
      dirty_82_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_83_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2808 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_83_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_83_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2808 & hit_way) begin // @[dcache.scala 102:23]
      dirty_83_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_84_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2811 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_84_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_84_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2811 & hit_way) begin // @[dcache.scala 102:23]
      dirty_84_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_85_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2814 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_85_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_85_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2814 & hit_way) begin // @[dcache.scala 102:23]
      dirty_85_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_86_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2817 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_86_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_86_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2817 & hit_way) begin // @[dcache.scala 102:23]
      dirty_86_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_87_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2820 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_87_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_87_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2820 & hit_way) begin // @[dcache.scala 102:23]
      dirty_87_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_88_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2823 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_88_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_88_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2823 & hit_way) begin // @[dcache.scala 102:23]
      dirty_88_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_89_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2826 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_89_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_89_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2826 & hit_way) begin // @[dcache.scala 102:23]
      dirty_89_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_90_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2829 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_90_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_90_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2829 & hit_way) begin // @[dcache.scala 102:23]
      dirty_90_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_91_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2832 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_91_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_91_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2832 & hit_way) begin // @[dcache.scala 102:23]
      dirty_91_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_92_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2835 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_92_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_92_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2835 & hit_way) begin // @[dcache.scala 102:23]
      dirty_92_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_93_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2838 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_93_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_93_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2838 & hit_way) begin // @[dcache.scala 102:23]
      dirty_93_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_94_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2841 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_94_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_94_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2841 & hit_way) begin // @[dcache.scala 102:23]
      dirty_94_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_95_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2844 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_95_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_95_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2844 & hit_way) begin // @[dcache.scala 102:23]
      dirty_95_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_96_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2847 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_96_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_96_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2847 & hit_way) begin // @[dcache.scala 102:23]
      dirty_96_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_97_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2850 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_97_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_97_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2850 & hit_way) begin // @[dcache.scala 102:23]
      dirty_97_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_98_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2853 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_98_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_98_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2853 & hit_way) begin // @[dcache.scala 102:23]
      dirty_98_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_99_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2856 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_99_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_99_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2856 & hit_way) begin // @[dcache.scala 102:23]
      dirty_99_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_100_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2859 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_100_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_100_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2859 & hit_way) begin // @[dcache.scala 102:23]
      dirty_100_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_101_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2862 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_101_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_101_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2862 & hit_way) begin // @[dcache.scala 102:23]
      dirty_101_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_102_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2865 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_102_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_102_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2865 & hit_way) begin // @[dcache.scala 102:23]
      dirty_102_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_103_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2868 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_103_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_103_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2868 & hit_way) begin // @[dcache.scala 102:23]
      dirty_103_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_104_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2871 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_104_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_104_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2871 & hit_way) begin // @[dcache.scala 102:23]
      dirty_104_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_105_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2874 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_105_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_105_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2874 & hit_way) begin // @[dcache.scala 102:23]
      dirty_105_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_106_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2877 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_106_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_106_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2877 & hit_way) begin // @[dcache.scala 102:23]
      dirty_106_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_107_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2880 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_107_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_107_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2880 & hit_way) begin // @[dcache.scala 102:23]
      dirty_107_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_108_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2883 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_108_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_108_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2883 & hit_way) begin // @[dcache.scala 102:23]
      dirty_108_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_109_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2886 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_109_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_109_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2886 & hit_way) begin // @[dcache.scala 102:23]
      dirty_109_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_110_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2889 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_110_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_110_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2889 & hit_way) begin // @[dcache.scala 102:23]
      dirty_110_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_111_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2892 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_111_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_111_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2892 & hit_way) begin // @[dcache.scala 102:23]
      dirty_111_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_112_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2895 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_112_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_112_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2895 & hit_way) begin // @[dcache.scala 102:23]
      dirty_112_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_113_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2898 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_113_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_113_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2898 & hit_way) begin // @[dcache.scala 102:23]
      dirty_113_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_114_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2901 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_114_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_114_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2901 & hit_way) begin // @[dcache.scala 102:23]
      dirty_114_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_115_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2904 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_115_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_115_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2904 & hit_way) begin // @[dcache.scala 102:23]
      dirty_115_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_116_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2907 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_116_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_116_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2907 & hit_way) begin // @[dcache.scala 102:23]
      dirty_116_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_117_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2910 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_117_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_117_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2910 & hit_way) begin // @[dcache.scala 102:23]
      dirty_117_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_118_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2913 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_118_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_118_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2913 & hit_way) begin // @[dcache.scala 102:23]
      dirty_118_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_119_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2916 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_119_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_119_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2916 & hit_way) begin // @[dcache.scala 102:23]
      dirty_119_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_120_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2919 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_120_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_120_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2919 & hit_way) begin // @[dcache.scala 102:23]
      dirty_120_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_121_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2922 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_121_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_121_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2922 & hit_way) begin // @[dcache.scala 102:23]
      dirty_121_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_122_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2925 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_122_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_122_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2925 & hit_way) begin // @[dcache.scala 102:23]
      dirty_122_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_123_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2928 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_123_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_123_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2928 & hit_way) begin // @[dcache.scala 102:23]
      dirty_123_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_124_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2931 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_124_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_124_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2931 & hit_way) begin // @[dcache.scala 102:23]
      dirty_124_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_125_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2934 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_125_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_125_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2934 & hit_way) begin // @[dcache.scala 102:23]
      dirty_125_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_126_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2937 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_126_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_126_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2937 & hit_way) begin // @[dcache.scala 102:23]
      dirty_126_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_127_0 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2940 & _GEN_4093) begin // @[dcache.scala 102:23]
      dirty_127_0 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 31:22]
      dirty_127_1 <= 1'h0; // @[dcache.scala 31:22]
    end else if (_GEN_2940 & hit_way) begin // @[dcache.scala 102:23]
      dirty_127_1 <= (_miss_T_2 & wmode & ~miss | _rstate_T_1 & wmode) & _valid_T_1 | _dirty_T_12; // @[dcache.scala 102:23]
    end
    if (reset) begin // @[dcache.scala 32:20]
      buf_ <= 128'h0; // @[dcache.scala 32:20]
    end else if (!(~_rstate_T_7 | uncache | io_uncache)) begin // @[dcache.scala 142:13]
      if (rcnt == addr[3]) begin // @[dcache.scala 143:13]
        buf_ <= _buf_T_7;
      end else begin
        buf_ <= _buf_T_9;
      end
    end
    if (reset) begin // @[dcache.scala 36:22]
      state <= 3'h0; // @[dcache.scala 36:22]
    end else if (3'h3 == state) begin // @[Mux.scala 81:58]
      state <= 3'h0;
    end else if (3'h2 == state) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[dcache.scala 78:22]
        state <= 3'h0;
      end else begin
        state <= _state_T_19;
      end
    end else if (3'h1 == state) begin // @[Mux.scala 81:58]
      state <= _state_T_6;
    end else begin
      state <= _state_T_22;
    end
    if (reset) begin // @[dcache.scala 37:23]
      rstate <= 3'h0; // @[dcache.scala 37:23]
    end else if (3'h6 == rstate) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[dcache.scala 86:19]
        rstate <= 3'h0;
      end else if (state != 3'h2) begin // @[dcache.scala 86:46]
        rstate <= 3'h0;
      end else begin
        rstate <= 3'h6;
      end
    end else if (3'h5 == rstate) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[dcache.scala 85:19]
        rstate <= 3'h0;
      end else begin
        rstate <= _rstate_T_12;
      end
    end else if (3'h4 == rstate) begin // @[Mux.scala 81:58]
      rstate <= _rstate_T_9;
    end else begin
      rstate <= _rstate_T_19;
    end
    if (reset) begin // @[dcache.scala 38:23]
      wstate <= 3'h0; // @[dcache.scala 38:23]
    end else if (3'h6 == wstate) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[dcache.scala 86:19]
        wstate <= 3'h0;
      end else if (state != 3'h2) begin // @[dcache.scala 86:46]
        wstate <= 3'h0;
      end else begin
        wstate <= 3'h6;
      end
    end else if (3'h5 == wstate) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[dcache.scala 92:19]
        wstate <= 3'h0;
      end else begin
        wstate <= _wstate_T_14;
      end
    end else if (3'h4 == wstate) begin // @[Mux.scala 81:58]
      wstate <= _wstate_T_11;
    end else begin
      wstate <= _wstate_T_21;
    end
    if (reset) begin // @[dcache.scala 41:21]
      addr <= 32'h0; // @[dcache.scala 41:21]
    end else if (_rmode_T_2 & ~io_uncache) begin // @[dcache.scala 105:14]
      addr <= io_in_ar_bits_addr;
    end else if (_wmode_T_2 & _addr_T_3) begin // @[dcache.scala 106:14]
      addr <= io_in_aw_bits_addr;
    end
    if (reset) begin // @[dcache.scala 42:22]
      wdata <= 64'h0; // @[dcache.scala 42:22]
    end else if (_rmode_T & _wdata_T_1) begin // @[dcache.scala 110:15]
      wdata <= io_in_w_bits_data;
    end
    if (reset) begin // @[dcache.scala 43:22]
      wstrb <= 8'h0; // @[dcache.scala 43:22]
    end else if (_wdata_T_2) begin // @[dcache.scala 111:15]
      wstrb <= io_in_w_bits_strb;
    end
    if (reset) begin // @[dcache.scala 44:24]
      uncache <= 1'h0; // @[dcache.scala 44:24]
    end else if (_rmode_T & req) begin // @[dcache.scala 108:16]
      uncache <= io_uncache;
    end
    if (reset) begin // @[dcache.scala 55:22]
      rmode <= 1'h0; // @[dcache.scala 55:22]
    end else begin
      rmode <= state == 3'h0 & _req_T | _rmode_T_4; // @[dcache.scala 57:9]
    end
    if (reset) begin // @[dcache.scala 56:22]
      wmode <= 1'h0; // @[dcache.scala 56:22]
    end else begin
      wmode <= _rmode_T & _req_T_1 | _wmode_T_4; // @[dcache.scala 58:9]
    end
    if (reset) begin // @[Reg.scala 35:20]
      way <= 1'h0; // @[Reg.scala 35:20]
    end else if (miss) begin // @[Reg.scala 36:18]
      way <= lfsr8_io_out[0]; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[dcache.scala 139:21]
      rcnt <= 1'h0; // @[dcache.scala 139:21]
    end else if (rstate == 3'h0) begin // @[dcache.scala 140:14]
      rcnt <= 1'h0;
    end else if (_rstate_T_7) begin // @[dcache.scala 140:42]
      rcnt <= rcnt + 1'h1;
    end
    if (reset) begin // @[dcache.scala 186:22]
      hit_num <= 32'h0; // @[dcache.scala 186:22]
    end else if (_io_in_r_bits_data_T_2) begin // @[dcache.scala 189:17]
      hit_num <= _hit_num_T_4;
    end
    if (reset) begin // @[dcache.scala 187:23]
      inst_num <= 32'h0; // @[dcache.scala 187:23]
    end else if (req) begin // @[dcache.scala 190:18]
      inst_num <= _inst_num_T_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cache_tag_0 = _RAND_0[41:0];
  _RAND_1 = {2{`RANDOM}};
  cache_tag_1 = _RAND_1[41:0];
  _RAND_2 = {2{`RANDOM}};
  cache_tag_2 = _RAND_2[41:0];
  _RAND_3 = {2{`RANDOM}};
  cache_tag_3 = _RAND_3[41:0];
  _RAND_4 = {2{`RANDOM}};
  cache_tag_4 = _RAND_4[41:0];
  _RAND_5 = {2{`RANDOM}};
  cache_tag_5 = _RAND_5[41:0];
  _RAND_6 = {2{`RANDOM}};
  cache_tag_6 = _RAND_6[41:0];
  _RAND_7 = {2{`RANDOM}};
  cache_tag_7 = _RAND_7[41:0];
  _RAND_8 = {2{`RANDOM}};
  cache_tag_8 = _RAND_8[41:0];
  _RAND_9 = {2{`RANDOM}};
  cache_tag_9 = _RAND_9[41:0];
  _RAND_10 = {2{`RANDOM}};
  cache_tag_10 = _RAND_10[41:0];
  _RAND_11 = {2{`RANDOM}};
  cache_tag_11 = _RAND_11[41:0];
  _RAND_12 = {2{`RANDOM}};
  cache_tag_12 = _RAND_12[41:0];
  _RAND_13 = {2{`RANDOM}};
  cache_tag_13 = _RAND_13[41:0];
  _RAND_14 = {2{`RANDOM}};
  cache_tag_14 = _RAND_14[41:0];
  _RAND_15 = {2{`RANDOM}};
  cache_tag_15 = _RAND_15[41:0];
  _RAND_16 = {2{`RANDOM}};
  cache_tag_16 = _RAND_16[41:0];
  _RAND_17 = {2{`RANDOM}};
  cache_tag_17 = _RAND_17[41:0];
  _RAND_18 = {2{`RANDOM}};
  cache_tag_18 = _RAND_18[41:0];
  _RAND_19 = {2{`RANDOM}};
  cache_tag_19 = _RAND_19[41:0];
  _RAND_20 = {2{`RANDOM}};
  cache_tag_20 = _RAND_20[41:0];
  _RAND_21 = {2{`RANDOM}};
  cache_tag_21 = _RAND_21[41:0];
  _RAND_22 = {2{`RANDOM}};
  cache_tag_22 = _RAND_22[41:0];
  _RAND_23 = {2{`RANDOM}};
  cache_tag_23 = _RAND_23[41:0];
  _RAND_24 = {2{`RANDOM}};
  cache_tag_24 = _RAND_24[41:0];
  _RAND_25 = {2{`RANDOM}};
  cache_tag_25 = _RAND_25[41:0];
  _RAND_26 = {2{`RANDOM}};
  cache_tag_26 = _RAND_26[41:0];
  _RAND_27 = {2{`RANDOM}};
  cache_tag_27 = _RAND_27[41:0];
  _RAND_28 = {2{`RANDOM}};
  cache_tag_28 = _RAND_28[41:0];
  _RAND_29 = {2{`RANDOM}};
  cache_tag_29 = _RAND_29[41:0];
  _RAND_30 = {2{`RANDOM}};
  cache_tag_30 = _RAND_30[41:0];
  _RAND_31 = {2{`RANDOM}};
  cache_tag_31 = _RAND_31[41:0];
  _RAND_32 = {2{`RANDOM}};
  cache_tag_32 = _RAND_32[41:0];
  _RAND_33 = {2{`RANDOM}};
  cache_tag_33 = _RAND_33[41:0];
  _RAND_34 = {2{`RANDOM}};
  cache_tag_34 = _RAND_34[41:0];
  _RAND_35 = {2{`RANDOM}};
  cache_tag_35 = _RAND_35[41:0];
  _RAND_36 = {2{`RANDOM}};
  cache_tag_36 = _RAND_36[41:0];
  _RAND_37 = {2{`RANDOM}};
  cache_tag_37 = _RAND_37[41:0];
  _RAND_38 = {2{`RANDOM}};
  cache_tag_38 = _RAND_38[41:0];
  _RAND_39 = {2{`RANDOM}};
  cache_tag_39 = _RAND_39[41:0];
  _RAND_40 = {2{`RANDOM}};
  cache_tag_40 = _RAND_40[41:0];
  _RAND_41 = {2{`RANDOM}};
  cache_tag_41 = _RAND_41[41:0];
  _RAND_42 = {2{`RANDOM}};
  cache_tag_42 = _RAND_42[41:0];
  _RAND_43 = {2{`RANDOM}};
  cache_tag_43 = _RAND_43[41:0];
  _RAND_44 = {2{`RANDOM}};
  cache_tag_44 = _RAND_44[41:0];
  _RAND_45 = {2{`RANDOM}};
  cache_tag_45 = _RAND_45[41:0];
  _RAND_46 = {2{`RANDOM}};
  cache_tag_46 = _RAND_46[41:0];
  _RAND_47 = {2{`RANDOM}};
  cache_tag_47 = _RAND_47[41:0];
  _RAND_48 = {2{`RANDOM}};
  cache_tag_48 = _RAND_48[41:0];
  _RAND_49 = {2{`RANDOM}};
  cache_tag_49 = _RAND_49[41:0];
  _RAND_50 = {2{`RANDOM}};
  cache_tag_50 = _RAND_50[41:0];
  _RAND_51 = {2{`RANDOM}};
  cache_tag_51 = _RAND_51[41:0];
  _RAND_52 = {2{`RANDOM}};
  cache_tag_52 = _RAND_52[41:0];
  _RAND_53 = {2{`RANDOM}};
  cache_tag_53 = _RAND_53[41:0];
  _RAND_54 = {2{`RANDOM}};
  cache_tag_54 = _RAND_54[41:0];
  _RAND_55 = {2{`RANDOM}};
  cache_tag_55 = _RAND_55[41:0];
  _RAND_56 = {2{`RANDOM}};
  cache_tag_56 = _RAND_56[41:0];
  _RAND_57 = {2{`RANDOM}};
  cache_tag_57 = _RAND_57[41:0];
  _RAND_58 = {2{`RANDOM}};
  cache_tag_58 = _RAND_58[41:0];
  _RAND_59 = {2{`RANDOM}};
  cache_tag_59 = _RAND_59[41:0];
  _RAND_60 = {2{`RANDOM}};
  cache_tag_60 = _RAND_60[41:0];
  _RAND_61 = {2{`RANDOM}};
  cache_tag_61 = _RAND_61[41:0];
  _RAND_62 = {2{`RANDOM}};
  cache_tag_62 = _RAND_62[41:0];
  _RAND_63 = {2{`RANDOM}};
  cache_tag_63 = _RAND_63[41:0];
  _RAND_64 = {2{`RANDOM}};
  cache_tag_64 = _RAND_64[41:0];
  _RAND_65 = {2{`RANDOM}};
  cache_tag_65 = _RAND_65[41:0];
  _RAND_66 = {2{`RANDOM}};
  cache_tag_66 = _RAND_66[41:0];
  _RAND_67 = {2{`RANDOM}};
  cache_tag_67 = _RAND_67[41:0];
  _RAND_68 = {2{`RANDOM}};
  cache_tag_68 = _RAND_68[41:0];
  _RAND_69 = {2{`RANDOM}};
  cache_tag_69 = _RAND_69[41:0];
  _RAND_70 = {2{`RANDOM}};
  cache_tag_70 = _RAND_70[41:0];
  _RAND_71 = {2{`RANDOM}};
  cache_tag_71 = _RAND_71[41:0];
  _RAND_72 = {2{`RANDOM}};
  cache_tag_72 = _RAND_72[41:0];
  _RAND_73 = {2{`RANDOM}};
  cache_tag_73 = _RAND_73[41:0];
  _RAND_74 = {2{`RANDOM}};
  cache_tag_74 = _RAND_74[41:0];
  _RAND_75 = {2{`RANDOM}};
  cache_tag_75 = _RAND_75[41:0];
  _RAND_76 = {2{`RANDOM}};
  cache_tag_76 = _RAND_76[41:0];
  _RAND_77 = {2{`RANDOM}};
  cache_tag_77 = _RAND_77[41:0];
  _RAND_78 = {2{`RANDOM}};
  cache_tag_78 = _RAND_78[41:0];
  _RAND_79 = {2{`RANDOM}};
  cache_tag_79 = _RAND_79[41:0];
  _RAND_80 = {2{`RANDOM}};
  cache_tag_80 = _RAND_80[41:0];
  _RAND_81 = {2{`RANDOM}};
  cache_tag_81 = _RAND_81[41:0];
  _RAND_82 = {2{`RANDOM}};
  cache_tag_82 = _RAND_82[41:0];
  _RAND_83 = {2{`RANDOM}};
  cache_tag_83 = _RAND_83[41:0];
  _RAND_84 = {2{`RANDOM}};
  cache_tag_84 = _RAND_84[41:0];
  _RAND_85 = {2{`RANDOM}};
  cache_tag_85 = _RAND_85[41:0];
  _RAND_86 = {2{`RANDOM}};
  cache_tag_86 = _RAND_86[41:0];
  _RAND_87 = {2{`RANDOM}};
  cache_tag_87 = _RAND_87[41:0];
  _RAND_88 = {2{`RANDOM}};
  cache_tag_88 = _RAND_88[41:0];
  _RAND_89 = {2{`RANDOM}};
  cache_tag_89 = _RAND_89[41:0];
  _RAND_90 = {2{`RANDOM}};
  cache_tag_90 = _RAND_90[41:0];
  _RAND_91 = {2{`RANDOM}};
  cache_tag_91 = _RAND_91[41:0];
  _RAND_92 = {2{`RANDOM}};
  cache_tag_92 = _RAND_92[41:0];
  _RAND_93 = {2{`RANDOM}};
  cache_tag_93 = _RAND_93[41:0];
  _RAND_94 = {2{`RANDOM}};
  cache_tag_94 = _RAND_94[41:0];
  _RAND_95 = {2{`RANDOM}};
  cache_tag_95 = _RAND_95[41:0];
  _RAND_96 = {2{`RANDOM}};
  cache_tag_96 = _RAND_96[41:0];
  _RAND_97 = {2{`RANDOM}};
  cache_tag_97 = _RAND_97[41:0];
  _RAND_98 = {2{`RANDOM}};
  cache_tag_98 = _RAND_98[41:0];
  _RAND_99 = {2{`RANDOM}};
  cache_tag_99 = _RAND_99[41:0];
  _RAND_100 = {2{`RANDOM}};
  cache_tag_100 = _RAND_100[41:0];
  _RAND_101 = {2{`RANDOM}};
  cache_tag_101 = _RAND_101[41:0];
  _RAND_102 = {2{`RANDOM}};
  cache_tag_102 = _RAND_102[41:0];
  _RAND_103 = {2{`RANDOM}};
  cache_tag_103 = _RAND_103[41:0];
  _RAND_104 = {2{`RANDOM}};
  cache_tag_104 = _RAND_104[41:0];
  _RAND_105 = {2{`RANDOM}};
  cache_tag_105 = _RAND_105[41:0];
  _RAND_106 = {2{`RANDOM}};
  cache_tag_106 = _RAND_106[41:0];
  _RAND_107 = {2{`RANDOM}};
  cache_tag_107 = _RAND_107[41:0];
  _RAND_108 = {2{`RANDOM}};
  cache_tag_108 = _RAND_108[41:0];
  _RAND_109 = {2{`RANDOM}};
  cache_tag_109 = _RAND_109[41:0];
  _RAND_110 = {2{`RANDOM}};
  cache_tag_110 = _RAND_110[41:0];
  _RAND_111 = {2{`RANDOM}};
  cache_tag_111 = _RAND_111[41:0];
  _RAND_112 = {2{`RANDOM}};
  cache_tag_112 = _RAND_112[41:0];
  _RAND_113 = {2{`RANDOM}};
  cache_tag_113 = _RAND_113[41:0];
  _RAND_114 = {2{`RANDOM}};
  cache_tag_114 = _RAND_114[41:0];
  _RAND_115 = {2{`RANDOM}};
  cache_tag_115 = _RAND_115[41:0];
  _RAND_116 = {2{`RANDOM}};
  cache_tag_116 = _RAND_116[41:0];
  _RAND_117 = {2{`RANDOM}};
  cache_tag_117 = _RAND_117[41:0];
  _RAND_118 = {2{`RANDOM}};
  cache_tag_118 = _RAND_118[41:0];
  _RAND_119 = {2{`RANDOM}};
  cache_tag_119 = _RAND_119[41:0];
  _RAND_120 = {2{`RANDOM}};
  cache_tag_120 = _RAND_120[41:0];
  _RAND_121 = {2{`RANDOM}};
  cache_tag_121 = _RAND_121[41:0];
  _RAND_122 = {2{`RANDOM}};
  cache_tag_122 = _RAND_122[41:0];
  _RAND_123 = {2{`RANDOM}};
  cache_tag_123 = _RAND_123[41:0];
  _RAND_124 = {2{`RANDOM}};
  cache_tag_124 = _RAND_124[41:0];
  _RAND_125 = {2{`RANDOM}};
  cache_tag_125 = _RAND_125[41:0];
  _RAND_126 = {2{`RANDOM}};
  cache_tag_126 = _RAND_126[41:0];
  _RAND_127 = {2{`RANDOM}};
  cache_tag_127 = _RAND_127[41:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_1_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_1_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_2_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_2_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_3_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_3_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_4_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_4_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_5_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_5_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_6_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_6_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_7_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_7_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_8_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_8_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_9_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_9_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_10_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_10_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_11_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_11_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_12_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_12_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_13_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_13_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_14_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_14_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_15_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_15_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_16_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_16_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_17_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_17_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_18_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_18_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_19_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_19_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_20_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_20_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_21_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_21_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_22_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_22_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_23_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_23_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_24_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_24_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_25_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_25_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_26_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_26_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_27_0 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_27_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_28_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_28_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_29_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_29_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_30_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_30_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_31_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_31_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_32_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_32_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_33_0 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_33_1 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_34_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_34_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_35_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_35_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_36_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_36_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_37_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_37_1 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_38_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_38_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_39_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_39_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_40_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_40_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_41_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_41_1 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_42_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_42_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_43_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_43_1 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_44_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_44_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_45_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_45_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_46_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_46_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_47_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_47_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_48_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_48_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_49_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_49_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_50_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_50_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_51_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_51_1 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_52_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_52_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_53_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_53_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_54_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_54_1 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_55_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_55_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_56_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_56_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_57_0 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_57_1 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_58_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_58_1 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_59_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_59_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_60_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_60_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_61_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_61_1 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_62_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_62_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_63_0 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_63_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_64_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_64_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_65_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_65_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_66_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_66_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_67_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_67_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_68_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_68_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_69_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_69_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_70_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_70_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_71_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_71_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_72_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_72_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_73_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_73_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_74_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_74_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_75_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_75_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_76_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_76_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_77_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_77_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_78_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_78_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_79_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_79_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_80_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_80_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_81_0 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_81_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_82_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_82_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_83_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_83_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_84_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_84_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_85_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_85_1 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_86_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_86_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_87_0 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_87_1 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_88_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_88_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_89_0 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_89_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_90_0 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_90_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_91_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_91_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_92_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_92_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_93_0 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_93_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_94_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_94_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_95_0 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_95_1 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_96_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_96_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_97_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_97_1 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_98_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_98_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_99_0 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_99_1 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_100_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_100_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_101_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_101_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_102_0 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_102_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_103_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_103_1 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_104_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_104_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_105_0 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_105_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_106_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_106_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_107_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_107_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_108_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_108_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_109_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_109_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_110_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_110_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_111_0 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_111_1 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_112_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_112_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_113_0 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_113_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_114_0 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_114_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_115_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_115_1 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_116_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_116_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_117_0 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_117_1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_118_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_118_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_119_0 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_119_1 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_120_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_120_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_121_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_121_1 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_122_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_122_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_123_0 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_123_1 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_124_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_124_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_125_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_125_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_126_0 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_126_1 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_127_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127_1 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  dirty_0_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  dirty_0_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dirty_1_0 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  dirty_1_1 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  dirty_2_0 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dirty_2_1 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  dirty_3_0 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  dirty_3_1 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dirty_4_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  dirty_4_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  dirty_5_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dirty_5_1 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  dirty_6_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  dirty_6_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dirty_7_0 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  dirty_7_1 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  dirty_8_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dirty_8_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  dirty_9_0 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  dirty_9_1 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dirty_10_0 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  dirty_10_1 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  dirty_11_0 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dirty_11_1 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  dirty_12_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  dirty_12_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dirty_13_0 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  dirty_13_1 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  dirty_14_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dirty_14_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  dirty_15_0 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  dirty_15_1 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dirty_16_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  dirty_16_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  dirty_17_0 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dirty_17_1 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  dirty_18_0 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  dirty_18_1 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dirty_19_0 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  dirty_19_1 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  dirty_20_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dirty_20_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  dirty_21_0 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  dirty_21_1 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dirty_22_0 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  dirty_22_1 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  dirty_23_0 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dirty_23_1 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  dirty_24_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  dirty_24_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dirty_25_0 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  dirty_25_1 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  dirty_26_0 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dirty_26_1 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  dirty_27_0 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  dirty_27_1 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dirty_28_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  dirty_28_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  dirty_29_0 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dirty_29_1 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  dirty_30_0 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  dirty_30_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dirty_31_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  dirty_31_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  dirty_32_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dirty_32_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  dirty_33_0 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  dirty_33_1 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dirty_34_0 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  dirty_34_1 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  dirty_35_0 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dirty_35_1 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  dirty_36_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  dirty_36_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dirty_37_0 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  dirty_37_1 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  dirty_38_0 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dirty_38_1 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  dirty_39_0 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  dirty_39_1 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dirty_40_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  dirty_40_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  dirty_41_0 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dirty_41_1 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  dirty_42_0 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  dirty_42_1 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dirty_43_0 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  dirty_43_1 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  dirty_44_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dirty_44_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  dirty_45_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  dirty_45_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dirty_46_0 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  dirty_46_1 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  dirty_47_0 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dirty_47_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  dirty_48_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  dirty_48_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dirty_49_0 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  dirty_49_1 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  dirty_50_0 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dirty_50_1 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  dirty_51_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  dirty_51_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dirty_52_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  dirty_52_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  dirty_53_0 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dirty_53_1 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  dirty_54_0 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  dirty_54_1 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dirty_55_0 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  dirty_55_1 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  dirty_56_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dirty_56_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  dirty_57_0 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  dirty_57_1 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dirty_58_0 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  dirty_58_1 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  dirty_59_0 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dirty_59_1 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  dirty_60_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  dirty_60_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dirty_61_0 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  dirty_61_1 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  dirty_62_0 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dirty_62_1 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  dirty_63_0 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  dirty_63_1 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_64_0 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_64_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_65_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  dirty_65_1 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  dirty_66_0 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  dirty_66_1 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  dirty_67_0 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  dirty_67_1 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  dirty_68_0 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  dirty_68_1 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  dirty_69_0 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  dirty_69_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dirty_70_0 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  dirty_70_1 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  dirty_71_0 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dirty_71_1 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  dirty_72_0 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  dirty_72_1 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dirty_73_0 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  dirty_73_1 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  dirty_74_0 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dirty_74_1 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  dirty_75_0 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  dirty_75_1 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dirty_76_0 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  dirty_76_1 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  dirty_77_0 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dirty_77_1 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  dirty_78_0 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  dirty_78_1 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dirty_79_0 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  dirty_79_1 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  dirty_80_0 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dirty_80_1 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  dirty_81_0 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  dirty_81_1 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dirty_82_0 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  dirty_82_1 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  dirty_83_0 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dirty_83_1 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  dirty_84_0 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  dirty_84_1 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dirty_85_0 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  dirty_85_1 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  dirty_86_0 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dirty_86_1 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  dirty_87_0 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  dirty_87_1 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dirty_88_0 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  dirty_88_1 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  dirty_89_0 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dirty_89_1 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  dirty_90_0 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  dirty_90_1 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dirty_91_0 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  dirty_91_1 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  dirty_92_0 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dirty_92_1 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  dirty_93_0 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  dirty_93_1 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dirty_94_0 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  dirty_94_1 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  dirty_95_0 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dirty_95_1 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  dirty_96_0 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  dirty_96_1 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dirty_97_0 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  dirty_97_1 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  dirty_98_0 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dirty_98_1 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  dirty_99_0 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  dirty_99_1 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dirty_100_0 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  dirty_100_1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  dirty_101_0 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dirty_101_1 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  dirty_102_0 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  dirty_102_1 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dirty_103_0 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  dirty_103_1 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  dirty_104_0 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dirty_104_1 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  dirty_105_0 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  dirty_105_1 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dirty_106_0 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  dirty_106_1 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  dirty_107_0 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dirty_107_1 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  dirty_108_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  dirty_108_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dirty_109_0 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  dirty_109_1 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  dirty_110_0 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dirty_110_1 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  dirty_111_0 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  dirty_111_1 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dirty_112_0 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  dirty_112_1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  dirty_113_0 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dirty_113_1 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  dirty_114_0 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  dirty_114_1 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dirty_115_0 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  dirty_115_1 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  dirty_116_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dirty_116_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  dirty_117_0 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  dirty_117_1 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dirty_118_0 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  dirty_118_1 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  dirty_119_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dirty_119_1 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  dirty_120_0 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  dirty_120_1 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dirty_121_0 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  dirty_121_1 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  dirty_122_0 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dirty_122_1 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  dirty_123_0 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  dirty_123_1 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dirty_124_0 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  dirty_124_1 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  dirty_125_0 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dirty_125_1 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  dirty_126_0 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  dirty_126_1 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dirty_127_0 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  dirty_127_1 = _RAND_639[0:0];
  _RAND_640 = {4{`RANDOM}};
  buf_ = _RAND_640[127:0];
  _RAND_641 = {1{`RANDOM}};
  state = _RAND_641[2:0];
  _RAND_642 = {1{`RANDOM}};
  rstate = _RAND_642[2:0];
  _RAND_643 = {1{`RANDOM}};
  wstate = _RAND_643[2:0];
  _RAND_644 = {1{`RANDOM}};
  addr = _RAND_644[31:0];
  _RAND_645 = {2{`RANDOM}};
  wdata = _RAND_645[63:0];
  _RAND_646 = {1{`RANDOM}};
  wstrb = _RAND_646[7:0];
  _RAND_647 = {1{`RANDOM}};
  uncache = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  rmode = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  wmode = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  way = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  rcnt = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  hit_num = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  inst_num = _RAND_653[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
