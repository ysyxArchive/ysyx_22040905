module ps2_keyboard(
  input        clock,
  input        io_ps2_clk,
  input        io_ps2_data,
  input        io_nextdata_n,
  output [7:0] io_data,
  output       io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg  rea; // @[ps2.scala 122:16]
  reg  buffer_0; // @[ps2.scala 130:19]
  reg  buffer_1; // @[ps2.scala 130:19]
  reg  buffer_2; // @[ps2.scala 130:19]
  reg  buffer_3; // @[ps2.scala 130:19]
  reg  buffer_4; // @[ps2.scala 130:19]
  reg  buffer_5; // @[ps2.scala 130:19]
  reg  buffer_6; // @[ps2.scala 130:19]
  reg  buffer_7; // @[ps2.scala 130:19]
  reg  buffer_8; // @[ps2.scala 130:19]
  reg  buffer_9; // @[ps2.scala 130:19]
  reg [7:0] fifo_0; // @[ps2.scala 131:17]
  reg [7:0] fifo_1; // @[ps2.scala 131:17]
  reg [7:0] fifo_2; // @[ps2.scala 131:17]
  reg [7:0] fifo_3; // @[ps2.scala 131:17]
  reg [7:0] fifo_4; // @[ps2.scala 131:17]
  reg [7:0] fifo_5; // @[ps2.scala 131:17]
  reg [7:0] fifo_6; // @[ps2.scala 131:17]
  reg [7:0] fifo_7; // @[ps2.scala 131:17]
  reg [2:0] w_ptr; // @[ps2.scala 132:18]
  reg [2:0] r_ptr; // @[ps2.scala 133:18]
  reg [3:0] count; // @[ps2.scala 134:18]
  reg [2:0] ps2_clk_sync; // @[ps2.scala 135:25]
  wire [1:0] ps2_clk_sync_hi = ps2_clk_sync[1:0]; // @[ps2.scala 137:35]
  wire  sampling = ps2_clk_sync[2] & ~ps2_clk_sync[1]; // @[ps2.scala 139:30]
  wire [2:0] _r_ptr_T_1 = r_ptr + 3'h1; // @[ps2.scala 149:29]
  wire  _GEN_0 = w_ptr == _r_ptr_T_1 ? 1'h0 : rea; // @[ps2.scala 150:42 ps2.scala 151:24 ps2.scala 122:16]
  wire  _GEN_3 = ~io_nextdata_n ? _GEN_0 : rea; // @[ps2.scala 148:38 ps2.scala 122:16]
  wire  _GEN_6 = rea ? _GEN_3 : rea; // @[ps2.scala 147:24 ps2.scala 122:16]
  wire [7:0] _fifo_T = {buffer_8,buffer_7,buffer_6,buffer_5,buffer_4,buffer_3,buffer_2,buffer_1}; // @[Cat.scala 30:58]
  wire [2:0] _w_ptr_T_1 = w_ptr + 3'h1; // @[ps2.scala 160:33]
  wire  _GEN_25 = ~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3
     ^ buffer_2 ^ buffer_1) | _GEN_6; // @[ps2.scala 158:162 ps2.scala 161:24]
  wire [3:0] _count_T_1 = count + 4'h1; // @[ps2.scala 167:29]
  wire [7:0] _GEN_106 = 3'h1 == r_ptr ? fifo_1 : fifo_0; // @[ps2.scala 171:12 ps2.scala 171:12]
  wire [7:0] _GEN_107 = 3'h2 == r_ptr ? fifo_2 : _GEN_106; // @[ps2.scala 171:12 ps2.scala 171:12]
  wire [7:0] _GEN_108 = 3'h3 == r_ptr ? fifo_3 : _GEN_107; // @[ps2.scala 171:12 ps2.scala 171:12]
  wire [7:0] _GEN_109 = 3'h4 == r_ptr ? fifo_4 : _GEN_108; // @[ps2.scala 171:12 ps2.scala 171:12]
  wire [7:0] _GEN_110 = 3'h5 == r_ptr ? fifo_5 : _GEN_109; // @[ps2.scala 171:12 ps2.scala 171:12]
  wire [7:0] _GEN_111 = 3'h6 == r_ptr ? fifo_6 : _GEN_110; // @[ps2.scala 171:12 ps2.scala 171:12]
  assign io_data = 3'h7 == r_ptr ? fifo_7 : _GEN_111; // @[ps2.scala 171:12 ps2.scala 171:12]
  assign io_ready = rea; // @[ps2.scala 140:24 ps2.scala 128:13]
  always @(posedge clock) begin
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        rea <= _GEN_25;
      end else begin
        rea <= _GEN_6;
      end
    end else begin
      rea <= _GEN_6;
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h0 == count) begin // @[ps2.scala 166:30]
          buffer_0 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h1 == count) begin // @[ps2.scala 166:30]
          buffer_1 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h2 == count) begin // @[ps2.scala 166:30]
          buffer_2 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h3 == count) begin // @[ps2.scala 166:30]
          buffer_3 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h4 == count) begin // @[ps2.scala 166:30]
          buffer_4 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h5 == count) begin // @[ps2.scala 166:30]
          buffer_5 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h6 == count) begin // @[ps2.scala 166:30]
          buffer_6 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h7 == count) begin // @[ps2.scala 166:30]
          buffer_7 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h8 == count) begin // @[ps2.scala 166:30]
          buffer_8 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (!(count == 4'ha)) begin // @[ps2.scala 157:31]
        if (4'h9 == count) begin // @[ps2.scala 166:30]
          buffer_9 <= io_ps2_data; // @[ps2.scala 166:30]
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h0 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_0 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h1 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_1 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h2 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_2 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h3 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_3 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h4 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_4 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h5 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_5 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h6 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_6 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          if (3'h7 == w_ptr) begin // @[ps2.scala 159:32]
            fifo_7 <= _fifo_T; // @[ps2.scala 159:32]
          end
        end
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        if (~buffer_0 & io_ps2_data & (buffer_9 ^ buffer_8 ^ buffer_7 ^ buffer_6 ^ buffer_5 ^ buffer_4 ^ buffer_3 ^
          buffer_2 ^ buffer_1)) begin // @[ps2.scala 158:162]
          w_ptr <= _w_ptr_T_1; // @[ps2.scala 160:26]
        end
      end
    end
    if (rea) begin // @[ps2.scala 147:24]
      if (~io_nextdata_n) begin // @[ps2.scala 148:38]
        r_ptr <= _r_ptr_T_1; // @[ps2.scala 149:22]
      end
    end
    if (sampling) begin // @[ps2.scala 156:29]
      if (count == 4'ha) begin // @[ps2.scala 157:31]
        count <= 4'h0; // @[ps2.scala 164:22]
      end else begin
        count <= _count_T_1; // @[ps2.scala 167:22]
      end
    end
    ps2_clk_sync <= {ps2_clk_sync_hi,io_ps2_clk}; // @[Cat.scala 30:58]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rea = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buffer_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  buffer_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  buffer_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buffer_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  buffer_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  fifo_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  fifo_1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  fifo_2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  fifo_3 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  fifo_4 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  fifo_5 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  fifo_6 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  fifo_7 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  w_ptr = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  r_ptr = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  count = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  ps2_clk_sync = _RAND_22[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ps2ascii(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [255:0] _GEN_21 = 8'h15 == io_in ? 256'h71 : 256'h0; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_22 = 8'h16 == io_in ? 256'h31 : _GEN_21; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_23 = 8'h17 == io_in ? 256'h0 : _GEN_22; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_24 = 8'h18 == io_in ? 256'h0 : _GEN_23; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_25 = 8'h19 == io_in ? 256'h0 : _GEN_24; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_26 = 8'h1a == io_in ? 256'h7a : _GEN_25; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_27 = 8'h1b == io_in ? 256'h73 : _GEN_26; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_28 = 8'h1c == io_in ? 256'h61 : _GEN_27; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_29 = 8'h1d == io_in ? 256'h77 : _GEN_28; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_30 = 8'h1e == io_in ? 256'h32 : _GEN_29; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_31 = 8'h1f == io_in ? 256'h0 : _GEN_30; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_32 = 8'h20 == io_in ? 256'h0 : _GEN_31; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_33 = 8'h21 == io_in ? 256'h63 : _GEN_32; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_34 = 8'h22 == io_in ? 256'h78 : _GEN_33; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_35 = 8'h23 == io_in ? 256'h64 : _GEN_34; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_36 = 8'h24 == io_in ? 256'h65 : _GEN_35; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_37 = 8'h25 == io_in ? 256'h34 : _GEN_36; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_38 = 8'h26 == io_in ? 256'h33 : _GEN_37; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_39 = 8'h27 == io_in ? 256'h0 : _GEN_38; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_40 = 8'h28 == io_in ? 256'h0 : _GEN_39; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_41 = 8'h29 == io_in ? 256'h0 : _GEN_40; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_42 = 8'h2a == io_in ? 256'h76 : _GEN_41; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_43 = 8'h2b == io_in ? 256'h66 : _GEN_42; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_44 = 8'h2c == io_in ? 256'h74 : _GEN_43; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_45 = 8'h2d == io_in ? 256'h72 : _GEN_44; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_46 = 8'h2e == io_in ? 256'h35 : _GEN_45; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_47 = 8'h2f == io_in ? 256'h0 : _GEN_46; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_48 = 8'h30 == io_in ? 256'h0 : _GEN_47; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_49 = 8'h31 == io_in ? 256'h6e : _GEN_48; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_50 = 8'h32 == io_in ? 256'h62 : _GEN_49; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_51 = 8'h33 == io_in ? 256'h68 : _GEN_50; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_52 = 8'h34 == io_in ? 256'h67 : _GEN_51; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_53 = 8'h35 == io_in ? 256'h79 : _GEN_52; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_54 = 8'h36 == io_in ? 256'h36 : _GEN_53; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_55 = 8'h37 == io_in ? 256'h0 : _GEN_54; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_56 = 8'h38 == io_in ? 256'h0 : _GEN_55; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_57 = 8'h39 == io_in ? 256'h0 : _GEN_56; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_58 = 8'h3a == io_in ? 256'h6d : _GEN_57; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_59 = 8'h3b == io_in ? 256'h6a : _GEN_58; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_60 = 8'h3c == io_in ? 256'h75 : _GEN_59; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_61 = 8'h3d == io_in ? 256'h37 : _GEN_60; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_62 = 8'h3e == io_in ? 256'h38 : _GEN_61; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_63 = 8'h3f == io_in ? 256'h0 : _GEN_62; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_64 = 8'h40 == io_in ? 256'h0 : _GEN_63; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_65 = 8'h41 == io_in ? 256'h0 : _GEN_64; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_66 = 8'h42 == io_in ? 256'h6b : _GEN_65; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_67 = 8'h43 == io_in ? 256'h69 : _GEN_66; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_68 = 8'h44 == io_in ? 256'h6f : _GEN_67; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_69 = 8'h45 == io_in ? 256'h30 : _GEN_68; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_70 = 8'h46 == io_in ? 256'h39 : _GEN_69; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_71 = 8'h47 == io_in ? 256'h0 : _GEN_70; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_72 = 8'h48 == io_in ? 256'h0 : _GEN_71; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_73 = 8'h49 == io_in ? 256'h0 : _GEN_72; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_74 = 8'h4a == io_in ? 256'h0 : _GEN_73; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_75 = 8'h4b == io_in ? 256'h6c : _GEN_74; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_76 = 8'h4c == io_in ? 256'h0 : _GEN_75; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_77 = 8'h4d == io_in ? 256'h70 : _GEN_76; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_78 = 8'h4e == io_in ? 256'h0 : _GEN_77; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_79 = 8'h4f == io_in ? 256'h0 : _GEN_78; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_80 = 8'h50 == io_in ? 256'h0 : _GEN_79; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_81 = 8'h51 == io_in ? 256'h0 : _GEN_80; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_82 = 8'h52 == io_in ? 256'h0 : _GEN_81; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_83 = 8'h53 == io_in ? 256'h0 : _GEN_82; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_84 = 8'h54 == io_in ? 256'h0 : _GEN_83; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_85 = 8'h55 == io_in ? 256'h0 : _GEN_84; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_86 = 8'h56 == io_in ? 256'h0 : _GEN_85; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_87 = 8'h57 == io_in ? 256'h0 : _GEN_86; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_88 = 8'h58 == io_in ? 256'h0 : _GEN_87; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_89 = 8'h59 == io_in ? 256'h0 : _GEN_88; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_90 = 8'h5a == io_in ? 256'h0 : _GEN_89; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_91 = 8'h5b == io_in ? 256'h0 : _GEN_90; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_92 = 8'h5c == io_in ? 256'h0 : _GEN_91; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_93 = 8'h5d == io_in ? 256'h0 : _GEN_92; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_94 = 8'h5e == io_in ? 256'h0 : _GEN_93; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_95 = 8'h5f == io_in ? 256'h0 : _GEN_94; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_96 = 8'h60 == io_in ? 256'h0 : _GEN_95; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_97 = 8'h61 == io_in ? 256'h0 : _GEN_96; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_98 = 8'h62 == io_in ? 256'h0 : _GEN_97; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_99 = 8'h63 == io_in ? 256'h0 : _GEN_98; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_100 = 8'h64 == io_in ? 256'h0 : _GEN_99; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_101 = 8'h65 == io_in ? 256'h0 : _GEN_100; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_102 = 8'h66 == io_in ? 256'h0 : _GEN_101; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_103 = 8'h67 == io_in ? 256'h0 : _GEN_102; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_104 = 8'h68 == io_in ? 256'h0 : _GEN_103; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_105 = 8'h69 == io_in ? 256'h0 : _GEN_104; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_106 = 8'h6a == io_in ? 256'h0 : _GEN_105; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_107 = 8'h6b == io_in ? 256'h0 : _GEN_106; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_108 = 8'h6c == io_in ? 256'h0 : _GEN_107; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_109 = 8'h6d == io_in ? 256'h0 : _GEN_108; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_110 = 8'h6e == io_in ? 256'h0 : _GEN_109; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_111 = 8'h6f == io_in ? 256'h0 : _GEN_110; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_112 = 8'h70 == io_in ? 256'h0 : _GEN_111; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_113 = 8'h71 == io_in ? 256'h0 : _GEN_112; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_114 = 8'h72 == io_in ? 256'h0 : _GEN_113; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_115 = 8'h73 == io_in ? 256'h0 : _GEN_114; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_116 = 8'h74 == io_in ? 256'h0 : _GEN_115; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_117 = 8'h75 == io_in ? 256'h0 : _GEN_116; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_118 = 8'h76 == io_in ? 256'h0 : _GEN_117; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_119 = 8'h77 == io_in ? 256'h0 : _GEN_118; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_120 = 8'h78 == io_in ? 256'h0 : _GEN_119; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_121 = 8'h79 == io_in ? 256'h0 : _GEN_120; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_122 = 8'h7a == io_in ? 256'h0 : _GEN_121; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_123 = 8'h7b == io_in ? 256'h0 : _GEN_122; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_124 = 8'h7c == io_in ? 256'h0 : _GEN_123; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_125 = 8'h7d == io_in ? 256'h0 : _GEN_124; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_126 = 8'h7e == io_in ? 256'h0 : _GEN_125; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_127 = 8'h7f == io_in ? 256'h0 : _GEN_126; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_128 = 8'h80 == io_in ? 256'h0 : _GEN_127; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_129 = 8'h81 == io_in ? 256'h0 : _GEN_128; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_130 = 8'h82 == io_in ? 256'h0 : _GEN_129; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_131 = 8'h83 == io_in ? 256'h0 : _GEN_130; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_132 = 8'h84 == io_in ? 256'h0 : _GEN_131; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_133 = 8'h85 == io_in ? 256'h0 : _GEN_132; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_134 = 8'h86 == io_in ? 256'h0 : _GEN_133; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_135 = 8'h87 == io_in ? 256'h0 : _GEN_134; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_136 = 8'h88 == io_in ? 256'h0 : _GEN_135; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_137 = 8'h89 == io_in ? 256'h0 : _GEN_136; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_138 = 8'h8a == io_in ? 256'h0 : _GEN_137; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_139 = 8'h8b == io_in ? 256'h0 : _GEN_138; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_140 = 8'h8c == io_in ? 256'h0 : _GEN_139; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_141 = 8'h8d == io_in ? 256'h0 : _GEN_140; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_142 = 8'h8e == io_in ? 256'h0 : _GEN_141; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_143 = 8'h8f == io_in ? 256'h0 : _GEN_142; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_144 = 8'h90 == io_in ? 256'h0 : _GEN_143; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_145 = 8'h91 == io_in ? 256'h0 : _GEN_144; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_146 = 8'h92 == io_in ? 256'h0 : _GEN_145; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_147 = 8'h93 == io_in ? 256'h0 : _GEN_146; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_148 = 8'h94 == io_in ? 256'h0 : _GEN_147; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_149 = 8'h95 == io_in ? 256'h0 : _GEN_148; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_150 = 8'h96 == io_in ? 256'h0 : _GEN_149; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_151 = 8'h97 == io_in ? 256'h0 : _GEN_150; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_152 = 8'h98 == io_in ? 256'h0 : _GEN_151; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_153 = 8'h99 == io_in ? 256'h0 : _GEN_152; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_154 = 8'h9a == io_in ? 256'h0 : _GEN_153; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_155 = 8'h9b == io_in ? 256'h0 : _GEN_154; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_156 = 8'h9c == io_in ? 256'h0 : _GEN_155; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_157 = 8'h9d == io_in ? 256'h0 : _GEN_156; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_158 = 8'h9e == io_in ? 256'h0 : _GEN_157; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_159 = 8'h9f == io_in ? 256'h0 : _GEN_158; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_160 = 8'ha0 == io_in ? 256'h0 : _GEN_159; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_161 = 8'ha1 == io_in ? 256'h0 : _GEN_160; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_162 = 8'ha2 == io_in ? 256'h0 : _GEN_161; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_163 = 8'ha3 == io_in ? 256'h0 : _GEN_162; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_164 = 8'ha4 == io_in ? 256'h0 : _GEN_163; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_165 = 8'ha5 == io_in ? 256'h0 : _GEN_164; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_166 = 8'ha6 == io_in ? 256'h0 : _GEN_165; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_167 = 8'ha7 == io_in ? 256'h0 : _GEN_166; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_168 = 8'ha8 == io_in ? 256'h0 : _GEN_167; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_169 = 8'ha9 == io_in ? 256'h0 : _GEN_168; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_170 = 8'haa == io_in ? 256'h0 : _GEN_169; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_171 = 8'hab == io_in ? 256'h0 : _GEN_170; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_172 = 8'hac == io_in ? 256'h0 : _GEN_171; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_173 = 8'had == io_in ? 256'h0 : _GEN_172; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_174 = 8'hae == io_in ? 256'h0 : _GEN_173; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_175 = 8'haf == io_in ? 256'h0 : _GEN_174; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_176 = 8'hb0 == io_in ? 256'h0 : _GEN_175; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_177 = 8'hb1 == io_in ? 256'h0 : _GEN_176; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_178 = 8'hb2 == io_in ? 256'h0 : _GEN_177; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_179 = 8'hb3 == io_in ? 256'h0 : _GEN_178; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_180 = 8'hb4 == io_in ? 256'h0 : _GEN_179; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_181 = 8'hb5 == io_in ? 256'h0 : _GEN_180; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_182 = 8'hb6 == io_in ? 256'h0 : _GEN_181; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_183 = 8'hb7 == io_in ? 256'h0 : _GEN_182; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_184 = 8'hb8 == io_in ? 256'h0 : _GEN_183; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_185 = 8'hb9 == io_in ? 256'h0 : _GEN_184; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_186 = 8'hba == io_in ? 256'h0 : _GEN_185; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_187 = 8'hbb == io_in ? 256'h0 : _GEN_186; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_188 = 8'hbc == io_in ? 256'h0 : _GEN_187; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_189 = 8'hbd == io_in ? 256'h0 : _GEN_188; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_190 = 8'hbe == io_in ? 256'h0 : _GEN_189; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_191 = 8'hbf == io_in ? 256'h0 : _GEN_190; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_192 = 8'hc0 == io_in ? 256'h0 : _GEN_191; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_193 = 8'hc1 == io_in ? 256'h0 : _GEN_192; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_194 = 8'hc2 == io_in ? 256'h0 : _GEN_193; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_195 = 8'hc3 == io_in ? 256'h0 : _GEN_194; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_196 = 8'hc4 == io_in ? 256'h0 : _GEN_195; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_197 = 8'hc5 == io_in ? 256'h0 : _GEN_196; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_198 = 8'hc6 == io_in ? 256'h0 : _GEN_197; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_199 = 8'hc7 == io_in ? 256'h0 : _GEN_198; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_200 = 8'hc8 == io_in ? 256'h0 : _GEN_199; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_201 = 8'hc9 == io_in ? 256'h0 : _GEN_200; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_202 = 8'hca == io_in ? 256'h0 : _GEN_201; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_203 = 8'hcb == io_in ? 256'h0 : _GEN_202; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_204 = 8'hcc == io_in ? 256'h0 : _GEN_203; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_205 = 8'hcd == io_in ? 256'h0 : _GEN_204; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_206 = 8'hce == io_in ? 256'h0 : _GEN_205; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_207 = 8'hcf == io_in ? 256'h0 : _GEN_206; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_208 = 8'hd0 == io_in ? 256'h0 : _GEN_207; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_209 = 8'hd1 == io_in ? 256'h0 : _GEN_208; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_210 = 8'hd2 == io_in ? 256'h0 : _GEN_209; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_211 = 8'hd3 == io_in ? 256'h0 : _GEN_210; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_212 = 8'hd4 == io_in ? 256'h0 : _GEN_211; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_213 = 8'hd5 == io_in ? 256'h0 : _GEN_212; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_214 = 8'hd6 == io_in ? 256'h0 : _GEN_213; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_215 = 8'hd7 == io_in ? 256'h0 : _GEN_214; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_216 = 8'hd8 == io_in ? 256'h0 : _GEN_215; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_217 = 8'hd9 == io_in ? 256'h0 : _GEN_216; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_218 = 8'hda == io_in ? 256'h0 : _GEN_217; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_219 = 8'hdb == io_in ? 256'h0 : _GEN_218; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_220 = 8'hdc == io_in ? 256'h0 : _GEN_219; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_221 = 8'hdd == io_in ? 256'h0 : _GEN_220; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_222 = 8'hde == io_in ? 256'h0 : _GEN_221; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_223 = 8'hdf == io_in ? 256'h0 : _GEN_222; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_224 = 8'he0 == io_in ? 256'h0 : _GEN_223; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_225 = 8'he1 == io_in ? 256'h0 : _GEN_224; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_226 = 8'he2 == io_in ? 256'h0 : _GEN_225; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_227 = 8'he3 == io_in ? 256'h0 : _GEN_226; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_228 = 8'he4 == io_in ? 256'h0 : _GEN_227; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_229 = 8'he5 == io_in ? 256'h0 : _GEN_228; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_230 = 8'he6 == io_in ? 256'h0 : _GEN_229; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_231 = 8'he7 == io_in ? 256'h0 : _GEN_230; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_232 = 8'he8 == io_in ? 256'h0 : _GEN_231; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_233 = 8'he9 == io_in ? 256'h0 : _GEN_232; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_234 = 8'hea == io_in ? 256'h0 : _GEN_233; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_235 = 8'heb == io_in ? 256'h0 : _GEN_234; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_236 = 8'hec == io_in ? 256'h0 : _GEN_235; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_237 = 8'hed == io_in ? 256'h0 : _GEN_236; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_238 = 8'hee == io_in ? 256'h0 : _GEN_237; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_239 = 8'hef == io_in ? 256'h0 : _GEN_238; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_240 = 8'hf0 == io_in ? 256'h0 : _GEN_239; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_241 = 8'hf1 == io_in ? 256'h0 : _GEN_240; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_242 = 8'hf2 == io_in ? 256'h0 : _GEN_241; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_243 = 8'hf3 == io_in ? 256'h0 : _GEN_242; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_244 = 8'hf4 == io_in ? 256'h0 : _GEN_243; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_245 = 8'hf5 == io_in ? 256'h0 : _GEN_244; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_246 = 8'hf6 == io_in ? 256'h0 : _GEN_245; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_247 = 8'hf7 == io_in ? 256'h0 : _GEN_246; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_248 = 8'hf8 == io_in ? 256'h0 : _GEN_247; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_249 = 8'hf9 == io_in ? 256'h0 : _GEN_248; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_250 = 8'hfa == io_in ? 256'h0 : _GEN_249; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_251 = 8'hfb == io_in ? 256'h0 : _GEN_250; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_252 = 8'hfc == io_in ? 256'h0 : _GEN_251; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_253 = 8'hfd == io_in ? 256'h0 : _GEN_252; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_254 = 8'hfe == io_in ? 256'h0 : _GEN_253; // @[ps2.scala 219:11 ps2.scala 219:11]
  wire [255:0] _GEN_255 = 8'hff == io_in ? 256'h0 : _GEN_254; // @[ps2.scala 219:11 ps2.scala 219:11]
  assign io_out = _GEN_255[7:0]; // @[ps2.scala 219:11]
endmodule
module seg(
  input        io_en,
  input  [3:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _GEN_0 = io_in == 4'hf ? 8'h8e : 8'hff; // @[ps2.scala 263:33 ps2.scala 264:19 ps2.scala 231:11]
  wire [7:0] _GEN_1 = io_in == 4'he ? 8'h86 : _GEN_0; // @[ps2.scala 261:33 ps2.scala 262:19]
  wire [7:0] _GEN_2 = io_in == 4'hd ? 8'ha1 : _GEN_1; // @[ps2.scala 259:33 ps2.scala 260:19]
  wire [7:0] _GEN_3 = io_in == 4'hc ? 8'hc6 : _GEN_2; // @[ps2.scala 257:33 ps2.scala 258:19]
  wire [7:0] _GEN_4 = io_in == 4'hb ? 8'h83 : _GEN_3; // @[ps2.scala 255:33 ps2.scala 256:19]
  wire [7:0] _GEN_5 = io_in == 4'ha ? 8'h88 : _GEN_4; // @[ps2.scala 253:33 ps2.scala 254:19]
  wire [7:0] _GEN_6 = io_in == 4'h9 ? 8'h90 : _GEN_5; // @[ps2.scala 251:32 ps2.scala 252:19]
  wire [7:0] _GEN_7 = io_in == 4'h8 ? 8'h80 : _GEN_6; // @[ps2.scala 249:32 ps2.scala 250:19]
  wire [7:0] _GEN_8 = io_in == 4'h7 ? 8'hf8 : _GEN_7; // @[ps2.scala 247:32 ps2.scala 248:19]
  wire [7:0] _GEN_9 = io_in == 4'h6 ? 8'h82 : _GEN_8; // @[ps2.scala 245:32 ps2.scala 246:19]
  wire [7:0] _GEN_10 = io_in == 4'h5 ? 8'h92 : _GEN_9; // @[ps2.scala 243:32 ps2.scala 244:19]
  wire [7:0] _GEN_11 = io_in == 4'h4 ? 8'h99 : _GEN_10; // @[ps2.scala 241:32 ps2.scala 242:19]
  wire [7:0] _GEN_12 = io_in == 4'h3 ? 8'hb0 : _GEN_11; // @[ps2.scala 239:32 ps2.scala 240:19]
  wire [7:0] _GEN_13 = io_in == 4'h2 ? 8'ha4 : _GEN_12; // @[ps2.scala 237:32 ps2.scala 238:19]
  wire [7:0] _GEN_14 = io_in == 4'h1 ? 8'hf9 : _GEN_13; // @[ps2.scala 235:32 ps2.scala 236:19]
  wire [7:0] _GEN_15 = io_in == 4'h0 ? 8'hc0 : _GEN_14; // @[ps2.scala 233:26 ps2.scala 234:19]
  assign io_out = io_en ? _GEN_15 : 8'hff; // @[ps2.scala 232:22 ps2.scala 267:15]
endmodule
module ps2(
  input        clock,
  input        reset,
  input        io_ps2_clk,
  input        io_ps2_data,
  output [7:0] io_ascii,
  output [1:0] io_now,
  output [7:0] io_bcd8seg_0,
  output [7:0] io_bcd8seg_1,
  output [7:0] io_bcd8seg_2,
  output [7:0] io_bcd8seg_3,
  output [7:0] io_bcd8seg_4,
  output [7:0] io_bcd8seg_5,
  output [7:0] io_bcd8seg_6,
  output [7:0] io_bcd8seg_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ps2_clock; // @[ps2.scala 17:19]
  wire  ps2_io_ps2_clk; // @[ps2.scala 17:19]
  wire  ps2_io_ps2_data; // @[ps2.scala 17:19]
  wire  ps2_io_nextdata_n; // @[ps2.scala 17:19]
  wire [7:0] ps2_io_data; // @[ps2.scala 17:19]
  wire  ps2_io_ready; // @[ps2.scala 17:19]
  wire [7:0] mm_io_in; // @[ps2.scala 73:18]
  wire [7:0] mm_io_out; // @[ps2.scala 73:18]
  wire  m0_io_en; // @[ps2.scala 78:18]
  wire [3:0] m0_io_in; // @[ps2.scala 78:18]
  wire [7:0] m0_io_out; // @[ps2.scala 78:18]
  wire  m1_io_en; // @[ps2.scala 82:18]
  wire [3:0] m1_io_in; // @[ps2.scala 82:18]
  wire [7:0] m1_io_out; // @[ps2.scala 82:18]
  wire  m2_io_en; // @[ps2.scala 86:18]
  wire [3:0] m2_io_in; // @[ps2.scala 86:18]
  wire [7:0] m2_io_out; // @[ps2.scala 86:18]
  wire  m3_io_en; // @[ps2.scala 90:18]
  wire [3:0] m3_io_in; // @[ps2.scala 90:18]
  wire [7:0] m3_io_out; // @[ps2.scala 90:18]
  wire  m4_io_en; // @[ps2.scala 94:18]
  wire [3:0] m4_io_in; // @[ps2.scala 94:18]
  wire [7:0] m4_io_out; // @[ps2.scala 94:18]
  wire  m5_io_en; // @[ps2.scala 98:18]
  wire [3:0] m5_io_in; // @[ps2.scala 98:18]
  wire [7:0] m5_io_out; // @[ps2.scala 98:18]
  wire  m6_io_en; // @[ps2.scala 102:18]
  wire [3:0] m6_io_in; // @[ps2.scala 102:18]
  wire [7:0] m6_io_out; // @[ps2.scala 102:18]
  wire  m7_io_en; // @[ps2.scala 106:18]
  wire [3:0] m7_io_in; // @[ps2.scala 106:18]
  wire [7:0] m7_io_out; // @[ps2.scala 106:18]
  reg [7:0] data; // @[ps2.scala 13:17]
  reg  ready; // @[ps2.scala 14:18]
  reg  nextdata; // @[ps2.scala 16:21]
  reg [3:0] now; // @[ps2.scala 31:20]
  reg [3:0] next; // @[ps2.scala 32:21]
  wire  _T = now == 4'h1; // @[ps2.scala 35:13]
  wire [1:0] _GEN_0 = ready ? 2'h2 : 2'h1; // @[ps2.scala 36:26 ps2.scala 37:17 ps2.scala 39:17]
  wire  _T_2 = now == 4'h2; // @[ps2.scala 41:19]
  wire  _T_3 = now == 4'h4; // @[ps2.scala 43:19]
  wire  _T_4 = now == 4'h8; // @[ps2.scala 45:19]
  reg [23:0] ps2segdata; // @[ps2.scala 50:27]
  wire [15:0] ps2segdata_hi = ps2segdata[15:0]; // @[ps2.scala 56:35]
  wire [23:0] _ps2segdata_T = {ps2segdata_hi,data}; // @[Cat.scala 30:58]
  wire  _GEN_6 = _T_2 ? nextdata : 1'h1; // @[ps2.scala 55:25 ps2.scala 16:21 ps2.scala 58:17]
  wire  _GEN_7 = _T_3 | _T_4 ? 1'h0 : _GEN_6; // @[ps2.scala 53:35 ps2.scala 54:17]
  reg [6:0] num; // @[ps2.scala 60:20]
  reg  segen; // @[ps2.scala 61:22]
  reg [1:0] ss; // @[ps2.scala 62:19]
  wire  ss_hi = ss[0]; // @[ps2.scala 68:15]
  wire [1:0] _ss_T = {ss_hi,segen}; // @[Cat.scala 30:58]
  wire [6:0] _num_T_1 = num + 7'h1; // @[ps2.scala 70:17]
  reg [7:0] ascii; // @[ps2.scala 72:22]
  wire [6:0] _GEN_1 = num % 7'ha; // @[ps2.scala 104:19]
  wire [6:0] _m6_io_in_T = _GEN_1[6:0]; // @[ps2.scala 104:19]
  wire [6:0] _m7_io_in_T = num / 7'ha; // @[ps2.scala 108:19]
  ps2_keyboard ps2 ( // @[ps2.scala 17:19]
    .clock(ps2_clock),
    .io_ps2_clk(ps2_io_ps2_clk),
    .io_ps2_data(ps2_io_ps2_data),
    .io_nextdata_n(ps2_io_nextdata_n),
    .io_data(ps2_io_data),
    .io_ready(ps2_io_ready)
  );
  ps2ascii mm ( // @[ps2.scala 73:18]
    .io_in(mm_io_in),
    .io_out(mm_io_out)
  );
  seg m0 ( // @[ps2.scala 78:18]
    .io_en(m0_io_en),
    .io_in(m0_io_in),
    .io_out(m0_io_out)
  );
  seg m1 ( // @[ps2.scala 82:18]
    .io_en(m1_io_en),
    .io_in(m1_io_in),
    .io_out(m1_io_out)
  );
  seg m2 ( // @[ps2.scala 86:18]
    .io_en(m2_io_en),
    .io_in(m2_io_in),
    .io_out(m2_io_out)
  );
  seg m3 ( // @[ps2.scala 90:18]
    .io_en(m3_io_en),
    .io_in(m3_io_in),
    .io_out(m3_io_out)
  );
  seg m4 ( // @[ps2.scala 94:18]
    .io_en(m4_io_en),
    .io_in(m4_io_in),
    .io_out(m4_io_out)
  );
  seg m5 ( // @[ps2.scala 98:18]
    .io_en(m5_io_en),
    .io_in(m5_io_in),
    .io_out(m5_io_out)
  );
  seg m6 ( // @[ps2.scala 102:18]
    .io_en(m6_io_en),
    .io_in(m6_io_in),
    .io_out(m6_io_out)
  );
  seg m7 ( // @[ps2.scala 106:18]
    .io_en(m7_io_en),
    .io_in(m7_io_in),
    .io_out(m7_io_out)
  );
  assign io_ascii = ascii; // @[ps2.scala 76:13]
  assign io_now = now[1:0]; // @[ps2.scala 33:11]
  assign io_bcd8seg_0 = m0_io_out; // @[ps2.scala 81:18]
  assign io_bcd8seg_1 = m1_io_out; // @[ps2.scala 85:18]
  assign io_bcd8seg_2 = m2_io_out; // @[ps2.scala 89:18]
  assign io_bcd8seg_3 = m3_io_out; // @[ps2.scala 93:18]
  assign io_bcd8seg_4 = m0_io_out; // @[ps2.scala 97:18]
  assign io_bcd8seg_5 = m0_io_out; // @[ps2.scala 101:18]
  assign io_bcd8seg_6 = m6_io_out; // @[ps2.scala 105:18]
  assign io_bcd8seg_7 = m7_io_out; // @[ps2.scala 109:18]
  assign ps2_clock = clock;
  assign ps2_io_ps2_clk = io_ps2_clk; // @[ps2.scala 19:19]
  assign ps2_io_ps2_data = io_ps2_data; // @[ps2.scala 20:20]
  assign ps2_io_nextdata_n = nextdata; // @[ps2.scala 21:22]
  assign mm_io_in = ps2segdata[7:0]; // @[ps2.scala 74:25]
  assign m0_io_en = segen; // @[ps2.scala 79:13]
  assign m0_io_in = ps2segdata[3:0]; // @[ps2.scala 80:25]
  assign m1_io_en = segen; // @[ps2.scala 83:13]
  assign m1_io_in = ps2segdata[7:4]; // @[ps2.scala 84:25]
  assign m2_io_en = segen; // @[ps2.scala 87:13]
  assign m2_io_in = ascii[3:0]; // @[ps2.scala 88:20]
  assign m3_io_en = segen; // @[ps2.scala 91:13]
  assign m3_io_in = ascii[7:4]; // @[ps2.scala 92:20]
  assign m4_io_en = 1'h0; // @[ps2.scala 95:13]
  assign m4_io_in = ps2segdata[3:0]; // @[ps2.scala 96:25]
  assign m5_io_en = 1'h0; // @[ps2.scala 99:13]
  assign m5_io_in = ps2segdata[7:4]; // @[ps2.scala 100:25]
  assign m6_io_en = 1'h1; // @[ps2.scala 103:13]
  assign m6_io_in = _m6_io_in_T[3:0]; // @[ps2.scala 104:30]
  assign m7_io_en = 1'h1; // @[ps2.scala 107:13]
  assign m7_io_in = _m7_io_in_T[3:0]; // @[ps2.scala 108:30]
  always @(posedge clock) begin
    data <= ps2_io_data; // @[ps2.scala 22:9]
    ready <= ps2_io_ready; // @[ps2.scala 23:10]
    nextdata <= _T | _GEN_7; // @[ps2.scala 51:19 ps2.scala 52:17]
    if (reset) begin // @[ps2.scala 31:20]
      now <= 4'h1; // @[ps2.scala 31:20]
    end else begin
      now <= next; // @[ps2.scala 34:8]
    end
    if (reset) begin // @[ps2.scala 32:21]
      next <= 4'h1; // @[ps2.scala 32:21]
    end else if (now == 4'h1) begin // @[ps2.scala 35:19]
      next <= {{2'd0}, _GEN_0};
    end else if (now == 4'h2) begin // @[ps2.scala 41:25]
      next <= 4'h4; // @[ps2.scala 42:13]
    end else if (now == 4'h4) begin // @[ps2.scala 43:25]
      next <= 4'h8; // @[ps2.scala 44:13]
    end else begin
      next <= 4'h1;
    end
    if (reset) begin // @[ps2.scala 50:27]
      ps2segdata <= 24'h0; // @[ps2.scala 50:27]
    end else if (!(_T)) begin // @[ps2.scala 51:19]
      if (!(_T_3 | _T_4)) begin // @[ps2.scala 53:35]
        if (_T_2) begin // @[ps2.scala 55:25]
          ps2segdata <= _ps2segdata_T; // @[ps2.scala 56:19]
        end
      end
    end
    if (reset) begin // @[ps2.scala 60:20]
      num <= 7'h0; // @[ps2.scala 60:20]
    end else if (ss == 2'h2) begin // @[ps2.scala 69:23]
      num <= _num_T_1; // @[ps2.scala 70:12]
    end
    if (reset) begin // @[ps2.scala 61:22]
      segen <= 1'h0; // @[ps2.scala 61:22]
    end else if (ps2segdata[23:16] == 8'hf0 & ps2segdata[7:0] == ps2segdata[15:8]) begin // @[ps2.scala 63:78]
      segen <= 1'h0; // @[ps2.scala 64:14]
    end else begin
      segen <= 1'h1; // @[ps2.scala 66:14]
    end
    if (reset) begin // @[ps2.scala 62:19]
      ss <= 2'h0; // @[ps2.scala 62:19]
    end else begin
      ss <= _ss_T; // @[ps2.scala 68:7]
    end
    if (reset) begin // @[ps2.scala 72:22]
      ascii <= 8'h0; // @[ps2.scala 72:22]
    end else begin
      ascii <= mm_io_out; // @[ps2.scala 75:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  ready = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  nextdata = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  now = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  next = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  ps2segdata = _RAND_5[23:0];
  _RAND_6 = {1{`RANDOM}};
  num = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  segen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ss = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ascii = _RAND_9[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vga_ctrl(
  input         clock,
  input         reset,
  input  [23:0] io_vga_data,
  output [9:0]  io_h_addr,
  output [9:0]  io_v_addr,
  output        io_hsync,
  output        io_vsync,
  output        io_valid,
  output [7:0]  io_vga_r,
  output [7:0]  io_vga_g,
  output [7:0]  io_vga_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] x_cnt; // @[vga.scala 98:22]
  reg [9:0] y_cnt; // @[vga.scala 99:22]
  wire  _T = x_cnt == 10'h320; // @[vga.scala 101:15]
  wire [9:0] _x_cnt_T_1 = x_cnt + 10'h1; // @[vga.scala 104:21]
  wire [9:0] _y_cnt_T_1 = y_cnt + 10'h1; // @[vga.scala 109:21]
  wire  h_valid = x_cnt > 10'h90 & x_cnt <= 10'h310; // @[vga.scala 113:39]
  wire  v_valid = y_cnt > 10'h23 & y_cnt <= 10'h203; // @[vga.scala 114:39]
  wire [9:0] _io_h_addr_T_1 = x_cnt - 10'h91; // @[vga.scala 116:33]
  wire [9:0] _io_v_addr_T_1 = y_cnt - 10'h24; // @[vga.scala 117:33]
  assign io_h_addr = h_valid ? _io_h_addr_T_1 : 10'h0; // @[vga.scala 116:19]
  assign io_v_addr = v_valid ? _io_v_addr_T_1 : 10'h0; // @[vga.scala 117:19]
  assign io_hsync = x_cnt > 10'h60; // @[vga.scala 111:21]
  assign io_vsync = y_cnt > 10'h2; // @[vga.scala 112:21]
  assign io_valid = h_valid & v_valid; // @[vga.scala 115:23]
  assign io_vga_r = io_vga_data[23:16]; // @[vga.scala 118:26]
  assign io_vga_g = io_vga_data[15:8]; // @[vga.scala 119:26]
  assign io_vga_b = io_vga_data[7:0]; // @[vga.scala 120:26]
  always @(posedge clock) begin
    if (reset) begin // @[vga.scala 98:22]
      x_cnt <= 10'h1; // @[vga.scala 98:22]
    end else if (x_cnt == 10'h320) begin // @[vga.scala 101:26]
      x_cnt <= 10'h1; // @[vga.scala 102:14]
    end else begin
      x_cnt <= _x_cnt_T_1; // @[vga.scala 104:14]
    end
    if (reset) begin // @[vga.scala 99:22]
      y_cnt <= 10'h1; // @[vga.scala 99:22]
    end else if (y_cnt == 10'h20d & _T) begin // @[vga.scala 106:47]
      y_cnt <= 10'h1; // @[vga.scala 107:14]
    end else if (_T) begin // @[vga.scala 108:32]
      y_cnt <= _y_cnt_T_1; // @[vga.scala 109:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_cnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  y_cnt = _RAND_1[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vmem(
  input         clock,
  input         reset,
  input  [1:0]  io_now,
  input  [7:0]  io_ascii,
  input  [9:0]  io_h_addr,
  input  [8:0]  io_v_addr,
  output [23:0] io_vga_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [287:0] _RAND_306;
  reg [287:0] _RAND_307;
  reg [287:0] _RAND_308;
  reg [287:0] _RAND_309;
  reg [287:0] _RAND_310;
  reg [287:0] _RAND_311;
  reg [287:0] _RAND_312;
  reg [287:0] _RAND_313;
  reg [287:0] _RAND_314;
  reg [287:0] _RAND_315;
  reg [287:0] _RAND_316;
  reg [287:0] _RAND_317;
  reg [287:0] _RAND_318;
  reg [287:0] _RAND_319;
  reg [287:0] _RAND_320;
  reg [287:0] _RAND_321;
  reg [287:0] _RAND_322;
  reg [287:0] _RAND_323;
  reg [287:0] _RAND_324;
  reg [287:0] _RAND_325;
  reg [287:0] _RAND_326;
  reg [287:0] _RAND_327;
  reg [287:0] _RAND_328;
  reg [287:0] _RAND_329;
  reg [287:0] _RAND_330;
  reg [287:0] _RAND_331;
  reg [287:0] _RAND_332;
  reg [287:0] _RAND_333;
  reg [287:0] _RAND_334;
  reg [287:0] _RAND_335;
  reg [287:0] _RAND_336;
  reg [287:0] _RAND_337;
  reg [287:0] _RAND_338;
  reg [287:0] _RAND_339;
  reg [287:0] _RAND_340;
  reg [287:0] _RAND_341;
  reg [287:0] _RAND_342;
  reg [287:0] _RAND_343;
  reg [287:0] _RAND_344;
  reg [287:0] _RAND_345;
  reg [287:0] _RAND_346;
  reg [287:0] _RAND_347;
  reg [287:0] _RAND_348;
  reg [287:0] _RAND_349;
  reg [287:0] _RAND_350;
  reg [287:0] _RAND_351;
  reg [287:0] _RAND_352;
  reg [287:0] _RAND_353;
  reg [287:0] _RAND_354;
  reg [287:0] _RAND_355;
  reg [287:0] _RAND_356;
  reg [287:0] _RAND_357;
  reg [287:0] _RAND_358;
  reg [287:0] _RAND_359;
  reg [287:0] _RAND_360;
  reg [287:0] _RAND_361;
  reg [287:0] _RAND_362;
  reg [287:0] _RAND_363;
  reg [287:0] _RAND_364;
  reg [287:0] _RAND_365;
  reg [287:0] _RAND_366;
  reg [287:0] _RAND_367;
  reg [287:0] _RAND_368;
  reg [287:0] _RAND_369;
  reg [287:0] _RAND_370;
  reg [287:0] _RAND_371;
  reg [287:0] _RAND_372;
  reg [287:0] _RAND_373;
  reg [287:0] _RAND_374;
  reg [287:0] _RAND_375;
  reg [287:0] _RAND_376;
  reg [287:0] _RAND_377;
  reg [287:0] _RAND_378;
  reg [287:0] _RAND_379;
  reg [287:0] _RAND_380;
  reg [287:0] _RAND_381;
  reg [287:0] _RAND_382;
  reg [287:0] _RAND_383;
  reg [287:0] _RAND_384;
  reg [287:0] _RAND_385;
  reg [287:0] _RAND_386;
  reg [287:0] _RAND_387;
  reg [287:0] _RAND_388;
  reg [287:0] _RAND_389;
  reg [287:0] _RAND_390;
  reg [287:0] _RAND_391;
  reg [287:0] _RAND_392;
  reg [287:0] _RAND_393;
  reg [287:0] _RAND_394;
  reg [287:0] _RAND_395;
  reg [287:0] _RAND_396;
  reg [287:0] _RAND_397;
  reg [287:0] _RAND_398;
  reg [287:0] _RAND_399;
  reg [287:0] _RAND_400;
  reg [287:0] _RAND_401;
  reg [287:0] _RAND_402;
  reg [287:0] _RAND_403;
  reg [287:0] _RAND_404;
  reg [287:0] _RAND_405;
  reg [287:0] _RAND_406;
  reg [287:0] _RAND_407;
  reg [287:0] _RAND_408;
  reg [287:0] _RAND_409;
  reg [287:0] _RAND_410;
  reg [287:0] _RAND_411;
  reg [287:0] _RAND_412;
  reg [287:0] _RAND_413;
  reg [287:0] _RAND_414;
  reg [287:0] _RAND_415;
  reg [287:0] _RAND_416;
  reg [287:0] _RAND_417;
  reg [287:0] _RAND_418;
  reg [287:0] _RAND_419;
  reg [287:0] _RAND_420;
  reg [287:0] _RAND_421;
  reg [287:0] _RAND_422;
  reg [287:0] _RAND_423;
  reg [287:0] _RAND_424;
  reg [287:0] _RAND_425;
  reg [287:0] _RAND_426;
  reg [287:0] _RAND_427;
  reg [287:0] _RAND_428;
  reg [287:0] _RAND_429;
  reg [287:0] _RAND_430;
  reg [287:0] _RAND_431;
  reg [287:0] _RAND_432;
  reg [287:0] _RAND_433;
  reg [287:0] _RAND_434;
  reg [287:0] _RAND_435;
  reg [287:0] _RAND_436;
  reg [287:0] _RAND_437;
  reg [287:0] _RAND_438;
  reg [287:0] _RAND_439;
  reg [287:0] _RAND_440;
  reg [287:0] _RAND_441;
  reg [287:0] _RAND_442;
  reg [287:0] _RAND_443;
  reg [287:0] _RAND_444;
  reg [287:0] _RAND_445;
  reg [287:0] _RAND_446;
  reg [287:0] _RAND_447;
  reg [287:0] _RAND_448;
  reg [287:0] _RAND_449;
  reg [287:0] _RAND_450;
  reg [287:0] _RAND_451;
  reg [287:0] _RAND_452;
  reg [287:0] _RAND_453;
  reg [287:0] _RAND_454;
  reg [287:0] _RAND_455;
  reg [287:0] _RAND_456;
  reg [287:0] _RAND_457;
  reg [287:0] _RAND_458;
  reg [287:0] _RAND_459;
  reg [287:0] _RAND_460;
  reg [287:0] _RAND_461;
  reg [287:0] _RAND_462;
  reg [287:0] _RAND_463;
  reg [287:0] _RAND_464;
  reg [287:0] _RAND_465;
  reg [287:0] _RAND_466;
  reg [287:0] _RAND_467;
  reg [287:0] _RAND_468;
  reg [287:0] _RAND_469;
  reg [287:0] _RAND_470;
  reg [287:0] _RAND_471;
  reg [287:0] _RAND_472;
  reg [287:0] _RAND_473;
  reg [287:0] _RAND_474;
  reg [287:0] _RAND_475;
  reg [287:0] _RAND_476;
  reg [287:0] _RAND_477;
  reg [287:0] _RAND_478;
  reg [287:0] _RAND_479;
  reg [287:0] _RAND_480;
  reg [287:0] _RAND_481;
  reg [287:0] _RAND_482;
  reg [287:0] _RAND_483;
  reg [287:0] _RAND_484;
  reg [287:0] _RAND_485;
  reg [287:0] _RAND_486;
  reg [287:0] _RAND_487;
  reg [287:0] _RAND_488;
  reg [287:0] _RAND_489;
  reg [287:0] _RAND_490;
  reg [287:0] _RAND_491;
  reg [287:0] _RAND_492;
  reg [287:0] _RAND_493;
  reg [287:0] _RAND_494;
  reg [287:0] _RAND_495;
  reg [287:0] _RAND_496;
  reg [287:0] _RAND_497;
  reg [287:0] _RAND_498;
  reg [287:0] _RAND_499;
  reg [287:0] _RAND_500;
  reg [287:0] _RAND_501;
  reg [287:0] _RAND_502;
  reg [287:0] _RAND_503;
  reg [287:0] _RAND_504;
  reg [287:0] _RAND_505;
  reg [287:0] _RAND_506;
  reg [287:0] _RAND_507;
  reg [287:0] _RAND_508;
  reg [287:0] _RAND_509;
  reg [287:0] _RAND_510;
  reg [287:0] _RAND_511;
  reg [287:0] _RAND_512;
  reg [287:0] _RAND_513;
  reg [287:0] _RAND_514;
  reg [287:0] _RAND_515;
  reg [287:0] _RAND_516;
  reg [287:0] _RAND_517;
  reg [287:0] _RAND_518;
  reg [287:0] _RAND_519;
  reg [287:0] _RAND_520;
  reg [287:0] _RAND_521;
  reg [287:0] _RAND_522;
  reg [287:0] _RAND_523;
  reg [287:0] _RAND_524;
  reg [287:0] _RAND_525;
  reg [287:0] _RAND_526;
  reg [287:0] _RAND_527;
  reg [287:0] _RAND_528;
  reg [287:0] _RAND_529;
  reg [287:0] _RAND_530;
  reg [287:0] _RAND_531;
  reg [287:0] _RAND_532;
  reg [287:0] _RAND_533;
  reg [287:0] _RAND_534;
  reg [287:0] _RAND_535;
  reg [287:0] _RAND_536;
  reg [287:0] _RAND_537;
  reg [287:0] _RAND_538;
  reg [287:0] _RAND_539;
  reg [287:0] _RAND_540;
  reg [287:0] _RAND_541;
  reg [287:0] _RAND_542;
  reg [287:0] _RAND_543;
  reg [287:0] _RAND_544;
  reg [287:0] _RAND_545;
  reg [287:0] _RAND_546;
  reg [287:0] _RAND_547;
  reg [287:0] _RAND_548;
  reg [287:0] _RAND_549;
  reg [287:0] _RAND_550;
  reg [287:0] _RAND_551;
  reg [287:0] _RAND_552;
  reg [287:0] _RAND_553;
  reg [287:0] _RAND_554;
  reg [287:0] _RAND_555;
  reg [287:0] _RAND_556;
  reg [287:0] _RAND_557;
  reg [287:0] _RAND_558;
  reg [287:0] _RAND_559;
  reg [287:0] _RAND_560;
  reg [287:0] _RAND_561;
  reg [287:0] _RAND_562;
  reg [287:0] _RAND_563;
  reg [287:0] _RAND_564;
  reg [287:0] _RAND_565;
  reg [287:0] _RAND_566;
  reg [287:0] _RAND_567;
  reg [287:0] _RAND_568;
  reg [287:0] _RAND_569;
  reg [287:0] _RAND_570;
  reg [287:0] _RAND_571;
  reg [287:0] _RAND_572;
  reg [287:0] _RAND_573;
  reg [287:0] _RAND_574;
  reg [287:0] _RAND_575;
  reg [287:0] _RAND_576;
  reg [287:0] _RAND_577;
  reg [287:0] _RAND_578;
  reg [287:0] _RAND_579;
  reg [287:0] _RAND_580;
  reg [287:0] _RAND_581;
  reg [287:0] _RAND_582;
  reg [287:0] _RAND_583;
  reg [287:0] _RAND_584;
  reg [287:0] _RAND_585;
  reg [287:0] _RAND_586;
  reg [287:0] _RAND_587;
  reg [287:0] _RAND_588;
  reg [287:0] _RAND_589;
  reg [287:0] _RAND_590;
  reg [287:0] _RAND_591;
  reg [287:0] _RAND_592;
  reg [287:0] _RAND_593;
  reg [287:0] _RAND_594;
  reg [287:0] _RAND_595;
  reg [287:0] _RAND_596;
  reg [287:0] _RAND_597;
  reg [287:0] _RAND_598;
  reg [287:0] _RAND_599;
  reg [287:0] _RAND_600;
  reg [287:0] _RAND_601;
  reg [287:0] _RAND_602;
  reg [287:0] _RAND_603;
  reg [287:0] _RAND_604;
  reg [287:0] _RAND_605;
  reg [287:0] _RAND_606;
  reg [287:0] _RAND_607;
  reg [287:0] _RAND_608;
  reg [287:0] _RAND_609;
  reg [287:0] _RAND_610;
  reg [287:0] _RAND_611;
  reg [287:0] _RAND_612;
  reg [287:0] _RAND_613;
  reg [287:0] _RAND_614;
  reg [287:0] _RAND_615;
  reg [287:0] _RAND_616;
  reg [287:0] _RAND_617;
  reg [287:0] _RAND_618;
  reg [287:0] _RAND_619;
  reg [287:0] _RAND_620;
  reg [287:0] _RAND_621;
  reg [287:0] _RAND_622;
  reg [287:0] _RAND_623;
  reg [287:0] _RAND_624;
  reg [287:0] _RAND_625;
  reg [287:0] _RAND_626;
  reg [287:0] _RAND_627;
  reg [287:0] _RAND_628;
  reg [287:0] _RAND_629;
  reg [287:0] _RAND_630;
  reg [287:0] _RAND_631;
  reg [287:0] _RAND_632;
  reg [287:0] _RAND_633;
  reg [287:0] _RAND_634;
  reg [287:0] _RAND_635;
  reg [287:0] _RAND_636;
  reg [287:0] _RAND_637;
  reg [287:0] _RAND_638;
  reg [287:0] _RAND_639;
  reg [287:0] _RAND_640;
  reg [287:0] _RAND_641;
  reg [287:0] _RAND_642;
  reg [287:0] _RAND_643;
  reg [287:0] _RAND_644;
  reg [287:0] _RAND_645;
  reg [287:0] _RAND_646;
  reg [287:0] _RAND_647;
  reg [287:0] _RAND_648;
  reg [287:0] _RAND_649;
  reg [287:0] _RAND_650;
  reg [287:0] _RAND_651;
  reg [287:0] _RAND_652;
  reg [287:0] _RAND_653;
  reg [287:0] _RAND_654;
  reg [287:0] _RAND_655;
  reg [287:0] _RAND_656;
  reg [287:0] _RAND_657;
  reg [287:0] _RAND_658;
  reg [287:0] _RAND_659;
  reg [287:0] _RAND_660;
  reg [287:0] _RAND_661;
  reg [287:0] _RAND_662;
  reg [287:0] _RAND_663;
  reg [287:0] _RAND_664;
  reg [287:0] _RAND_665;
  reg [287:0] _RAND_666;
  reg [287:0] _RAND_667;
  reg [287:0] _RAND_668;
  reg [287:0] _RAND_669;
  reg [287:0] _RAND_670;
  reg [287:0] _RAND_671;
  reg [287:0] _RAND_672;
  reg [287:0] _RAND_673;
  reg [287:0] _RAND_674;
  reg [287:0] _RAND_675;
  reg [287:0] _RAND_676;
  reg [287:0] _RAND_677;
  reg [287:0] _RAND_678;
  reg [287:0] _RAND_679;
  reg [287:0] _RAND_680;
  reg [287:0] _RAND_681;
  reg [287:0] _RAND_682;
  reg [287:0] _RAND_683;
  reg [287:0] _RAND_684;
  reg [287:0] _RAND_685;
  reg [287:0] _RAND_686;
  reg [287:0] _RAND_687;
  reg [287:0] _RAND_688;
  reg [287:0] _RAND_689;
  reg [287:0] _RAND_690;
  reg [287:0] _RAND_691;
  reg [287:0] _RAND_692;
  reg [287:0] _RAND_693;
  reg [287:0] _RAND_694;
  reg [287:0] _RAND_695;
  reg [287:0] _RAND_696;
  reg [287:0] _RAND_697;
  reg [287:0] _RAND_698;
  reg [287:0] _RAND_699;
  reg [287:0] _RAND_700;
  reg [287:0] _RAND_701;
  reg [287:0] _RAND_702;
  reg [287:0] _RAND_703;
  reg [287:0] _RAND_704;
  reg [287:0] _RAND_705;
  reg [287:0] _RAND_706;
  reg [287:0] _RAND_707;
  reg [287:0] _RAND_708;
  reg [287:0] _RAND_709;
  reg [287:0] _RAND_710;
  reg [287:0] _RAND_711;
  reg [287:0] _RAND_712;
  reg [287:0] _RAND_713;
  reg [287:0] _RAND_714;
  reg [287:0] _RAND_715;
  reg [287:0] _RAND_716;
  reg [287:0] _RAND_717;
  reg [287:0] _RAND_718;
  reg [287:0] _RAND_719;
  reg [287:0] _RAND_720;
  reg [287:0] _RAND_721;
  reg [287:0] _RAND_722;
  reg [287:0] _RAND_723;
  reg [287:0] _RAND_724;
  reg [287:0] _RAND_725;
  reg [287:0] _RAND_726;
  reg [287:0] _RAND_727;
  reg [287:0] _RAND_728;
  reg [287:0] _RAND_729;
  reg [287:0] _RAND_730;
  reg [287:0] _RAND_731;
  reg [287:0] _RAND_732;
  reg [287:0] _RAND_733;
  reg [287:0] _RAND_734;
  reg [287:0] _RAND_735;
  reg [287:0] _RAND_736;
  reg [287:0] _RAND_737;
  reg [287:0] _RAND_738;
  reg [287:0] _RAND_739;
  reg [287:0] _RAND_740;
  reg [287:0] _RAND_741;
  reg [287:0] _RAND_742;
  reg [287:0] _RAND_743;
  reg [287:0] _RAND_744;
  reg [287:0] _RAND_745;
  reg [287:0] _RAND_746;
  reg [287:0] _RAND_747;
  reg [287:0] _RAND_748;
  reg [287:0] _RAND_749;
  reg [287:0] _RAND_750;
  reg [287:0] _RAND_751;
  reg [287:0] _RAND_752;
  reg [287:0] _RAND_753;
  reg [287:0] _RAND_754;
  reg [287:0] _RAND_755;
  reg [287:0] _RAND_756;
  reg [287:0] _RAND_757;
  reg [287:0] _RAND_758;
  reg [287:0] _RAND_759;
  reg [287:0] _RAND_760;
  reg [287:0] _RAND_761;
  reg [287:0] _RAND_762;
  reg [287:0] _RAND_763;
  reg [287:0] _RAND_764;
  reg [287:0] _RAND_765;
  reg [287:0] _RAND_766;
  reg [287:0] _RAND_767;
  reg [287:0] _RAND_768;
  reg [287:0] _RAND_769;
  reg [287:0] _RAND_770;
  reg [287:0] _RAND_771;
  reg [287:0] _RAND_772;
  reg [287:0] _RAND_773;
  reg [287:0] _RAND_774;
  reg [287:0] _RAND_775;
  reg [287:0] _RAND_776;
  reg [287:0] _RAND_777;
  reg [287:0] _RAND_778;
  reg [287:0] _RAND_779;
  reg [287:0] _RAND_780;
  reg [287:0] _RAND_781;
  reg [287:0] _RAND_782;
  reg [287:0] _RAND_783;
  reg [287:0] _RAND_784;
  reg [287:0] _RAND_785;
  reg [287:0] _RAND_786;
  reg [287:0] _RAND_787;
  reg [287:0] _RAND_788;
  reg [287:0] _RAND_789;
  reg [287:0] _RAND_790;
  reg [287:0] _RAND_791;
  reg [287:0] _RAND_792;
  reg [287:0] _RAND_793;
  reg [287:0] _RAND_794;
  reg [287:0] _RAND_795;
  reg [287:0] _RAND_796;
  reg [287:0] _RAND_797;
  reg [287:0] _RAND_798;
  reg [287:0] _RAND_799;
  reg [287:0] _RAND_800;
  reg [287:0] _RAND_801;
  reg [287:0] _RAND_802;
  reg [287:0] _RAND_803;
  reg [287:0] _RAND_804;
  reg [287:0] _RAND_805;
  reg [287:0] _RAND_806;
  reg [287:0] _RAND_807;
  reg [287:0] _RAND_808;
  reg [287:0] _RAND_809;
  reg [287:0] _RAND_810;
  reg [287:0] _RAND_811;
  reg [287:0] _RAND_812;
  reg [287:0] _RAND_813;
  reg [287:0] _RAND_814;
  reg [287:0] _RAND_815;
  reg [287:0] _RAND_816;
  reg [287:0] _RAND_817;
  reg [287:0] _RAND_818;
  reg [287:0] _RAND_819;
  reg [287:0] _RAND_820;
  reg [287:0] _RAND_821;
  reg [287:0] _RAND_822;
  reg [287:0] _RAND_823;
  reg [287:0] _RAND_824;
  reg [287:0] _RAND_825;
  reg [287:0] _RAND_826;
  reg [287:0] _RAND_827;
  reg [287:0] _RAND_828;
  reg [287:0] _RAND_829;
  reg [287:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
`endif // RANDOMIZE_REG_INIT
  reg [11:0] vga_mem [0:4095]; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_1_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_1_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_2_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_2_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_3_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_3_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_4_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_4_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_5_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_5_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_6_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_6_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_7_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_7_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_8_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_8_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_9_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_9_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_10_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_10_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_11_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_11_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_12_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_12_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_13_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_13_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_14_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_14_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_15_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_15_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_16_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_16_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_17_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_17_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_18_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_18_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_19_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_19_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_20_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_20_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_21_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_21_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_22_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_22_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_23_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_23_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_24_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_24_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_25_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_25_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_26_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_26_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_27_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_27_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_28_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_28_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_29_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_29_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_30_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_30_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_31_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_31_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_32_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_32_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_33_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_33_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_34_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_34_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_35_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_35_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_36_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_36_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_37_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_37_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_38_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_38_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_39_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_39_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_40_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_40_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_41_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_41_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_42_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_42_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_43_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_43_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_44_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_44_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_45_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_45_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_46_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_46_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_47_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_47_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_48_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_48_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_49_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_49_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_50_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_50_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_51_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_51_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_52_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_52_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_53_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_53_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_54_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_54_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_55_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_55_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_56_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_56_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_57_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_57_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_58_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_58_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_59_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_59_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_60_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_60_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_61_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_61_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_62_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_62_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_63_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_63_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_64_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_64_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_65_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_65_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_66_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_66_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_67_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_67_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_68_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_68_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_69_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_69_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_70_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_70_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_71_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_71_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_72_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_72_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_73_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_73_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_74_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_74_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_75_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_75_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_76_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_76_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_77_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_77_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_78_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_78_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_79_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_79_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_80_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_80_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_81_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_81_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_82_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_82_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_83_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_83_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_84_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_84_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_85_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_85_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_86_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_86_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_87_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_87_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_88_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_88_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_89_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_89_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_90_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_90_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_91_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_91_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_92_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_92_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_93_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_93_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_94_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_94_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_95_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_95_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_96_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_96_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_97_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_97_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_98_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_98_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_99_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_99_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_100_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_100_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_101_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_101_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_102_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_102_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_103_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_103_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_104_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_104_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_105_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_105_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_106_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_106_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_107_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_107_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_108_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_108_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_109_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_109_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_110_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_110_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_111_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_111_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_112_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_112_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_113_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_113_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_114_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_114_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_115_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_115_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_116_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_116_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_117_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_117_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_118_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_118_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_119_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_119_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_120_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_120_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_121_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_121_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_122_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_122_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_123_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_123_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_124_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_124_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_125_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_125_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_126_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_126_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_127_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_127_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_128_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_128_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_129_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_129_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_130_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_130_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_131_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_131_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_132_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_132_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_133_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_133_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_134_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_134_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_135_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_135_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_136_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_136_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_137_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_137_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_138_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_138_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_139_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_139_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_140_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_140_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_141_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_141_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_142_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_142_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_143_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_143_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_144_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_144_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_145_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_145_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_146_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_146_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_147_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_147_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_148_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_148_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_149_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_149_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_150_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_150_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_151_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_151_addr; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_152_data; // @[vga.scala 50:30]
  wire [11:0] vga_mem_ram_MPORT_152_addr; // @[vga.scala 50:30]
  reg  vga_mem_ram_MPORT_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_addr_pipe_0;
  reg  vga_mem_ram_MPORT_1_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_1_addr_pipe_0;
  reg  vga_mem_ram_MPORT_2_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_2_addr_pipe_0;
  reg  vga_mem_ram_MPORT_3_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_3_addr_pipe_0;
  reg  vga_mem_ram_MPORT_4_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_4_addr_pipe_0;
  reg  vga_mem_ram_MPORT_5_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_5_addr_pipe_0;
  reg  vga_mem_ram_MPORT_6_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_6_addr_pipe_0;
  reg  vga_mem_ram_MPORT_7_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_7_addr_pipe_0;
  reg  vga_mem_ram_MPORT_8_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_8_addr_pipe_0;
  reg  vga_mem_ram_MPORT_9_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_9_addr_pipe_0;
  reg  vga_mem_ram_MPORT_10_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_10_addr_pipe_0;
  reg  vga_mem_ram_MPORT_11_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_11_addr_pipe_0;
  reg  vga_mem_ram_MPORT_12_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_12_addr_pipe_0;
  reg  vga_mem_ram_MPORT_13_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_13_addr_pipe_0;
  reg  vga_mem_ram_MPORT_14_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_14_addr_pipe_0;
  reg  vga_mem_ram_MPORT_15_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_15_addr_pipe_0;
  reg  vga_mem_ram_MPORT_16_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_16_addr_pipe_0;
  reg  vga_mem_ram_MPORT_17_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_17_addr_pipe_0;
  reg  vga_mem_ram_MPORT_18_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_18_addr_pipe_0;
  reg  vga_mem_ram_MPORT_19_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_19_addr_pipe_0;
  reg  vga_mem_ram_MPORT_20_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_20_addr_pipe_0;
  reg  vga_mem_ram_MPORT_21_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_21_addr_pipe_0;
  reg  vga_mem_ram_MPORT_22_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_22_addr_pipe_0;
  reg  vga_mem_ram_MPORT_23_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_23_addr_pipe_0;
  reg  vga_mem_ram_MPORT_24_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_24_addr_pipe_0;
  reg  vga_mem_ram_MPORT_25_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_25_addr_pipe_0;
  reg  vga_mem_ram_MPORT_26_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_26_addr_pipe_0;
  reg  vga_mem_ram_MPORT_27_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_27_addr_pipe_0;
  reg  vga_mem_ram_MPORT_28_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_28_addr_pipe_0;
  reg  vga_mem_ram_MPORT_29_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_29_addr_pipe_0;
  reg  vga_mem_ram_MPORT_30_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_30_addr_pipe_0;
  reg  vga_mem_ram_MPORT_31_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_31_addr_pipe_0;
  reg  vga_mem_ram_MPORT_32_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_32_addr_pipe_0;
  reg  vga_mem_ram_MPORT_33_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_33_addr_pipe_0;
  reg  vga_mem_ram_MPORT_34_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_34_addr_pipe_0;
  reg  vga_mem_ram_MPORT_35_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_35_addr_pipe_0;
  reg  vga_mem_ram_MPORT_36_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_36_addr_pipe_0;
  reg  vga_mem_ram_MPORT_37_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_37_addr_pipe_0;
  reg  vga_mem_ram_MPORT_38_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_38_addr_pipe_0;
  reg  vga_mem_ram_MPORT_39_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_39_addr_pipe_0;
  reg  vga_mem_ram_MPORT_40_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_40_addr_pipe_0;
  reg  vga_mem_ram_MPORT_41_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_41_addr_pipe_0;
  reg  vga_mem_ram_MPORT_42_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_42_addr_pipe_0;
  reg  vga_mem_ram_MPORT_43_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_43_addr_pipe_0;
  reg  vga_mem_ram_MPORT_44_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_44_addr_pipe_0;
  reg  vga_mem_ram_MPORT_45_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_45_addr_pipe_0;
  reg  vga_mem_ram_MPORT_46_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_46_addr_pipe_0;
  reg  vga_mem_ram_MPORT_47_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_47_addr_pipe_0;
  reg  vga_mem_ram_MPORT_48_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_48_addr_pipe_0;
  reg  vga_mem_ram_MPORT_49_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_49_addr_pipe_0;
  reg  vga_mem_ram_MPORT_50_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_50_addr_pipe_0;
  reg  vga_mem_ram_MPORT_51_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_51_addr_pipe_0;
  reg  vga_mem_ram_MPORT_52_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_52_addr_pipe_0;
  reg  vga_mem_ram_MPORT_53_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_53_addr_pipe_0;
  reg  vga_mem_ram_MPORT_54_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_54_addr_pipe_0;
  reg  vga_mem_ram_MPORT_55_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_55_addr_pipe_0;
  reg  vga_mem_ram_MPORT_56_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_56_addr_pipe_0;
  reg  vga_mem_ram_MPORT_57_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_57_addr_pipe_0;
  reg  vga_mem_ram_MPORT_58_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_58_addr_pipe_0;
  reg  vga_mem_ram_MPORT_59_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_59_addr_pipe_0;
  reg  vga_mem_ram_MPORT_60_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_60_addr_pipe_0;
  reg  vga_mem_ram_MPORT_61_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_61_addr_pipe_0;
  reg  vga_mem_ram_MPORT_62_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_62_addr_pipe_0;
  reg  vga_mem_ram_MPORT_63_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_63_addr_pipe_0;
  reg  vga_mem_ram_MPORT_64_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_64_addr_pipe_0;
  reg  vga_mem_ram_MPORT_65_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_65_addr_pipe_0;
  reg  vga_mem_ram_MPORT_66_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_66_addr_pipe_0;
  reg  vga_mem_ram_MPORT_67_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_67_addr_pipe_0;
  reg  vga_mem_ram_MPORT_68_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_68_addr_pipe_0;
  reg  vga_mem_ram_MPORT_69_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_69_addr_pipe_0;
  reg  vga_mem_ram_MPORT_70_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_70_addr_pipe_0;
  reg  vga_mem_ram_MPORT_71_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_71_addr_pipe_0;
  reg  vga_mem_ram_MPORT_72_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_72_addr_pipe_0;
  reg  vga_mem_ram_MPORT_73_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_73_addr_pipe_0;
  reg  vga_mem_ram_MPORT_74_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_74_addr_pipe_0;
  reg  vga_mem_ram_MPORT_75_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_75_addr_pipe_0;
  reg  vga_mem_ram_MPORT_76_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_76_addr_pipe_0;
  reg  vga_mem_ram_MPORT_77_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_77_addr_pipe_0;
  reg  vga_mem_ram_MPORT_78_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_78_addr_pipe_0;
  reg  vga_mem_ram_MPORT_79_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_79_addr_pipe_0;
  reg  vga_mem_ram_MPORT_80_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_80_addr_pipe_0;
  reg  vga_mem_ram_MPORT_81_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_81_addr_pipe_0;
  reg  vga_mem_ram_MPORT_82_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_82_addr_pipe_0;
  reg  vga_mem_ram_MPORT_83_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_83_addr_pipe_0;
  reg  vga_mem_ram_MPORT_84_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_84_addr_pipe_0;
  reg  vga_mem_ram_MPORT_85_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_85_addr_pipe_0;
  reg  vga_mem_ram_MPORT_86_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_86_addr_pipe_0;
  reg  vga_mem_ram_MPORT_87_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_87_addr_pipe_0;
  reg  vga_mem_ram_MPORT_88_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_88_addr_pipe_0;
  reg  vga_mem_ram_MPORT_89_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_89_addr_pipe_0;
  reg  vga_mem_ram_MPORT_90_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_90_addr_pipe_0;
  reg  vga_mem_ram_MPORT_91_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_91_addr_pipe_0;
  reg  vga_mem_ram_MPORT_92_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_92_addr_pipe_0;
  reg  vga_mem_ram_MPORT_93_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_93_addr_pipe_0;
  reg  vga_mem_ram_MPORT_94_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_94_addr_pipe_0;
  reg  vga_mem_ram_MPORT_95_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_95_addr_pipe_0;
  reg  vga_mem_ram_MPORT_96_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_96_addr_pipe_0;
  reg  vga_mem_ram_MPORT_97_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_97_addr_pipe_0;
  reg  vga_mem_ram_MPORT_98_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_98_addr_pipe_0;
  reg  vga_mem_ram_MPORT_99_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_99_addr_pipe_0;
  reg  vga_mem_ram_MPORT_100_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_100_addr_pipe_0;
  reg  vga_mem_ram_MPORT_101_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_101_addr_pipe_0;
  reg  vga_mem_ram_MPORT_102_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_102_addr_pipe_0;
  reg  vga_mem_ram_MPORT_103_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_103_addr_pipe_0;
  reg  vga_mem_ram_MPORT_104_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_104_addr_pipe_0;
  reg  vga_mem_ram_MPORT_105_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_105_addr_pipe_0;
  reg  vga_mem_ram_MPORT_106_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_106_addr_pipe_0;
  reg  vga_mem_ram_MPORT_107_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_107_addr_pipe_0;
  reg  vga_mem_ram_MPORT_108_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_108_addr_pipe_0;
  reg  vga_mem_ram_MPORT_109_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_109_addr_pipe_0;
  reg  vga_mem_ram_MPORT_110_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_110_addr_pipe_0;
  reg  vga_mem_ram_MPORT_111_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_111_addr_pipe_0;
  reg  vga_mem_ram_MPORT_112_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_112_addr_pipe_0;
  reg  vga_mem_ram_MPORT_113_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_113_addr_pipe_0;
  reg  vga_mem_ram_MPORT_114_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_114_addr_pipe_0;
  reg  vga_mem_ram_MPORT_115_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_115_addr_pipe_0;
  reg  vga_mem_ram_MPORT_116_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_116_addr_pipe_0;
  reg  vga_mem_ram_MPORT_117_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_117_addr_pipe_0;
  reg  vga_mem_ram_MPORT_118_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_118_addr_pipe_0;
  reg  vga_mem_ram_MPORT_119_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_119_addr_pipe_0;
  reg  vga_mem_ram_MPORT_120_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_120_addr_pipe_0;
  reg  vga_mem_ram_MPORT_121_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_121_addr_pipe_0;
  reg  vga_mem_ram_MPORT_122_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_122_addr_pipe_0;
  reg  vga_mem_ram_MPORT_123_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_123_addr_pipe_0;
  reg  vga_mem_ram_MPORT_124_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_124_addr_pipe_0;
  reg  vga_mem_ram_MPORT_125_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_125_addr_pipe_0;
  reg  vga_mem_ram_MPORT_126_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_126_addr_pipe_0;
  reg  vga_mem_ram_MPORT_127_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_127_addr_pipe_0;
  reg  vga_mem_ram_MPORT_128_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_128_addr_pipe_0;
  reg  vga_mem_ram_MPORT_129_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_129_addr_pipe_0;
  reg  vga_mem_ram_MPORT_130_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_130_addr_pipe_0;
  reg  vga_mem_ram_MPORT_131_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_131_addr_pipe_0;
  reg  vga_mem_ram_MPORT_132_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_132_addr_pipe_0;
  reg  vga_mem_ram_MPORT_133_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_133_addr_pipe_0;
  reg  vga_mem_ram_MPORT_134_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_134_addr_pipe_0;
  reg  vga_mem_ram_MPORT_135_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_135_addr_pipe_0;
  reg  vga_mem_ram_MPORT_136_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_136_addr_pipe_0;
  reg  vga_mem_ram_MPORT_137_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_137_addr_pipe_0;
  reg  vga_mem_ram_MPORT_138_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_138_addr_pipe_0;
  reg  vga_mem_ram_MPORT_139_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_139_addr_pipe_0;
  reg  vga_mem_ram_MPORT_140_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_140_addr_pipe_0;
  reg  vga_mem_ram_MPORT_141_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_141_addr_pipe_0;
  reg  vga_mem_ram_MPORT_142_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_142_addr_pipe_0;
  reg  vga_mem_ram_MPORT_143_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_143_addr_pipe_0;
  reg  vga_mem_ram_MPORT_144_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_144_addr_pipe_0;
  reg  vga_mem_ram_MPORT_145_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_145_addr_pipe_0;
  reg  vga_mem_ram_MPORT_146_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_146_addr_pipe_0;
  reg  vga_mem_ram_MPORT_147_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_147_addr_pipe_0;
  reg  vga_mem_ram_MPORT_148_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_148_addr_pipe_0;
  reg  vga_mem_ram_MPORT_149_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_149_addr_pipe_0;
  reg  vga_mem_ram_MPORT_150_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_150_addr_pipe_0;
  reg  vga_mem_ram_MPORT_151_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_151_addr_pipe_0;
  reg  vga_mem_ram_MPORT_152_en_pipe_0;
  reg [11:0] vga_mem_ram_MPORT_152_addr_pipe_0;
  reg [287:0] ram_0; // @[vga.scala 46:20]
  reg [287:0] ram_1; // @[vga.scala 46:20]
  reg [287:0] ram_2; // @[vga.scala 46:20]
  reg [287:0] ram_3; // @[vga.scala 46:20]
  reg [287:0] ram_4; // @[vga.scala 46:20]
  reg [287:0] ram_5; // @[vga.scala 46:20]
  reg [287:0] ram_6; // @[vga.scala 46:20]
  reg [287:0] ram_7; // @[vga.scala 46:20]
  reg [287:0] ram_8; // @[vga.scala 46:20]
  reg [287:0] ram_9; // @[vga.scala 46:20]
  reg [287:0] ram_10; // @[vga.scala 46:20]
  reg [287:0] ram_11; // @[vga.scala 46:20]
  reg [287:0] ram_12; // @[vga.scala 46:20]
  reg [287:0] ram_13; // @[vga.scala 46:20]
  reg [287:0] ram_14; // @[vga.scala 46:20]
  reg [287:0] ram_15; // @[vga.scala 46:20]
  reg [287:0] ram_16; // @[vga.scala 46:20]
  reg [287:0] ram_17; // @[vga.scala 46:20]
  reg [287:0] ram_18; // @[vga.scala 46:20]
  reg [287:0] ram_19; // @[vga.scala 46:20]
  reg [287:0] ram_20; // @[vga.scala 46:20]
  reg [287:0] ram_21; // @[vga.scala 46:20]
  reg [287:0] ram_22; // @[vga.scala 46:20]
  reg [287:0] ram_23; // @[vga.scala 46:20]
  reg [287:0] ram_24; // @[vga.scala 46:20]
  reg [287:0] ram_25; // @[vga.scala 46:20]
  reg [287:0] ram_26; // @[vga.scala 46:20]
  reg [287:0] ram_27; // @[vga.scala 46:20]
  reg [287:0] ram_28; // @[vga.scala 46:20]
  reg [287:0] ram_29; // @[vga.scala 46:20]
  reg [287:0] ram_30; // @[vga.scala 46:20]
  reg [287:0] ram_31; // @[vga.scala 46:20]
  reg [287:0] ram_32; // @[vga.scala 46:20]
  reg [287:0] ram_33; // @[vga.scala 46:20]
  reg [287:0] ram_34; // @[vga.scala 46:20]
  reg [287:0] ram_35; // @[vga.scala 46:20]
  reg [287:0] ram_36; // @[vga.scala 46:20]
  reg [287:0] ram_37; // @[vga.scala 46:20]
  reg [287:0] ram_38; // @[vga.scala 46:20]
  reg [287:0] ram_39; // @[vga.scala 46:20]
  reg [287:0] ram_40; // @[vga.scala 46:20]
  reg [287:0] ram_41; // @[vga.scala 46:20]
  reg [287:0] ram_42; // @[vga.scala 46:20]
  reg [287:0] ram_43; // @[vga.scala 46:20]
  reg [287:0] ram_44; // @[vga.scala 46:20]
  reg [287:0] ram_45; // @[vga.scala 46:20]
  reg [287:0] ram_46; // @[vga.scala 46:20]
  reg [287:0] ram_47; // @[vga.scala 46:20]
  reg [287:0] ram_48; // @[vga.scala 46:20]
  reg [287:0] ram_49; // @[vga.scala 46:20]
  reg [287:0] ram_50; // @[vga.scala 46:20]
  reg [287:0] ram_51; // @[vga.scala 46:20]
  reg [287:0] ram_52; // @[vga.scala 46:20]
  reg [287:0] ram_53; // @[vga.scala 46:20]
  reg [287:0] ram_54; // @[vga.scala 46:20]
  reg [287:0] ram_55; // @[vga.scala 46:20]
  reg [287:0] ram_56; // @[vga.scala 46:20]
  reg [287:0] ram_57; // @[vga.scala 46:20]
  reg [287:0] ram_58; // @[vga.scala 46:20]
  reg [287:0] ram_59; // @[vga.scala 46:20]
  reg [287:0] ram_60; // @[vga.scala 46:20]
  reg [287:0] ram_61; // @[vga.scala 46:20]
  reg [287:0] ram_62; // @[vga.scala 46:20]
  reg [287:0] ram_63; // @[vga.scala 46:20]
  reg [287:0] ram_64; // @[vga.scala 46:20]
  reg [287:0] ram_65; // @[vga.scala 46:20]
  reg [287:0] ram_66; // @[vga.scala 46:20]
  reg [287:0] ram_67; // @[vga.scala 46:20]
  reg [287:0] ram_68; // @[vga.scala 46:20]
  reg [287:0] ram_69; // @[vga.scala 46:20]
  reg [287:0] ram_70; // @[vga.scala 46:20]
  reg [287:0] ram_71; // @[vga.scala 46:20]
  reg [287:0] ram_72; // @[vga.scala 46:20]
  reg [287:0] ram_73; // @[vga.scala 46:20]
  reg [287:0] ram_74; // @[vga.scala 46:20]
  reg [287:0] ram_75; // @[vga.scala 46:20]
  reg [287:0] ram_76; // @[vga.scala 46:20]
  reg [287:0] ram_77; // @[vga.scala 46:20]
  reg [287:0] ram_78; // @[vga.scala 46:20]
  reg [287:0] ram_79; // @[vga.scala 46:20]
  reg [287:0] ram_80; // @[vga.scala 46:20]
  reg [287:0] ram_81; // @[vga.scala 46:20]
  reg [287:0] ram_82; // @[vga.scala 46:20]
  reg [287:0] ram_83; // @[vga.scala 46:20]
  reg [287:0] ram_84; // @[vga.scala 46:20]
  reg [287:0] ram_85; // @[vga.scala 46:20]
  reg [287:0] ram_86; // @[vga.scala 46:20]
  reg [287:0] ram_87; // @[vga.scala 46:20]
  reg [287:0] ram_88; // @[vga.scala 46:20]
  reg [287:0] ram_89; // @[vga.scala 46:20]
  reg [287:0] ram_90; // @[vga.scala 46:20]
  reg [287:0] ram_91; // @[vga.scala 46:20]
  reg [287:0] ram_92; // @[vga.scala 46:20]
  reg [287:0] ram_93; // @[vga.scala 46:20]
  reg [287:0] ram_94; // @[vga.scala 46:20]
  reg [287:0] ram_95; // @[vga.scala 46:20]
  reg [287:0] ram_96; // @[vga.scala 46:20]
  reg [287:0] ram_97; // @[vga.scala 46:20]
  reg [287:0] ram_98; // @[vga.scala 46:20]
  reg [287:0] ram_99; // @[vga.scala 46:20]
  reg [287:0] ram_100; // @[vga.scala 46:20]
  reg [287:0] ram_101; // @[vga.scala 46:20]
  reg [287:0] ram_102; // @[vga.scala 46:20]
  reg [287:0] ram_103; // @[vga.scala 46:20]
  reg [287:0] ram_104; // @[vga.scala 46:20]
  reg [287:0] ram_105; // @[vga.scala 46:20]
  reg [287:0] ram_106; // @[vga.scala 46:20]
  reg [287:0] ram_107; // @[vga.scala 46:20]
  reg [287:0] ram_108; // @[vga.scala 46:20]
  reg [287:0] ram_109; // @[vga.scala 46:20]
  reg [287:0] ram_110; // @[vga.scala 46:20]
  reg [287:0] ram_111; // @[vga.scala 46:20]
  reg [287:0] ram_112; // @[vga.scala 46:20]
  reg [287:0] ram_113; // @[vga.scala 46:20]
  reg [287:0] ram_114; // @[vga.scala 46:20]
  reg [287:0] ram_115; // @[vga.scala 46:20]
  reg [287:0] ram_116; // @[vga.scala 46:20]
  reg [287:0] ram_117; // @[vga.scala 46:20]
  reg [287:0] ram_118; // @[vga.scala 46:20]
  reg [287:0] ram_119; // @[vga.scala 46:20]
  reg [287:0] ram_120; // @[vga.scala 46:20]
  reg [287:0] ram_121; // @[vga.scala 46:20]
  reg [287:0] ram_122; // @[vga.scala 46:20]
  reg [287:0] ram_123; // @[vga.scala 46:20]
  reg [287:0] ram_124; // @[vga.scala 46:20]
  reg [287:0] ram_125; // @[vga.scala 46:20]
  reg [287:0] ram_126; // @[vga.scala 46:20]
  reg [287:0] ram_127; // @[vga.scala 46:20]
  reg [287:0] ram_128; // @[vga.scala 46:20]
  reg [287:0] ram_129; // @[vga.scala 46:20]
  reg [287:0] ram_130; // @[vga.scala 46:20]
  reg [287:0] ram_131; // @[vga.scala 46:20]
  reg [287:0] ram_132; // @[vga.scala 46:20]
  reg [287:0] ram_133; // @[vga.scala 46:20]
  reg [287:0] ram_134; // @[vga.scala 46:20]
  reg [287:0] ram_135; // @[vga.scala 46:20]
  reg [287:0] ram_136; // @[vga.scala 46:20]
  reg [287:0] ram_137; // @[vga.scala 46:20]
  reg [287:0] ram_138; // @[vga.scala 46:20]
  reg [287:0] ram_139; // @[vga.scala 46:20]
  reg [287:0] ram_140; // @[vga.scala 46:20]
  reg [287:0] ram_141; // @[vga.scala 46:20]
  reg [287:0] ram_142; // @[vga.scala 46:20]
  reg [287:0] ram_143; // @[vga.scala 46:20]
  reg [287:0] ram_144; // @[vga.scala 46:20]
  reg [287:0] ram_145; // @[vga.scala 46:20]
  reg [287:0] ram_146; // @[vga.scala 46:20]
  reg [287:0] ram_147; // @[vga.scala 46:20]
  reg [287:0] ram_148; // @[vga.scala 46:20]
  reg [287:0] ram_149; // @[vga.scala 46:20]
  reg [287:0] ram_150; // @[vga.scala 46:20]
  reg [287:0] ram_151; // @[vga.scala 46:20]
  reg [287:0] ram_152; // @[vga.scala 46:20]
  reg [287:0] ram_153; // @[vga.scala 46:20]
  reg [287:0] ram_154; // @[vga.scala 46:20]
  reg [287:0] ram_155; // @[vga.scala 46:20]
  reg [287:0] ram_156; // @[vga.scala 46:20]
  reg [287:0] ram_157; // @[vga.scala 46:20]
  reg [287:0] ram_158; // @[vga.scala 46:20]
  reg [287:0] ram_159; // @[vga.scala 46:20]
  reg [287:0] ram_160; // @[vga.scala 46:20]
  reg [287:0] ram_161; // @[vga.scala 46:20]
  reg [287:0] ram_162; // @[vga.scala 46:20]
  reg [287:0] ram_163; // @[vga.scala 46:20]
  reg [287:0] ram_164; // @[vga.scala 46:20]
  reg [287:0] ram_165; // @[vga.scala 46:20]
  reg [287:0] ram_166; // @[vga.scala 46:20]
  reg [287:0] ram_167; // @[vga.scala 46:20]
  reg [287:0] ram_168; // @[vga.scala 46:20]
  reg [287:0] ram_169; // @[vga.scala 46:20]
  reg [287:0] ram_170; // @[vga.scala 46:20]
  reg [287:0] ram_171; // @[vga.scala 46:20]
  reg [287:0] ram_172; // @[vga.scala 46:20]
  reg [287:0] ram_173; // @[vga.scala 46:20]
  reg [287:0] ram_174; // @[vga.scala 46:20]
  reg [287:0] ram_175; // @[vga.scala 46:20]
  reg [287:0] ram_176; // @[vga.scala 46:20]
  reg [287:0] ram_177; // @[vga.scala 46:20]
  reg [287:0] ram_178; // @[vga.scala 46:20]
  reg [287:0] ram_179; // @[vga.scala 46:20]
  reg [287:0] ram_180; // @[vga.scala 46:20]
  reg [287:0] ram_181; // @[vga.scala 46:20]
  reg [287:0] ram_182; // @[vga.scala 46:20]
  reg [287:0] ram_183; // @[vga.scala 46:20]
  reg [287:0] ram_184; // @[vga.scala 46:20]
  reg [287:0] ram_185; // @[vga.scala 46:20]
  reg [287:0] ram_186; // @[vga.scala 46:20]
  reg [287:0] ram_187; // @[vga.scala 46:20]
  reg [287:0] ram_188; // @[vga.scala 46:20]
  reg [287:0] ram_189; // @[vga.scala 46:20]
  reg [287:0] ram_190; // @[vga.scala 46:20]
  reg [287:0] ram_191; // @[vga.scala 46:20]
  reg [287:0] ram_192; // @[vga.scala 46:20]
  reg [287:0] ram_193; // @[vga.scala 46:20]
  reg [287:0] ram_194; // @[vga.scala 46:20]
  reg [287:0] ram_195; // @[vga.scala 46:20]
  reg [287:0] ram_196; // @[vga.scala 46:20]
  reg [287:0] ram_197; // @[vga.scala 46:20]
  reg [287:0] ram_198; // @[vga.scala 46:20]
  reg [287:0] ram_199; // @[vga.scala 46:20]
  reg [287:0] ram_200; // @[vga.scala 46:20]
  reg [287:0] ram_201; // @[vga.scala 46:20]
  reg [287:0] ram_202; // @[vga.scala 46:20]
  reg [287:0] ram_203; // @[vga.scala 46:20]
  reg [287:0] ram_204; // @[vga.scala 46:20]
  reg [287:0] ram_205; // @[vga.scala 46:20]
  reg [287:0] ram_206; // @[vga.scala 46:20]
  reg [287:0] ram_207; // @[vga.scala 46:20]
  reg [287:0] ram_208; // @[vga.scala 46:20]
  reg [287:0] ram_209; // @[vga.scala 46:20]
  reg [287:0] ram_210; // @[vga.scala 46:20]
  reg [287:0] ram_211; // @[vga.scala 46:20]
  reg [287:0] ram_212; // @[vga.scala 46:20]
  reg [287:0] ram_213; // @[vga.scala 46:20]
  reg [287:0] ram_214; // @[vga.scala 46:20]
  reg [287:0] ram_215; // @[vga.scala 46:20]
  reg [287:0] ram_216; // @[vga.scala 46:20]
  reg [287:0] ram_217; // @[vga.scala 46:20]
  reg [287:0] ram_218; // @[vga.scala 46:20]
  reg [287:0] ram_219; // @[vga.scala 46:20]
  reg [287:0] ram_220; // @[vga.scala 46:20]
  reg [287:0] ram_221; // @[vga.scala 46:20]
  reg [287:0] ram_222; // @[vga.scala 46:20]
  reg [287:0] ram_223; // @[vga.scala 46:20]
  reg [287:0] ram_224; // @[vga.scala 46:20]
  reg [287:0] ram_225; // @[vga.scala 46:20]
  reg [287:0] ram_226; // @[vga.scala 46:20]
  reg [287:0] ram_227; // @[vga.scala 46:20]
  reg [287:0] ram_228; // @[vga.scala 46:20]
  reg [287:0] ram_229; // @[vga.scala 46:20]
  reg [287:0] ram_230; // @[vga.scala 46:20]
  reg [287:0] ram_231; // @[vga.scala 46:20]
  reg [287:0] ram_232; // @[vga.scala 46:20]
  reg [287:0] ram_233; // @[vga.scala 46:20]
  reg [287:0] ram_234; // @[vga.scala 46:20]
  reg [287:0] ram_235; // @[vga.scala 46:20]
  reg [287:0] ram_236; // @[vga.scala 46:20]
  reg [287:0] ram_237; // @[vga.scala 46:20]
  reg [287:0] ram_238; // @[vga.scala 46:20]
  reg [287:0] ram_239; // @[vga.scala 46:20]
  reg [287:0] ram_240; // @[vga.scala 46:20]
  reg [287:0] ram_241; // @[vga.scala 46:20]
  reg [287:0] ram_242; // @[vga.scala 46:20]
  reg [287:0] ram_243; // @[vga.scala 46:20]
  reg [287:0] ram_244; // @[vga.scala 46:20]
  reg [287:0] ram_245; // @[vga.scala 46:20]
  reg [287:0] ram_246; // @[vga.scala 46:20]
  reg [287:0] ram_247; // @[vga.scala 46:20]
  reg [287:0] ram_248; // @[vga.scala 46:20]
  reg [287:0] ram_249; // @[vga.scala 46:20]
  reg [287:0] ram_250; // @[vga.scala 46:20]
  reg [287:0] ram_251; // @[vga.scala 46:20]
  reg [287:0] ram_252; // @[vga.scala 46:20]
  reg [287:0] ram_253; // @[vga.scala 46:20]
  reg [287:0] ram_254; // @[vga.scala 46:20]
  reg [287:0] ram_255; // @[vga.scala 46:20]
  reg [287:0] ram_256; // @[vga.scala 46:20]
  reg [287:0] ram_257; // @[vga.scala 46:20]
  reg [287:0] ram_258; // @[vga.scala 46:20]
  reg [287:0] ram_259; // @[vga.scala 46:20]
  reg [287:0] ram_260; // @[vga.scala 46:20]
  reg [287:0] ram_261; // @[vga.scala 46:20]
  reg [287:0] ram_262; // @[vga.scala 46:20]
  reg [287:0] ram_263; // @[vga.scala 46:20]
  reg [287:0] ram_264; // @[vga.scala 46:20]
  reg [287:0] ram_265; // @[vga.scala 46:20]
  reg [287:0] ram_266; // @[vga.scala 46:20]
  reg [287:0] ram_267; // @[vga.scala 46:20]
  reg [287:0] ram_268; // @[vga.scala 46:20]
  reg [287:0] ram_269; // @[vga.scala 46:20]
  reg [287:0] ram_270; // @[vga.scala 46:20]
  reg [287:0] ram_271; // @[vga.scala 46:20]
  reg [287:0] ram_272; // @[vga.scala 46:20]
  reg [287:0] ram_273; // @[vga.scala 46:20]
  reg [287:0] ram_274; // @[vga.scala 46:20]
  reg [287:0] ram_275; // @[vga.scala 46:20]
  reg [287:0] ram_276; // @[vga.scala 46:20]
  reg [287:0] ram_277; // @[vga.scala 46:20]
  reg [287:0] ram_278; // @[vga.scala 46:20]
  reg [287:0] ram_279; // @[vga.scala 46:20]
  reg [287:0] ram_280; // @[vga.scala 46:20]
  reg [287:0] ram_281; // @[vga.scala 46:20]
  reg [287:0] ram_282; // @[vga.scala 46:20]
  reg [287:0] ram_283; // @[vga.scala 46:20]
  reg [287:0] ram_284; // @[vga.scala 46:20]
  reg [287:0] ram_285; // @[vga.scala 46:20]
  reg [287:0] ram_286; // @[vga.scala 46:20]
  reg [287:0] ram_287; // @[vga.scala 46:20]
  reg [287:0] ram_288; // @[vga.scala 46:20]
  reg [287:0] ram_289; // @[vga.scala 46:20]
  reg [287:0] ram_290; // @[vga.scala 46:20]
  reg [287:0] ram_291; // @[vga.scala 46:20]
  reg [287:0] ram_292; // @[vga.scala 46:20]
  reg [287:0] ram_293; // @[vga.scala 46:20]
  reg [287:0] ram_294; // @[vga.scala 46:20]
  reg [287:0] ram_295; // @[vga.scala 46:20]
  reg [287:0] ram_296; // @[vga.scala 46:20]
  reg [287:0] ram_297; // @[vga.scala 46:20]
  reg [287:0] ram_298; // @[vga.scala 46:20]
  reg [287:0] ram_299; // @[vga.scala 46:20]
  reg [287:0] ram_300; // @[vga.scala 46:20]
  reg [287:0] ram_301; // @[vga.scala 46:20]
  reg [287:0] ram_302; // @[vga.scala 46:20]
  reg [287:0] ram_303; // @[vga.scala 46:20]
  reg [287:0] ram_304; // @[vga.scala 46:20]
  reg [287:0] ram_305; // @[vga.scala 46:20]
  reg [287:0] ram_306; // @[vga.scala 46:20]
  reg [287:0] ram_307; // @[vga.scala 46:20]
  reg [287:0] ram_308; // @[vga.scala 46:20]
  reg [287:0] ram_309; // @[vga.scala 46:20]
  reg [287:0] ram_310; // @[vga.scala 46:20]
  reg [287:0] ram_311; // @[vga.scala 46:20]
  reg [287:0] ram_312; // @[vga.scala 46:20]
  reg [287:0] ram_313; // @[vga.scala 46:20]
  reg [287:0] ram_314; // @[vga.scala 46:20]
  reg [287:0] ram_315; // @[vga.scala 46:20]
  reg [287:0] ram_316; // @[vga.scala 46:20]
  reg [287:0] ram_317; // @[vga.scala 46:20]
  reg [287:0] ram_318; // @[vga.scala 46:20]
  reg [287:0] ram_319; // @[vga.scala 46:20]
  reg [287:0] ram_320; // @[vga.scala 46:20]
  reg [287:0] ram_321; // @[vga.scala 46:20]
  reg [287:0] ram_322; // @[vga.scala 46:20]
  reg [287:0] ram_323; // @[vga.scala 46:20]
  reg [287:0] ram_324; // @[vga.scala 46:20]
  reg [287:0] ram_325; // @[vga.scala 46:20]
  reg [287:0] ram_326; // @[vga.scala 46:20]
  reg [287:0] ram_327; // @[vga.scala 46:20]
  reg [287:0] ram_328; // @[vga.scala 46:20]
  reg [287:0] ram_329; // @[vga.scala 46:20]
  reg [287:0] ram_330; // @[vga.scala 46:20]
  reg [287:0] ram_331; // @[vga.scala 46:20]
  reg [287:0] ram_332; // @[vga.scala 46:20]
  reg [287:0] ram_333; // @[vga.scala 46:20]
  reg [287:0] ram_334; // @[vga.scala 46:20]
  reg [287:0] ram_335; // @[vga.scala 46:20]
  reg [287:0] ram_336; // @[vga.scala 46:20]
  reg [287:0] ram_337; // @[vga.scala 46:20]
  reg [287:0] ram_338; // @[vga.scala 46:20]
  reg [287:0] ram_339; // @[vga.scala 46:20]
  reg [287:0] ram_340; // @[vga.scala 46:20]
  reg [287:0] ram_341; // @[vga.scala 46:20]
  reg [287:0] ram_342; // @[vga.scala 46:20]
  reg [287:0] ram_343; // @[vga.scala 46:20]
  reg [287:0] ram_344; // @[vga.scala 46:20]
  reg [287:0] ram_345; // @[vga.scala 46:20]
  reg [287:0] ram_346; // @[vga.scala 46:20]
  reg [287:0] ram_347; // @[vga.scala 46:20]
  reg [287:0] ram_348; // @[vga.scala 46:20]
  reg [287:0] ram_349; // @[vga.scala 46:20]
  reg [287:0] ram_350; // @[vga.scala 46:20]
  reg [287:0] ram_351; // @[vga.scala 46:20]
  reg [287:0] ram_352; // @[vga.scala 46:20]
  reg [287:0] ram_353; // @[vga.scala 46:20]
  reg [287:0] ram_354; // @[vga.scala 46:20]
  reg [287:0] ram_355; // @[vga.scala 46:20]
  reg [287:0] ram_356; // @[vga.scala 46:20]
  reg [287:0] ram_357; // @[vga.scala 46:20]
  reg [287:0] ram_358; // @[vga.scala 46:20]
  reg [287:0] ram_359; // @[vga.scala 46:20]
  reg [287:0] ram_360; // @[vga.scala 46:20]
  reg [287:0] ram_361; // @[vga.scala 46:20]
  reg [287:0] ram_362; // @[vga.scala 46:20]
  reg [287:0] ram_363; // @[vga.scala 46:20]
  reg [287:0] ram_364; // @[vga.scala 46:20]
  reg [287:0] ram_365; // @[vga.scala 46:20]
  reg [287:0] ram_366; // @[vga.scala 46:20]
  reg [287:0] ram_367; // @[vga.scala 46:20]
  reg [287:0] ram_368; // @[vga.scala 46:20]
  reg [287:0] ram_369; // @[vga.scala 46:20]
  reg [287:0] ram_370; // @[vga.scala 46:20]
  reg [287:0] ram_371; // @[vga.scala 46:20]
  reg [287:0] ram_372; // @[vga.scala 46:20]
  reg [287:0] ram_373; // @[vga.scala 46:20]
  reg [287:0] ram_374; // @[vga.scala 46:20]
  reg [287:0] ram_375; // @[vga.scala 46:20]
  reg [287:0] ram_376; // @[vga.scala 46:20]
  reg [287:0] ram_377; // @[vga.scala 46:20]
  reg [287:0] ram_378; // @[vga.scala 46:20]
  reg [287:0] ram_379; // @[vga.scala 46:20]
  reg [287:0] ram_380; // @[vga.scala 46:20]
  reg [287:0] ram_381; // @[vga.scala 46:20]
  reg [287:0] ram_382; // @[vga.scala 46:20]
  reg [287:0] ram_383; // @[vga.scala 46:20]
  reg [287:0] ram_384; // @[vga.scala 46:20]
  reg [287:0] ram_385; // @[vga.scala 46:20]
  reg [287:0] ram_386; // @[vga.scala 46:20]
  reg [287:0] ram_387; // @[vga.scala 46:20]
  reg [287:0] ram_388; // @[vga.scala 46:20]
  reg [287:0] ram_389; // @[vga.scala 46:20]
  reg [287:0] ram_390; // @[vga.scala 46:20]
  reg [287:0] ram_391; // @[vga.scala 46:20]
  reg [287:0] ram_392; // @[vga.scala 46:20]
  reg [287:0] ram_393; // @[vga.scala 46:20]
  reg [287:0] ram_394; // @[vga.scala 46:20]
  reg [287:0] ram_395; // @[vga.scala 46:20]
  reg [287:0] ram_396; // @[vga.scala 46:20]
  reg [287:0] ram_397; // @[vga.scala 46:20]
  reg [287:0] ram_398; // @[vga.scala 46:20]
  reg [287:0] ram_399; // @[vga.scala 46:20]
  reg [287:0] ram_400; // @[vga.scala 46:20]
  reg [287:0] ram_401; // @[vga.scala 46:20]
  reg [287:0] ram_402; // @[vga.scala 46:20]
  reg [287:0] ram_403; // @[vga.scala 46:20]
  reg [287:0] ram_404; // @[vga.scala 46:20]
  reg [287:0] ram_405; // @[vga.scala 46:20]
  reg [287:0] ram_406; // @[vga.scala 46:20]
  reg [287:0] ram_407; // @[vga.scala 46:20]
  reg [287:0] ram_408; // @[vga.scala 46:20]
  reg [287:0] ram_409; // @[vga.scala 46:20]
  reg [287:0] ram_410; // @[vga.scala 46:20]
  reg [287:0] ram_411; // @[vga.scala 46:20]
  reg [287:0] ram_412; // @[vga.scala 46:20]
  reg [287:0] ram_413; // @[vga.scala 46:20]
  reg [287:0] ram_414; // @[vga.scala 46:20]
  reg [287:0] ram_415; // @[vga.scala 46:20]
  reg [287:0] ram_416; // @[vga.scala 46:20]
  reg [287:0] ram_417; // @[vga.scala 46:20]
  reg [287:0] ram_418; // @[vga.scala 46:20]
  reg [287:0] ram_419; // @[vga.scala 46:20]
  reg [287:0] ram_420; // @[vga.scala 46:20]
  reg [287:0] ram_421; // @[vga.scala 46:20]
  reg [287:0] ram_422; // @[vga.scala 46:20]
  reg [287:0] ram_423; // @[vga.scala 46:20]
  reg [287:0] ram_424; // @[vga.scala 46:20]
  reg [287:0] ram_425; // @[vga.scala 46:20]
  reg [287:0] ram_426; // @[vga.scala 46:20]
  reg [287:0] ram_427; // @[vga.scala 46:20]
  reg [287:0] ram_428; // @[vga.scala 46:20]
  reg [287:0] ram_429; // @[vga.scala 46:20]
  reg [287:0] ram_430; // @[vga.scala 46:20]
  reg [287:0] ram_431; // @[vga.scala 46:20]
  reg [287:0] ram_432; // @[vga.scala 46:20]
  reg [287:0] ram_433; // @[vga.scala 46:20]
  reg [287:0] ram_434; // @[vga.scala 46:20]
  reg [287:0] ram_435; // @[vga.scala 46:20]
  reg [287:0] ram_436; // @[vga.scala 46:20]
  reg [287:0] ram_437; // @[vga.scala 46:20]
  reg [287:0] ram_438; // @[vga.scala 46:20]
  reg [287:0] ram_439; // @[vga.scala 46:20]
  reg [287:0] ram_440; // @[vga.scala 46:20]
  reg [287:0] ram_441; // @[vga.scala 46:20]
  reg [287:0] ram_442; // @[vga.scala 46:20]
  reg [287:0] ram_443; // @[vga.scala 46:20]
  reg [287:0] ram_444; // @[vga.scala 46:20]
  reg [287:0] ram_445; // @[vga.scala 46:20]
  reg [287:0] ram_446; // @[vga.scala 46:20]
  reg [287:0] ram_447; // @[vga.scala 46:20]
  reg [287:0] ram_448; // @[vga.scala 46:20]
  reg [287:0] ram_449; // @[vga.scala 46:20]
  reg [287:0] ram_450; // @[vga.scala 46:20]
  reg [287:0] ram_451; // @[vga.scala 46:20]
  reg [287:0] ram_452; // @[vga.scala 46:20]
  reg [287:0] ram_453; // @[vga.scala 46:20]
  reg [287:0] ram_454; // @[vga.scala 46:20]
  reg [287:0] ram_455; // @[vga.scala 46:20]
  reg [287:0] ram_456; // @[vga.scala 46:20]
  reg [287:0] ram_457; // @[vga.scala 46:20]
  reg [287:0] ram_458; // @[vga.scala 46:20]
  reg [287:0] ram_459; // @[vga.scala 46:20]
  reg [287:0] ram_460; // @[vga.scala 46:20]
  reg [287:0] ram_461; // @[vga.scala 46:20]
  reg [287:0] ram_462; // @[vga.scala 46:20]
  reg [287:0] ram_463; // @[vga.scala 46:20]
  reg [287:0] ram_464; // @[vga.scala 46:20]
  reg [287:0] ram_465; // @[vga.scala 46:20]
  reg [287:0] ram_466; // @[vga.scala 46:20]
  reg [287:0] ram_467; // @[vga.scala 46:20]
  reg [287:0] ram_468; // @[vga.scala 46:20]
  reg [287:0] ram_469; // @[vga.scala 46:20]
  reg [287:0] ram_470; // @[vga.scala 46:20]
  reg [287:0] ram_471; // @[vga.scala 46:20]
  reg [287:0] ram_472; // @[vga.scala 46:20]
  reg [287:0] ram_473; // @[vga.scala 46:20]
  reg [287:0] ram_474; // @[vga.scala 46:20]
  reg [287:0] ram_475; // @[vga.scala 46:20]
  reg [287:0] ram_476; // @[vga.scala 46:20]
  reg [287:0] ram_477; // @[vga.scala 46:20]
  reg [287:0] ram_478; // @[vga.scala 46:20]
  reg [287:0] ram_479; // @[vga.scala 46:20]
  reg [287:0] ram_480; // @[vga.scala 46:20]
  reg [287:0] ram_481; // @[vga.scala 46:20]
  reg [287:0] ram_482; // @[vga.scala 46:20]
  reg [287:0] ram_483; // @[vga.scala 46:20]
  reg [287:0] ram_484; // @[vga.scala 46:20]
  reg [287:0] ram_485; // @[vga.scala 46:20]
  reg [287:0] ram_486; // @[vga.scala 46:20]
  reg [287:0] ram_487; // @[vga.scala 46:20]
  reg [287:0] ram_488; // @[vga.scala 46:20]
  reg [287:0] ram_489; // @[vga.scala 46:20]
  reg [287:0] ram_490; // @[vga.scala 46:20]
  reg [287:0] ram_491; // @[vga.scala 46:20]
  reg [287:0] ram_492; // @[vga.scala 46:20]
  reg [287:0] ram_493; // @[vga.scala 46:20]
  reg [287:0] ram_494; // @[vga.scala 46:20]
  reg [287:0] ram_495; // @[vga.scala 46:20]
  reg [287:0] ram_496; // @[vga.scala 46:20]
  reg [287:0] ram_497; // @[vga.scala 46:20]
  reg [287:0] ram_498; // @[vga.scala 46:20]
  reg [287:0] ram_499; // @[vga.scala 46:20]
  reg [287:0] ram_500; // @[vga.scala 46:20]
  reg [287:0] ram_501; // @[vga.scala 46:20]
  reg [287:0] ram_502; // @[vga.scala 46:20]
  reg [287:0] ram_503; // @[vga.scala 46:20]
  reg [287:0] ram_504; // @[vga.scala 46:20]
  reg [287:0] ram_505; // @[vga.scala 46:20]
  reg [287:0] ram_506; // @[vga.scala 46:20]
  reg [287:0] ram_507; // @[vga.scala 46:20]
  reg [287:0] ram_508; // @[vga.scala 46:20]
  reg [287:0] ram_509; // @[vga.scala 46:20]
  reg [287:0] ram_510; // @[vga.scala 46:20]
  reg [287:0] ram_511; // @[vga.scala 46:20]
  reg [287:0] ram_512; // @[vga.scala 46:20]
  reg [287:0] ram_513; // @[vga.scala 46:20]
  reg [287:0] ram_514; // @[vga.scala 46:20]
  reg [287:0] ram_515; // @[vga.scala 46:20]
  reg [287:0] ram_516; // @[vga.scala 46:20]
  reg [287:0] ram_517; // @[vga.scala 46:20]
  reg [287:0] ram_518; // @[vga.scala 46:20]
  reg [287:0] ram_519; // @[vga.scala 46:20]
  reg [287:0] ram_520; // @[vga.scala 46:20]
  reg [287:0] ram_521; // @[vga.scala 46:20]
  reg [287:0] ram_522; // @[vga.scala 46:20]
  reg [287:0] ram_523; // @[vga.scala 46:20]
  reg [287:0] ram_524; // @[vga.scala 46:20]
  reg [9:0] h; // @[vga.scala 47:18]
  reg [8:0] v; // @[vga.scala 48:18]
  wire  _T_1 = v == 9'h120; // @[vga.scala 54:25]
  wire [9:0] _h_T_1 = h + 10'h10; // @[vga.scala 57:13]
  wire [10:0] _T_6 = {{1'd0}, h}; // @[vga.scala 64:14]
  wire [12:0] _ram_T_2 = 5'h10 * io_ascii; // @[vga.scala 64:73]
  wire  ram_hi_hi_hi_lo = vga_mem_ram_MPORT_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo = vga_mem_ram_MPORT_1_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi = vga_mem_ram_MPORT_2_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo = vga_mem_ram_MPORT_3_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi = vga_mem_ram_MPORT_4_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo = vga_mem_ram_MPORT_5_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo = vga_mem_ram_MPORT_6_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi = vga_mem_ram_MPORT_7_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo = vga_mem_ram_MPORT_8_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_20 = {278'h0,ram_hi_hi_hi_lo,ram_hi_hi_lo,ram_hi_lo_hi,ram_hi_lo_lo,ram_lo_hi_hi_hi,
    ram_lo_hi_hi_lo,ram_lo_hi_lo,ram_lo_lo_hi,ram_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [12:0] _ram_T_21 = v * 4'h9; // @[vga.scala 64:305]
  wire [12:0] _ram_T_23 = 13'h116 - _ram_T_21; // @[vga.scala 64:303]
  wire [8477:0] _GEN_19060 = {{8191'd0}, _ram_T_20}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_24 = _GEN_19060 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_4 = 10'h1 == _T_6[9:0] ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5 = 10'h2 == _T_6[9:0] ? ram_2 : _GEN_4; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6 = 10'h3 == _T_6[9:0] ? ram_3 : _GEN_5; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7 = 10'h4 == _T_6[9:0] ? ram_4 : _GEN_6; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8 = 10'h5 == _T_6[9:0] ? ram_5 : _GEN_7; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9 = 10'h6 == _T_6[9:0] ? ram_6 : _GEN_8; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10 = 10'h7 == _T_6[9:0] ? ram_7 : _GEN_9; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11 = 10'h8 == _T_6[9:0] ? ram_8 : _GEN_10; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12 = 10'h9 == _T_6[9:0] ? ram_9 : _GEN_11; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13 = 10'ha == _T_6[9:0] ? ram_10 : _GEN_12; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14 = 10'hb == _T_6[9:0] ? ram_11 : _GEN_13; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15 = 10'hc == _T_6[9:0] ? ram_12 : _GEN_14; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16 = 10'hd == _T_6[9:0] ? ram_13 : _GEN_15; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17 = 10'he == _T_6[9:0] ? ram_14 : _GEN_16; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_18 = 10'hf == _T_6[9:0] ? ram_15 : _GEN_17; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_19 = 10'h10 == _T_6[9:0] ? ram_16 : _GEN_18; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_20 = 10'h11 == _T_6[9:0] ? ram_17 : _GEN_19; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_21 = 10'h12 == _T_6[9:0] ? ram_18 : _GEN_20; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_22 = 10'h13 == _T_6[9:0] ? ram_19 : _GEN_21; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_23 = 10'h14 == _T_6[9:0] ? ram_20 : _GEN_22; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_24 = 10'h15 == _T_6[9:0] ? ram_21 : _GEN_23; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_25 = 10'h16 == _T_6[9:0] ? ram_22 : _GEN_24; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_26 = 10'h17 == _T_6[9:0] ? ram_23 : _GEN_25; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_27 = 10'h18 == _T_6[9:0] ? ram_24 : _GEN_26; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_28 = 10'h19 == _T_6[9:0] ? ram_25 : _GEN_27; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_29 = 10'h1a == _T_6[9:0] ? ram_26 : _GEN_28; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_30 = 10'h1b == _T_6[9:0] ? ram_27 : _GEN_29; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_31 = 10'h1c == _T_6[9:0] ? ram_28 : _GEN_30; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_32 = 10'h1d == _T_6[9:0] ? ram_29 : _GEN_31; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_33 = 10'h1e == _T_6[9:0] ? ram_30 : _GEN_32; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_34 = 10'h1f == _T_6[9:0] ? ram_31 : _GEN_33; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_35 = 10'h20 == _T_6[9:0] ? ram_32 : _GEN_34; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_36 = 10'h21 == _T_6[9:0] ? ram_33 : _GEN_35; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_37 = 10'h22 == _T_6[9:0] ? ram_34 : _GEN_36; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_38 = 10'h23 == _T_6[9:0] ? ram_35 : _GEN_37; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_39 = 10'h24 == _T_6[9:0] ? ram_36 : _GEN_38; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_40 = 10'h25 == _T_6[9:0] ? ram_37 : _GEN_39; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_41 = 10'h26 == _T_6[9:0] ? ram_38 : _GEN_40; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_42 = 10'h27 == _T_6[9:0] ? ram_39 : _GEN_41; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_43 = 10'h28 == _T_6[9:0] ? ram_40 : _GEN_42; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_44 = 10'h29 == _T_6[9:0] ? ram_41 : _GEN_43; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_45 = 10'h2a == _T_6[9:0] ? ram_42 : _GEN_44; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_46 = 10'h2b == _T_6[9:0] ? ram_43 : _GEN_45; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_47 = 10'h2c == _T_6[9:0] ? ram_44 : _GEN_46; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_48 = 10'h2d == _T_6[9:0] ? ram_45 : _GEN_47; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_49 = 10'h2e == _T_6[9:0] ? ram_46 : _GEN_48; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_50 = 10'h2f == _T_6[9:0] ? ram_47 : _GEN_49; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_51 = 10'h30 == _T_6[9:0] ? ram_48 : _GEN_50; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_52 = 10'h31 == _T_6[9:0] ? ram_49 : _GEN_51; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_53 = 10'h32 == _T_6[9:0] ? ram_50 : _GEN_52; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_54 = 10'h33 == _T_6[9:0] ? ram_51 : _GEN_53; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_55 = 10'h34 == _T_6[9:0] ? ram_52 : _GEN_54; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_56 = 10'h35 == _T_6[9:0] ? ram_53 : _GEN_55; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_57 = 10'h36 == _T_6[9:0] ? ram_54 : _GEN_56; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_58 = 10'h37 == _T_6[9:0] ? ram_55 : _GEN_57; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_59 = 10'h38 == _T_6[9:0] ? ram_56 : _GEN_58; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_60 = 10'h39 == _T_6[9:0] ? ram_57 : _GEN_59; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_61 = 10'h3a == _T_6[9:0] ? ram_58 : _GEN_60; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_62 = 10'h3b == _T_6[9:0] ? ram_59 : _GEN_61; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_63 = 10'h3c == _T_6[9:0] ? ram_60 : _GEN_62; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_64 = 10'h3d == _T_6[9:0] ? ram_61 : _GEN_63; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_65 = 10'h3e == _T_6[9:0] ? ram_62 : _GEN_64; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_66 = 10'h3f == _T_6[9:0] ? ram_63 : _GEN_65; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_67 = 10'h40 == _T_6[9:0] ? ram_64 : _GEN_66; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_68 = 10'h41 == _T_6[9:0] ? ram_65 : _GEN_67; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_69 = 10'h42 == _T_6[9:0] ? ram_66 : _GEN_68; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_70 = 10'h43 == _T_6[9:0] ? ram_67 : _GEN_69; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_71 = 10'h44 == _T_6[9:0] ? ram_68 : _GEN_70; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_72 = 10'h45 == _T_6[9:0] ? ram_69 : _GEN_71; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_73 = 10'h46 == _T_6[9:0] ? ram_70 : _GEN_72; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_74 = 10'h47 == _T_6[9:0] ? ram_71 : _GEN_73; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_75 = 10'h48 == _T_6[9:0] ? ram_72 : _GEN_74; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_76 = 10'h49 == _T_6[9:0] ? ram_73 : _GEN_75; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_77 = 10'h4a == _T_6[9:0] ? ram_74 : _GEN_76; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_78 = 10'h4b == _T_6[9:0] ? ram_75 : _GEN_77; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_79 = 10'h4c == _T_6[9:0] ? ram_76 : _GEN_78; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_80 = 10'h4d == _T_6[9:0] ? ram_77 : _GEN_79; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_81 = 10'h4e == _T_6[9:0] ? ram_78 : _GEN_80; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_82 = 10'h4f == _T_6[9:0] ? ram_79 : _GEN_81; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_83 = 10'h50 == _T_6[9:0] ? ram_80 : _GEN_82; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_84 = 10'h51 == _T_6[9:0] ? ram_81 : _GEN_83; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_85 = 10'h52 == _T_6[9:0] ? ram_82 : _GEN_84; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_86 = 10'h53 == _T_6[9:0] ? ram_83 : _GEN_85; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_87 = 10'h54 == _T_6[9:0] ? ram_84 : _GEN_86; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_88 = 10'h55 == _T_6[9:0] ? ram_85 : _GEN_87; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_89 = 10'h56 == _T_6[9:0] ? ram_86 : _GEN_88; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_90 = 10'h57 == _T_6[9:0] ? ram_87 : _GEN_89; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_91 = 10'h58 == _T_6[9:0] ? ram_88 : _GEN_90; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_92 = 10'h59 == _T_6[9:0] ? ram_89 : _GEN_91; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_93 = 10'h5a == _T_6[9:0] ? ram_90 : _GEN_92; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_94 = 10'h5b == _T_6[9:0] ? ram_91 : _GEN_93; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_95 = 10'h5c == _T_6[9:0] ? ram_92 : _GEN_94; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_96 = 10'h5d == _T_6[9:0] ? ram_93 : _GEN_95; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_97 = 10'h5e == _T_6[9:0] ? ram_94 : _GEN_96; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_98 = 10'h5f == _T_6[9:0] ? ram_95 : _GEN_97; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_99 = 10'h60 == _T_6[9:0] ? ram_96 : _GEN_98; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_100 = 10'h61 == _T_6[9:0] ? ram_97 : _GEN_99; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_101 = 10'h62 == _T_6[9:0] ? ram_98 : _GEN_100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_102 = 10'h63 == _T_6[9:0] ? ram_99 : _GEN_101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_103 = 10'h64 == _T_6[9:0] ? ram_100 : _GEN_102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_104 = 10'h65 == _T_6[9:0] ? ram_101 : _GEN_103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_105 = 10'h66 == _T_6[9:0] ? ram_102 : _GEN_104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_106 = 10'h67 == _T_6[9:0] ? ram_103 : _GEN_105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_107 = 10'h68 == _T_6[9:0] ? ram_104 : _GEN_106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_108 = 10'h69 == _T_6[9:0] ? ram_105 : _GEN_107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_109 = 10'h6a == _T_6[9:0] ? ram_106 : _GEN_108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_110 = 10'h6b == _T_6[9:0] ? ram_107 : _GEN_109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_111 = 10'h6c == _T_6[9:0] ? ram_108 : _GEN_110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_112 = 10'h6d == _T_6[9:0] ? ram_109 : _GEN_111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_113 = 10'h6e == _T_6[9:0] ? ram_110 : _GEN_112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_114 = 10'h6f == _T_6[9:0] ? ram_111 : _GEN_113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_115 = 10'h70 == _T_6[9:0] ? ram_112 : _GEN_114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_116 = 10'h71 == _T_6[9:0] ? ram_113 : _GEN_115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_117 = 10'h72 == _T_6[9:0] ? ram_114 : _GEN_116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_118 = 10'h73 == _T_6[9:0] ? ram_115 : _GEN_117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_119 = 10'h74 == _T_6[9:0] ? ram_116 : _GEN_118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_120 = 10'h75 == _T_6[9:0] ? ram_117 : _GEN_119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_121 = 10'h76 == _T_6[9:0] ? ram_118 : _GEN_120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_122 = 10'h77 == _T_6[9:0] ? ram_119 : _GEN_121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_123 = 10'h78 == _T_6[9:0] ? ram_120 : _GEN_122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_124 = 10'h79 == _T_6[9:0] ? ram_121 : _GEN_123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_125 = 10'h7a == _T_6[9:0] ? ram_122 : _GEN_124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_126 = 10'h7b == _T_6[9:0] ? ram_123 : _GEN_125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_127 = 10'h7c == _T_6[9:0] ? ram_124 : _GEN_126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_128 = 10'h7d == _T_6[9:0] ? ram_125 : _GEN_127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_129 = 10'h7e == _T_6[9:0] ? ram_126 : _GEN_128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_130 = 10'h7f == _T_6[9:0] ? ram_127 : _GEN_129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_131 = 10'h80 == _T_6[9:0] ? ram_128 : _GEN_130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_132 = 10'h81 == _T_6[9:0] ? ram_129 : _GEN_131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_133 = 10'h82 == _T_6[9:0] ? ram_130 : _GEN_132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_134 = 10'h83 == _T_6[9:0] ? ram_131 : _GEN_133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_135 = 10'h84 == _T_6[9:0] ? ram_132 : _GEN_134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_136 = 10'h85 == _T_6[9:0] ? ram_133 : _GEN_135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_137 = 10'h86 == _T_6[9:0] ? ram_134 : _GEN_136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_138 = 10'h87 == _T_6[9:0] ? ram_135 : _GEN_137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_139 = 10'h88 == _T_6[9:0] ? ram_136 : _GEN_138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_140 = 10'h89 == _T_6[9:0] ? ram_137 : _GEN_139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_141 = 10'h8a == _T_6[9:0] ? ram_138 : _GEN_140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_142 = 10'h8b == _T_6[9:0] ? ram_139 : _GEN_141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_143 = 10'h8c == _T_6[9:0] ? ram_140 : _GEN_142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_144 = 10'h8d == _T_6[9:0] ? ram_141 : _GEN_143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_145 = 10'h8e == _T_6[9:0] ? ram_142 : _GEN_144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_146 = 10'h8f == _T_6[9:0] ? ram_143 : _GEN_145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_147 = 10'h90 == _T_6[9:0] ? ram_144 : _GEN_146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_148 = 10'h91 == _T_6[9:0] ? ram_145 : _GEN_147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_149 = 10'h92 == _T_6[9:0] ? ram_146 : _GEN_148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_150 = 10'h93 == _T_6[9:0] ? ram_147 : _GEN_149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_151 = 10'h94 == _T_6[9:0] ? ram_148 : _GEN_150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_152 = 10'h95 == _T_6[9:0] ? ram_149 : _GEN_151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_153 = 10'h96 == _T_6[9:0] ? ram_150 : _GEN_152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_154 = 10'h97 == _T_6[9:0] ? ram_151 : _GEN_153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_155 = 10'h98 == _T_6[9:0] ? ram_152 : _GEN_154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_156 = 10'h99 == _T_6[9:0] ? ram_153 : _GEN_155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_157 = 10'h9a == _T_6[9:0] ? ram_154 : _GEN_156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_158 = 10'h9b == _T_6[9:0] ? ram_155 : _GEN_157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_159 = 10'h9c == _T_6[9:0] ? ram_156 : _GEN_158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_160 = 10'h9d == _T_6[9:0] ? ram_157 : _GEN_159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_161 = 10'h9e == _T_6[9:0] ? ram_158 : _GEN_160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_162 = 10'h9f == _T_6[9:0] ? ram_159 : _GEN_161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_163 = 10'ha0 == _T_6[9:0] ? ram_160 : _GEN_162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_164 = 10'ha1 == _T_6[9:0] ? ram_161 : _GEN_163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_165 = 10'ha2 == _T_6[9:0] ? ram_162 : _GEN_164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_166 = 10'ha3 == _T_6[9:0] ? ram_163 : _GEN_165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_167 = 10'ha4 == _T_6[9:0] ? ram_164 : _GEN_166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_168 = 10'ha5 == _T_6[9:0] ? ram_165 : _GEN_167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_169 = 10'ha6 == _T_6[9:0] ? ram_166 : _GEN_168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_170 = 10'ha7 == _T_6[9:0] ? ram_167 : _GEN_169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_171 = 10'ha8 == _T_6[9:0] ? ram_168 : _GEN_170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_172 = 10'ha9 == _T_6[9:0] ? ram_169 : _GEN_171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_173 = 10'haa == _T_6[9:0] ? ram_170 : _GEN_172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_174 = 10'hab == _T_6[9:0] ? ram_171 : _GEN_173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_175 = 10'hac == _T_6[9:0] ? ram_172 : _GEN_174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_176 = 10'had == _T_6[9:0] ? ram_173 : _GEN_175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_177 = 10'hae == _T_6[9:0] ? ram_174 : _GEN_176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_178 = 10'haf == _T_6[9:0] ? ram_175 : _GEN_177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_179 = 10'hb0 == _T_6[9:0] ? ram_176 : _GEN_178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_180 = 10'hb1 == _T_6[9:0] ? ram_177 : _GEN_179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_181 = 10'hb2 == _T_6[9:0] ? ram_178 : _GEN_180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_182 = 10'hb3 == _T_6[9:0] ? ram_179 : _GEN_181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_183 = 10'hb4 == _T_6[9:0] ? ram_180 : _GEN_182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_184 = 10'hb5 == _T_6[9:0] ? ram_181 : _GEN_183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_185 = 10'hb6 == _T_6[9:0] ? ram_182 : _GEN_184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_186 = 10'hb7 == _T_6[9:0] ? ram_183 : _GEN_185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_187 = 10'hb8 == _T_6[9:0] ? ram_184 : _GEN_186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_188 = 10'hb9 == _T_6[9:0] ? ram_185 : _GEN_187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_189 = 10'hba == _T_6[9:0] ? ram_186 : _GEN_188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_190 = 10'hbb == _T_6[9:0] ? ram_187 : _GEN_189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_191 = 10'hbc == _T_6[9:0] ? ram_188 : _GEN_190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_192 = 10'hbd == _T_6[9:0] ? ram_189 : _GEN_191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_193 = 10'hbe == _T_6[9:0] ? ram_190 : _GEN_192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_194 = 10'hbf == _T_6[9:0] ? ram_191 : _GEN_193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_195 = 10'hc0 == _T_6[9:0] ? ram_192 : _GEN_194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_196 = 10'hc1 == _T_6[9:0] ? ram_193 : _GEN_195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_197 = 10'hc2 == _T_6[9:0] ? ram_194 : _GEN_196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_198 = 10'hc3 == _T_6[9:0] ? ram_195 : _GEN_197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_199 = 10'hc4 == _T_6[9:0] ? ram_196 : _GEN_198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_200 = 10'hc5 == _T_6[9:0] ? ram_197 : _GEN_199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_201 = 10'hc6 == _T_6[9:0] ? ram_198 : _GEN_200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_202 = 10'hc7 == _T_6[9:0] ? ram_199 : _GEN_201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_203 = 10'hc8 == _T_6[9:0] ? ram_200 : _GEN_202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_204 = 10'hc9 == _T_6[9:0] ? ram_201 : _GEN_203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_205 = 10'hca == _T_6[9:0] ? ram_202 : _GEN_204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_206 = 10'hcb == _T_6[9:0] ? ram_203 : _GEN_205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_207 = 10'hcc == _T_6[9:0] ? ram_204 : _GEN_206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_208 = 10'hcd == _T_6[9:0] ? ram_205 : _GEN_207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_209 = 10'hce == _T_6[9:0] ? ram_206 : _GEN_208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_210 = 10'hcf == _T_6[9:0] ? ram_207 : _GEN_209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_211 = 10'hd0 == _T_6[9:0] ? ram_208 : _GEN_210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_212 = 10'hd1 == _T_6[9:0] ? ram_209 : _GEN_211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_213 = 10'hd2 == _T_6[9:0] ? ram_210 : _GEN_212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_214 = 10'hd3 == _T_6[9:0] ? ram_211 : _GEN_213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_215 = 10'hd4 == _T_6[9:0] ? ram_212 : _GEN_214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_216 = 10'hd5 == _T_6[9:0] ? ram_213 : _GEN_215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_217 = 10'hd6 == _T_6[9:0] ? ram_214 : _GEN_216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_218 = 10'hd7 == _T_6[9:0] ? ram_215 : _GEN_217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_219 = 10'hd8 == _T_6[9:0] ? ram_216 : _GEN_218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_220 = 10'hd9 == _T_6[9:0] ? ram_217 : _GEN_219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_221 = 10'hda == _T_6[9:0] ? ram_218 : _GEN_220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_222 = 10'hdb == _T_6[9:0] ? ram_219 : _GEN_221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_223 = 10'hdc == _T_6[9:0] ? ram_220 : _GEN_222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_224 = 10'hdd == _T_6[9:0] ? ram_221 : _GEN_223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_225 = 10'hde == _T_6[9:0] ? ram_222 : _GEN_224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_226 = 10'hdf == _T_6[9:0] ? ram_223 : _GEN_225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_227 = 10'he0 == _T_6[9:0] ? ram_224 : _GEN_226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_228 = 10'he1 == _T_6[9:0] ? ram_225 : _GEN_227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_229 = 10'he2 == _T_6[9:0] ? ram_226 : _GEN_228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_230 = 10'he3 == _T_6[9:0] ? ram_227 : _GEN_229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_231 = 10'he4 == _T_6[9:0] ? ram_228 : _GEN_230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_232 = 10'he5 == _T_6[9:0] ? ram_229 : _GEN_231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_233 = 10'he6 == _T_6[9:0] ? ram_230 : _GEN_232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_234 = 10'he7 == _T_6[9:0] ? ram_231 : _GEN_233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_235 = 10'he8 == _T_6[9:0] ? ram_232 : _GEN_234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_236 = 10'he9 == _T_6[9:0] ? ram_233 : _GEN_235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_237 = 10'hea == _T_6[9:0] ? ram_234 : _GEN_236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_238 = 10'heb == _T_6[9:0] ? ram_235 : _GEN_237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_239 = 10'hec == _T_6[9:0] ? ram_236 : _GEN_238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_240 = 10'hed == _T_6[9:0] ? ram_237 : _GEN_239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_241 = 10'hee == _T_6[9:0] ? ram_238 : _GEN_240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_242 = 10'hef == _T_6[9:0] ? ram_239 : _GEN_241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_243 = 10'hf0 == _T_6[9:0] ? ram_240 : _GEN_242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_244 = 10'hf1 == _T_6[9:0] ? ram_241 : _GEN_243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_245 = 10'hf2 == _T_6[9:0] ? ram_242 : _GEN_244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_246 = 10'hf3 == _T_6[9:0] ? ram_243 : _GEN_245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_247 = 10'hf4 == _T_6[9:0] ? ram_244 : _GEN_246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_248 = 10'hf5 == _T_6[9:0] ? ram_245 : _GEN_247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_249 = 10'hf6 == _T_6[9:0] ? ram_246 : _GEN_248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_250 = 10'hf7 == _T_6[9:0] ? ram_247 : _GEN_249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_251 = 10'hf8 == _T_6[9:0] ? ram_248 : _GEN_250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_252 = 10'hf9 == _T_6[9:0] ? ram_249 : _GEN_251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_253 = 10'hfa == _T_6[9:0] ? ram_250 : _GEN_252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_254 = 10'hfb == _T_6[9:0] ? ram_251 : _GEN_253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_255 = 10'hfc == _T_6[9:0] ? ram_252 : _GEN_254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_256 = 10'hfd == _T_6[9:0] ? ram_253 : _GEN_255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_257 = 10'hfe == _T_6[9:0] ? ram_254 : _GEN_256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_258 = 10'hff == _T_6[9:0] ? ram_255 : _GEN_257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_259 = 10'h100 == _T_6[9:0] ? ram_256 : _GEN_258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_260 = 10'h101 == _T_6[9:0] ? ram_257 : _GEN_259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_261 = 10'h102 == _T_6[9:0] ? ram_258 : _GEN_260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_262 = 10'h103 == _T_6[9:0] ? ram_259 : _GEN_261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_263 = 10'h104 == _T_6[9:0] ? ram_260 : _GEN_262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_264 = 10'h105 == _T_6[9:0] ? ram_261 : _GEN_263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_265 = 10'h106 == _T_6[9:0] ? ram_262 : _GEN_264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_266 = 10'h107 == _T_6[9:0] ? ram_263 : _GEN_265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_267 = 10'h108 == _T_6[9:0] ? ram_264 : _GEN_266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_268 = 10'h109 == _T_6[9:0] ? ram_265 : _GEN_267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_269 = 10'h10a == _T_6[9:0] ? ram_266 : _GEN_268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_270 = 10'h10b == _T_6[9:0] ? ram_267 : _GEN_269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_271 = 10'h10c == _T_6[9:0] ? ram_268 : _GEN_270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_272 = 10'h10d == _T_6[9:0] ? ram_269 : _GEN_271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_273 = 10'h10e == _T_6[9:0] ? ram_270 : _GEN_272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_274 = 10'h10f == _T_6[9:0] ? ram_271 : _GEN_273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_275 = 10'h110 == _T_6[9:0] ? ram_272 : _GEN_274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_276 = 10'h111 == _T_6[9:0] ? ram_273 : _GEN_275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_277 = 10'h112 == _T_6[9:0] ? ram_274 : _GEN_276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_278 = 10'h113 == _T_6[9:0] ? ram_275 : _GEN_277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_279 = 10'h114 == _T_6[9:0] ? ram_276 : _GEN_278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_280 = 10'h115 == _T_6[9:0] ? ram_277 : _GEN_279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_281 = 10'h116 == _T_6[9:0] ? ram_278 : _GEN_280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_282 = 10'h117 == _T_6[9:0] ? ram_279 : _GEN_281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_283 = 10'h118 == _T_6[9:0] ? ram_280 : _GEN_282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_284 = 10'h119 == _T_6[9:0] ? ram_281 : _GEN_283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_285 = 10'h11a == _T_6[9:0] ? ram_282 : _GEN_284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_286 = 10'h11b == _T_6[9:0] ? ram_283 : _GEN_285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_287 = 10'h11c == _T_6[9:0] ? ram_284 : _GEN_286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_288 = 10'h11d == _T_6[9:0] ? ram_285 : _GEN_287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_289 = 10'h11e == _T_6[9:0] ? ram_286 : _GEN_288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_290 = 10'h11f == _T_6[9:0] ? ram_287 : _GEN_289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_291 = 10'h120 == _T_6[9:0] ? ram_288 : _GEN_290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_292 = 10'h121 == _T_6[9:0] ? ram_289 : _GEN_291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_293 = 10'h122 == _T_6[9:0] ? ram_290 : _GEN_292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_294 = 10'h123 == _T_6[9:0] ? ram_291 : _GEN_293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_295 = 10'h124 == _T_6[9:0] ? ram_292 : _GEN_294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_296 = 10'h125 == _T_6[9:0] ? ram_293 : _GEN_295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_297 = 10'h126 == _T_6[9:0] ? ram_294 : _GEN_296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_298 = 10'h127 == _T_6[9:0] ? ram_295 : _GEN_297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_299 = 10'h128 == _T_6[9:0] ? ram_296 : _GEN_298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_300 = 10'h129 == _T_6[9:0] ? ram_297 : _GEN_299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_301 = 10'h12a == _T_6[9:0] ? ram_298 : _GEN_300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_302 = 10'h12b == _T_6[9:0] ? ram_299 : _GEN_301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_303 = 10'h12c == _T_6[9:0] ? ram_300 : _GEN_302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_304 = 10'h12d == _T_6[9:0] ? ram_301 : _GEN_303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_305 = 10'h12e == _T_6[9:0] ? ram_302 : _GEN_304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_306 = 10'h12f == _T_6[9:0] ? ram_303 : _GEN_305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_307 = 10'h130 == _T_6[9:0] ? ram_304 : _GEN_306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_308 = 10'h131 == _T_6[9:0] ? ram_305 : _GEN_307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_309 = 10'h132 == _T_6[9:0] ? ram_306 : _GEN_308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_310 = 10'h133 == _T_6[9:0] ? ram_307 : _GEN_309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_311 = 10'h134 == _T_6[9:0] ? ram_308 : _GEN_310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_312 = 10'h135 == _T_6[9:0] ? ram_309 : _GEN_311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_313 = 10'h136 == _T_6[9:0] ? ram_310 : _GEN_312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_314 = 10'h137 == _T_6[9:0] ? ram_311 : _GEN_313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_315 = 10'h138 == _T_6[9:0] ? ram_312 : _GEN_314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_316 = 10'h139 == _T_6[9:0] ? ram_313 : _GEN_315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_317 = 10'h13a == _T_6[9:0] ? ram_314 : _GEN_316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_318 = 10'h13b == _T_6[9:0] ? ram_315 : _GEN_317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_319 = 10'h13c == _T_6[9:0] ? ram_316 : _GEN_318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_320 = 10'h13d == _T_6[9:0] ? ram_317 : _GEN_319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_321 = 10'h13e == _T_6[9:0] ? ram_318 : _GEN_320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_322 = 10'h13f == _T_6[9:0] ? ram_319 : _GEN_321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_323 = 10'h140 == _T_6[9:0] ? ram_320 : _GEN_322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_324 = 10'h141 == _T_6[9:0] ? ram_321 : _GEN_323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_325 = 10'h142 == _T_6[9:0] ? ram_322 : _GEN_324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_326 = 10'h143 == _T_6[9:0] ? ram_323 : _GEN_325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_327 = 10'h144 == _T_6[9:0] ? ram_324 : _GEN_326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_328 = 10'h145 == _T_6[9:0] ? ram_325 : _GEN_327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_329 = 10'h146 == _T_6[9:0] ? ram_326 : _GEN_328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_330 = 10'h147 == _T_6[9:0] ? ram_327 : _GEN_329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_331 = 10'h148 == _T_6[9:0] ? ram_328 : _GEN_330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_332 = 10'h149 == _T_6[9:0] ? ram_329 : _GEN_331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_333 = 10'h14a == _T_6[9:0] ? ram_330 : _GEN_332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_334 = 10'h14b == _T_6[9:0] ? ram_331 : _GEN_333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_335 = 10'h14c == _T_6[9:0] ? ram_332 : _GEN_334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_336 = 10'h14d == _T_6[9:0] ? ram_333 : _GEN_335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_337 = 10'h14e == _T_6[9:0] ? ram_334 : _GEN_336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_338 = 10'h14f == _T_6[9:0] ? ram_335 : _GEN_337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_339 = 10'h150 == _T_6[9:0] ? ram_336 : _GEN_338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_340 = 10'h151 == _T_6[9:0] ? ram_337 : _GEN_339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_341 = 10'h152 == _T_6[9:0] ? ram_338 : _GEN_340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_342 = 10'h153 == _T_6[9:0] ? ram_339 : _GEN_341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_343 = 10'h154 == _T_6[9:0] ? ram_340 : _GEN_342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_344 = 10'h155 == _T_6[9:0] ? ram_341 : _GEN_343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_345 = 10'h156 == _T_6[9:0] ? ram_342 : _GEN_344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_346 = 10'h157 == _T_6[9:0] ? ram_343 : _GEN_345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_347 = 10'h158 == _T_6[9:0] ? ram_344 : _GEN_346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_348 = 10'h159 == _T_6[9:0] ? ram_345 : _GEN_347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_349 = 10'h15a == _T_6[9:0] ? ram_346 : _GEN_348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_350 = 10'h15b == _T_6[9:0] ? ram_347 : _GEN_349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_351 = 10'h15c == _T_6[9:0] ? ram_348 : _GEN_350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_352 = 10'h15d == _T_6[9:0] ? ram_349 : _GEN_351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_353 = 10'h15e == _T_6[9:0] ? ram_350 : _GEN_352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_354 = 10'h15f == _T_6[9:0] ? ram_351 : _GEN_353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_355 = 10'h160 == _T_6[9:0] ? ram_352 : _GEN_354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_356 = 10'h161 == _T_6[9:0] ? ram_353 : _GEN_355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_357 = 10'h162 == _T_6[9:0] ? ram_354 : _GEN_356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_358 = 10'h163 == _T_6[9:0] ? ram_355 : _GEN_357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_359 = 10'h164 == _T_6[9:0] ? ram_356 : _GEN_358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_360 = 10'h165 == _T_6[9:0] ? ram_357 : _GEN_359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_361 = 10'h166 == _T_6[9:0] ? ram_358 : _GEN_360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_362 = 10'h167 == _T_6[9:0] ? ram_359 : _GEN_361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_363 = 10'h168 == _T_6[9:0] ? ram_360 : _GEN_362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_364 = 10'h169 == _T_6[9:0] ? ram_361 : _GEN_363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_365 = 10'h16a == _T_6[9:0] ? ram_362 : _GEN_364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_366 = 10'h16b == _T_6[9:0] ? ram_363 : _GEN_365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_367 = 10'h16c == _T_6[9:0] ? ram_364 : _GEN_366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_368 = 10'h16d == _T_6[9:0] ? ram_365 : _GEN_367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_369 = 10'h16e == _T_6[9:0] ? ram_366 : _GEN_368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_370 = 10'h16f == _T_6[9:0] ? ram_367 : _GEN_369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_371 = 10'h170 == _T_6[9:0] ? ram_368 : _GEN_370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_372 = 10'h171 == _T_6[9:0] ? ram_369 : _GEN_371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_373 = 10'h172 == _T_6[9:0] ? ram_370 : _GEN_372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_374 = 10'h173 == _T_6[9:0] ? ram_371 : _GEN_373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_375 = 10'h174 == _T_6[9:0] ? ram_372 : _GEN_374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_376 = 10'h175 == _T_6[9:0] ? ram_373 : _GEN_375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_377 = 10'h176 == _T_6[9:0] ? ram_374 : _GEN_376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_378 = 10'h177 == _T_6[9:0] ? ram_375 : _GEN_377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_379 = 10'h178 == _T_6[9:0] ? ram_376 : _GEN_378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_380 = 10'h179 == _T_6[9:0] ? ram_377 : _GEN_379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_381 = 10'h17a == _T_6[9:0] ? ram_378 : _GEN_380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_382 = 10'h17b == _T_6[9:0] ? ram_379 : _GEN_381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_383 = 10'h17c == _T_6[9:0] ? ram_380 : _GEN_382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_384 = 10'h17d == _T_6[9:0] ? ram_381 : _GEN_383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_385 = 10'h17e == _T_6[9:0] ? ram_382 : _GEN_384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_386 = 10'h17f == _T_6[9:0] ? ram_383 : _GEN_385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_387 = 10'h180 == _T_6[9:0] ? ram_384 : _GEN_386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_388 = 10'h181 == _T_6[9:0] ? ram_385 : _GEN_387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_389 = 10'h182 == _T_6[9:0] ? ram_386 : _GEN_388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_390 = 10'h183 == _T_6[9:0] ? ram_387 : _GEN_389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_391 = 10'h184 == _T_6[9:0] ? ram_388 : _GEN_390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_392 = 10'h185 == _T_6[9:0] ? ram_389 : _GEN_391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_393 = 10'h186 == _T_6[9:0] ? ram_390 : _GEN_392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_394 = 10'h187 == _T_6[9:0] ? ram_391 : _GEN_393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_395 = 10'h188 == _T_6[9:0] ? ram_392 : _GEN_394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_396 = 10'h189 == _T_6[9:0] ? ram_393 : _GEN_395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_397 = 10'h18a == _T_6[9:0] ? ram_394 : _GEN_396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_398 = 10'h18b == _T_6[9:0] ? ram_395 : _GEN_397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_399 = 10'h18c == _T_6[9:0] ? ram_396 : _GEN_398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_400 = 10'h18d == _T_6[9:0] ? ram_397 : _GEN_399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_401 = 10'h18e == _T_6[9:0] ? ram_398 : _GEN_400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_402 = 10'h18f == _T_6[9:0] ? ram_399 : _GEN_401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_403 = 10'h190 == _T_6[9:0] ? ram_400 : _GEN_402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_404 = 10'h191 == _T_6[9:0] ? ram_401 : _GEN_403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_405 = 10'h192 == _T_6[9:0] ? ram_402 : _GEN_404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_406 = 10'h193 == _T_6[9:0] ? ram_403 : _GEN_405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_407 = 10'h194 == _T_6[9:0] ? ram_404 : _GEN_406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_408 = 10'h195 == _T_6[9:0] ? ram_405 : _GEN_407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_409 = 10'h196 == _T_6[9:0] ? ram_406 : _GEN_408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_410 = 10'h197 == _T_6[9:0] ? ram_407 : _GEN_409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_411 = 10'h198 == _T_6[9:0] ? ram_408 : _GEN_410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_412 = 10'h199 == _T_6[9:0] ? ram_409 : _GEN_411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_413 = 10'h19a == _T_6[9:0] ? ram_410 : _GEN_412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_414 = 10'h19b == _T_6[9:0] ? ram_411 : _GEN_413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_415 = 10'h19c == _T_6[9:0] ? ram_412 : _GEN_414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_416 = 10'h19d == _T_6[9:0] ? ram_413 : _GEN_415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_417 = 10'h19e == _T_6[9:0] ? ram_414 : _GEN_416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_418 = 10'h19f == _T_6[9:0] ? ram_415 : _GEN_417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_419 = 10'h1a0 == _T_6[9:0] ? ram_416 : _GEN_418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_420 = 10'h1a1 == _T_6[9:0] ? ram_417 : _GEN_419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_421 = 10'h1a2 == _T_6[9:0] ? ram_418 : _GEN_420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_422 = 10'h1a3 == _T_6[9:0] ? ram_419 : _GEN_421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_423 = 10'h1a4 == _T_6[9:0] ? ram_420 : _GEN_422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_424 = 10'h1a5 == _T_6[9:0] ? ram_421 : _GEN_423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_425 = 10'h1a6 == _T_6[9:0] ? ram_422 : _GEN_424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_426 = 10'h1a7 == _T_6[9:0] ? ram_423 : _GEN_425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_427 = 10'h1a8 == _T_6[9:0] ? ram_424 : _GEN_426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_428 = 10'h1a9 == _T_6[9:0] ? ram_425 : _GEN_427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_429 = 10'h1aa == _T_6[9:0] ? ram_426 : _GEN_428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_430 = 10'h1ab == _T_6[9:0] ? ram_427 : _GEN_429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_431 = 10'h1ac == _T_6[9:0] ? ram_428 : _GEN_430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_432 = 10'h1ad == _T_6[9:0] ? ram_429 : _GEN_431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_433 = 10'h1ae == _T_6[9:0] ? ram_430 : _GEN_432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_434 = 10'h1af == _T_6[9:0] ? ram_431 : _GEN_433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_435 = 10'h1b0 == _T_6[9:0] ? ram_432 : _GEN_434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_436 = 10'h1b1 == _T_6[9:0] ? ram_433 : _GEN_435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_437 = 10'h1b2 == _T_6[9:0] ? ram_434 : _GEN_436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_438 = 10'h1b3 == _T_6[9:0] ? ram_435 : _GEN_437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_439 = 10'h1b4 == _T_6[9:0] ? ram_436 : _GEN_438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_440 = 10'h1b5 == _T_6[9:0] ? ram_437 : _GEN_439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_441 = 10'h1b6 == _T_6[9:0] ? ram_438 : _GEN_440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_442 = 10'h1b7 == _T_6[9:0] ? ram_439 : _GEN_441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_443 = 10'h1b8 == _T_6[9:0] ? ram_440 : _GEN_442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_444 = 10'h1b9 == _T_6[9:0] ? ram_441 : _GEN_443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_445 = 10'h1ba == _T_6[9:0] ? ram_442 : _GEN_444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_446 = 10'h1bb == _T_6[9:0] ? ram_443 : _GEN_445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_447 = 10'h1bc == _T_6[9:0] ? ram_444 : _GEN_446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_448 = 10'h1bd == _T_6[9:0] ? ram_445 : _GEN_447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_449 = 10'h1be == _T_6[9:0] ? ram_446 : _GEN_448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_450 = 10'h1bf == _T_6[9:0] ? ram_447 : _GEN_449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_451 = 10'h1c0 == _T_6[9:0] ? ram_448 : _GEN_450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_452 = 10'h1c1 == _T_6[9:0] ? ram_449 : _GEN_451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_453 = 10'h1c2 == _T_6[9:0] ? ram_450 : _GEN_452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_454 = 10'h1c3 == _T_6[9:0] ? ram_451 : _GEN_453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_455 = 10'h1c4 == _T_6[9:0] ? ram_452 : _GEN_454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_456 = 10'h1c5 == _T_6[9:0] ? ram_453 : _GEN_455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_457 = 10'h1c6 == _T_6[9:0] ? ram_454 : _GEN_456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_458 = 10'h1c7 == _T_6[9:0] ? ram_455 : _GEN_457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_459 = 10'h1c8 == _T_6[9:0] ? ram_456 : _GEN_458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_460 = 10'h1c9 == _T_6[9:0] ? ram_457 : _GEN_459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_461 = 10'h1ca == _T_6[9:0] ? ram_458 : _GEN_460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_462 = 10'h1cb == _T_6[9:0] ? ram_459 : _GEN_461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_463 = 10'h1cc == _T_6[9:0] ? ram_460 : _GEN_462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_464 = 10'h1cd == _T_6[9:0] ? ram_461 : _GEN_463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_465 = 10'h1ce == _T_6[9:0] ? ram_462 : _GEN_464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_466 = 10'h1cf == _T_6[9:0] ? ram_463 : _GEN_465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_467 = 10'h1d0 == _T_6[9:0] ? ram_464 : _GEN_466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_468 = 10'h1d1 == _T_6[9:0] ? ram_465 : _GEN_467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_469 = 10'h1d2 == _T_6[9:0] ? ram_466 : _GEN_468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_470 = 10'h1d3 == _T_6[9:0] ? ram_467 : _GEN_469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_471 = 10'h1d4 == _T_6[9:0] ? ram_468 : _GEN_470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_472 = 10'h1d5 == _T_6[9:0] ? ram_469 : _GEN_471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_473 = 10'h1d6 == _T_6[9:0] ? ram_470 : _GEN_472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_474 = 10'h1d7 == _T_6[9:0] ? ram_471 : _GEN_473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_475 = 10'h1d8 == _T_6[9:0] ? ram_472 : _GEN_474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_476 = 10'h1d9 == _T_6[9:0] ? ram_473 : _GEN_475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_477 = 10'h1da == _T_6[9:0] ? ram_474 : _GEN_476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_478 = 10'h1db == _T_6[9:0] ? ram_475 : _GEN_477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_479 = 10'h1dc == _T_6[9:0] ? ram_476 : _GEN_478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_480 = 10'h1dd == _T_6[9:0] ? ram_477 : _GEN_479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_481 = 10'h1de == _T_6[9:0] ? ram_478 : _GEN_480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_482 = 10'h1df == _T_6[9:0] ? ram_479 : _GEN_481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_483 = 10'h1e0 == _T_6[9:0] ? ram_480 : _GEN_482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_484 = 10'h1e1 == _T_6[9:0] ? ram_481 : _GEN_483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_485 = 10'h1e2 == _T_6[9:0] ? ram_482 : _GEN_484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_486 = 10'h1e3 == _T_6[9:0] ? ram_483 : _GEN_485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_487 = 10'h1e4 == _T_6[9:0] ? ram_484 : _GEN_486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_488 = 10'h1e5 == _T_6[9:0] ? ram_485 : _GEN_487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_489 = 10'h1e6 == _T_6[9:0] ? ram_486 : _GEN_488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_490 = 10'h1e7 == _T_6[9:0] ? ram_487 : _GEN_489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_491 = 10'h1e8 == _T_6[9:0] ? ram_488 : _GEN_490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_492 = 10'h1e9 == _T_6[9:0] ? ram_489 : _GEN_491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_493 = 10'h1ea == _T_6[9:0] ? ram_490 : _GEN_492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_494 = 10'h1eb == _T_6[9:0] ? ram_491 : _GEN_493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_495 = 10'h1ec == _T_6[9:0] ? ram_492 : _GEN_494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_496 = 10'h1ed == _T_6[9:0] ? ram_493 : _GEN_495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_497 = 10'h1ee == _T_6[9:0] ? ram_494 : _GEN_496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_498 = 10'h1ef == _T_6[9:0] ? ram_495 : _GEN_497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_499 = 10'h1f0 == _T_6[9:0] ? ram_496 : _GEN_498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_500 = 10'h1f1 == _T_6[9:0] ? ram_497 : _GEN_499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_501 = 10'h1f2 == _T_6[9:0] ? ram_498 : _GEN_500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_502 = 10'h1f3 == _T_6[9:0] ? ram_499 : _GEN_501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_503 = 10'h1f4 == _T_6[9:0] ? ram_500 : _GEN_502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_504 = 10'h1f5 == _T_6[9:0] ? ram_501 : _GEN_503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_505 = 10'h1f6 == _T_6[9:0] ? ram_502 : _GEN_504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_506 = 10'h1f7 == _T_6[9:0] ? ram_503 : _GEN_505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_507 = 10'h1f8 == _T_6[9:0] ? ram_504 : _GEN_506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_508 = 10'h1f9 == _T_6[9:0] ? ram_505 : _GEN_507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_509 = 10'h1fa == _T_6[9:0] ? ram_506 : _GEN_508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_510 = 10'h1fb == _T_6[9:0] ? ram_507 : _GEN_509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_511 = 10'h1fc == _T_6[9:0] ? ram_508 : _GEN_510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_512 = 10'h1fd == _T_6[9:0] ? ram_509 : _GEN_511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_513 = 10'h1fe == _T_6[9:0] ? ram_510 : _GEN_512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_514 = 10'h1ff == _T_6[9:0] ? ram_511 : _GEN_513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_515 = 10'h200 == _T_6[9:0] ? ram_512 : _GEN_514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_516 = 10'h201 == _T_6[9:0] ? ram_513 : _GEN_515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_517 = 10'h202 == _T_6[9:0] ? ram_514 : _GEN_516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_518 = 10'h203 == _T_6[9:0] ? ram_515 : _GEN_517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_519 = 10'h204 == _T_6[9:0] ? ram_516 : _GEN_518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_520 = 10'h205 == _T_6[9:0] ? ram_517 : _GEN_519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_521 = 10'h206 == _T_6[9:0] ? ram_518 : _GEN_520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_522 = 10'h207 == _T_6[9:0] ? ram_519 : _GEN_521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_523 = 10'h208 == _T_6[9:0] ? ram_520 : _GEN_522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_524 = 10'h209 == _T_6[9:0] ? ram_521 : _GEN_523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_525 = 10'h20a == _T_6[9:0] ? ram_522 : _GEN_524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_526 = 10'h20b == _T_6[9:0] ? ram_523 : _GEN_525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_527 = 10'h20c == _T_6[9:0] ? ram_524 : _GEN_526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19061 = {{8190'd0}, _GEN_527}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_25 = _GEN_19061 ^ _ram_T_24; // @[vga.scala 64:41]
  wire [287:0] _GEN_528 = 10'h0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_0; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_529 = 10'h1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_1; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_530 = 10'h2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_2; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_531 = 10'h3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_3; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_532 = 10'h4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_4; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_533 = 10'h5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_5; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_534 = 10'h6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_6; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_535 = 10'h7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_7; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_536 = 10'h8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_8; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_537 = 10'h9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_9; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_538 = 10'ha == _T_6[9:0] ? _ram_T_25[287:0] : ram_10; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_539 = 10'hb == _T_6[9:0] ? _ram_T_25[287:0] : ram_11; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_540 = 10'hc == _T_6[9:0] ? _ram_T_25[287:0] : ram_12; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_541 = 10'hd == _T_6[9:0] ? _ram_T_25[287:0] : ram_13; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_542 = 10'he == _T_6[9:0] ? _ram_T_25[287:0] : ram_14; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_543 = 10'hf == _T_6[9:0] ? _ram_T_25[287:0] : ram_15; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_544 = 10'h10 == _T_6[9:0] ? _ram_T_25[287:0] : ram_16; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_545 = 10'h11 == _T_6[9:0] ? _ram_T_25[287:0] : ram_17; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_546 = 10'h12 == _T_6[9:0] ? _ram_T_25[287:0] : ram_18; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_547 = 10'h13 == _T_6[9:0] ? _ram_T_25[287:0] : ram_19; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_548 = 10'h14 == _T_6[9:0] ? _ram_T_25[287:0] : ram_20; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_549 = 10'h15 == _T_6[9:0] ? _ram_T_25[287:0] : ram_21; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_550 = 10'h16 == _T_6[9:0] ? _ram_T_25[287:0] : ram_22; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_551 = 10'h17 == _T_6[9:0] ? _ram_T_25[287:0] : ram_23; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_552 = 10'h18 == _T_6[9:0] ? _ram_T_25[287:0] : ram_24; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_553 = 10'h19 == _T_6[9:0] ? _ram_T_25[287:0] : ram_25; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_554 = 10'h1a == _T_6[9:0] ? _ram_T_25[287:0] : ram_26; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_555 = 10'h1b == _T_6[9:0] ? _ram_T_25[287:0] : ram_27; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_556 = 10'h1c == _T_6[9:0] ? _ram_T_25[287:0] : ram_28; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_557 = 10'h1d == _T_6[9:0] ? _ram_T_25[287:0] : ram_29; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_558 = 10'h1e == _T_6[9:0] ? _ram_T_25[287:0] : ram_30; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_559 = 10'h1f == _T_6[9:0] ? _ram_T_25[287:0] : ram_31; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_560 = 10'h20 == _T_6[9:0] ? _ram_T_25[287:0] : ram_32; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_561 = 10'h21 == _T_6[9:0] ? _ram_T_25[287:0] : ram_33; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_562 = 10'h22 == _T_6[9:0] ? _ram_T_25[287:0] : ram_34; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_563 = 10'h23 == _T_6[9:0] ? _ram_T_25[287:0] : ram_35; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_564 = 10'h24 == _T_6[9:0] ? _ram_T_25[287:0] : ram_36; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_565 = 10'h25 == _T_6[9:0] ? _ram_T_25[287:0] : ram_37; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_566 = 10'h26 == _T_6[9:0] ? _ram_T_25[287:0] : ram_38; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_567 = 10'h27 == _T_6[9:0] ? _ram_T_25[287:0] : ram_39; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_568 = 10'h28 == _T_6[9:0] ? _ram_T_25[287:0] : ram_40; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_569 = 10'h29 == _T_6[9:0] ? _ram_T_25[287:0] : ram_41; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_570 = 10'h2a == _T_6[9:0] ? _ram_T_25[287:0] : ram_42; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_571 = 10'h2b == _T_6[9:0] ? _ram_T_25[287:0] : ram_43; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_572 = 10'h2c == _T_6[9:0] ? _ram_T_25[287:0] : ram_44; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_573 = 10'h2d == _T_6[9:0] ? _ram_T_25[287:0] : ram_45; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_574 = 10'h2e == _T_6[9:0] ? _ram_T_25[287:0] : ram_46; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_575 = 10'h2f == _T_6[9:0] ? _ram_T_25[287:0] : ram_47; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_576 = 10'h30 == _T_6[9:0] ? _ram_T_25[287:0] : ram_48; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_577 = 10'h31 == _T_6[9:0] ? _ram_T_25[287:0] : ram_49; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_578 = 10'h32 == _T_6[9:0] ? _ram_T_25[287:0] : ram_50; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_579 = 10'h33 == _T_6[9:0] ? _ram_T_25[287:0] : ram_51; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_580 = 10'h34 == _T_6[9:0] ? _ram_T_25[287:0] : ram_52; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_581 = 10'h35 == _T_6[9:0] ? _ram_T_25[287:0] : ram_53; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_582 = 10'h36 == _T_6[9:0] ? _ram_T_25[287:0] : ram_54; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_583 = 10'h37 == _T_6[9:0] ? _ram_T_25[287:0] : ram_55; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_584 = 10'h38 == _T_6[9:0] ? _ram_T_25[287:0] : ram_56; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_585 = 10'h39 == _T_6[9:0] ? _ram_T_25[287:0] : ram_57; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_586 = 10'h3a == _T_6[9:0] ? _ram_T_25[287:0] : ram_58; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_587 = 10'h3b == _T_6[9:0] ? _ram_T_25[287:0] : ram_59; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_588 = 10'h3c == _T_6[9:0] ? _ram_T_25[287:0] : ram_60; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_589 = 10'h3d == _T_6[9:0] ? _ram_T_25[287:0] : ram_61; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_590 = 10'h3e == _T_6[9:0] ? _ram_T_25[287:0] : ram_62; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_591 = 10'h3f == _T_6[9:0] ? _ram_T_25[287:0] : ram_63; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_592 = 10'h40 == _T_6[9:0] ? _ram_T_25[287:0] : ram_64; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_593 = 10'h41 == _T_6[9:0] ? _ram_T_25[287:0] : ram_65; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_594 = 10'h42 == _T_6[9:0] ? _ram_T_25[287:0] : ram_66; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_595 = 10'h43 == _T_6[9:0] ? _ram_T_25[287:0] : ram_67; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_596 = 10'h44 == _T_6[9:0] ? _ram_T_25[287:0] : ram_68; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_597 = 10'h45 == _T_6[9:0] ? _ram_T_25[287:0] : ram_69; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_598 = 10'h46 == _T_6[9:0] ? _ram_T_25[287:0] : ram_70; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_599 = 10'h47 == _T_6[9:0] ? _ram_T_25[287:0] : ram_71; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_600 = 10'h48 == _T_6[9:0] ? _ram_T_25[287:0] : ram_72; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_601 = 10'h49 == _T_6[9:0] ? _ram_T_25[287:0] : ram_73; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_602 = 10'h4a == _T_6[9:0] ? _ram_T_25[287:0] : ram_74; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_603 = 10'h4b == _T_6[9:0] ? _ram_T_25[287:0] : ram_75; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_604 = 10'h4c == _T_6[9:0] ? _ram_T_25[287:0] : ram_76; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_605 = 10'h4d == _T_6[9:0] ? _ram_T_25[287:0] : ram_77; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_606 = 10'h4e == _T_6[9:0] ? _ram_T_25[287:0] : ram_78; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_607 = 10'h4f == _T_6[9:0] ? _ram_T_25[287:0] : ram_79; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_608 = 10'h50 == _T_6[9:0] ? _ram_T_25[287:0] : ram_80; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_609 = 10'h51 == _T_6[9:0] ? _ram_T_25[287:0] : ram_81; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_610 = 10'h52 == _T_6[9:0] ? _ram_T_25[287:0] : ram_82; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_611 = 10'h53 == _T_6[9:0] ? _ram_T_25[287:0] : ram_83; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_612 = 10'h54 == _T_6[9:0] ? _ram_T_25[287:0] : ram_84; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_613 = 10'h55 == _T_6[9:0] ? _ram_T_25[287:0] : ram_85; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_614 = 10'h56 == _T_6[9:0] ? _ram_T_25[287:0] : ram_86; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_615 = 10'h57 == _T_6[9:0] ? _ram_T_25[287:0] : ram_87; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_616 = 10'h58 == _T_6[9:0] ? _ram_T_25[287:0] : ram_88; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_617 = 10'h59 == _T_6[9:0] ? _ram_T_25[287:0] : ram_89; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_618 = 10'h5a == _T_6[9:0] ? _ram_T_25[287:0] : ram_90; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_619 = 10'h5b == _T_6[9:0] ? _ram_T_25[287:0] : ram_91; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_620 = 10'h5c == _T_6[9:0] ? _ram_T_25[287:0] : ram_92; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_621 = 10'h5d == _T_6[9:0] ? _ram_T_25[287:0] : ram_93; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_622 = 10'h5e == _T_6[9:0] ? _ram_T_25[287:0] : ram_94; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_623 = 10'h5f == _T_6[9:0] ? _ram_T_25[287:0] : ram_95; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_624 = 10'h60 == _T_6[9:0] ? _ram_T_25[287:0] : ram_96; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_625 = 10'h61 == _T_6[9:0] ? _ram_T_25[287:0] : ram_97; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_626 = 10'h62 == _T_6[9:0] ? _ram_T_25[287:0] : ram_98; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_627 = 10'h63 == _T_6[9:0] ? _ram_T_25[287:0] : ram_99; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_628 = 10'h64 == _T_6[9:0] ? _ram_T_25[287:0] : ram_100; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_629 = 10'h65 == _T_6[9:0] ? _ram_T_25[287:0] : ram_101; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_630 = 10'h66 == _T_6[9:0] ? _ram_T_25[287:0] : ram_102; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_631 = 10'h67 == _T_6[9:0] ? _ram_T_25[287:0] : ram_103; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_632 = 10'h68 == _T_6[9:0] ? _ram_T_25[287:0] : ram_104; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_633 = 10'h69 == _T_6[9:0] ? _ram_T_25[287:0] : ram_105; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_634 = 10'h6a == _T_6[9:0] ? _ram_T_25[287:0] : ram_106; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_635 = 10'h6b == _T_6[9:0] ? _ram_T_25[287:0] : ram_107; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_636 = 10'h6c == _T_6[9:0] ? _ram_T_25[287:0] : ram_108; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_637 = 10'h6d == _T_6[9:0] ? _ram_T_25[287:0] : ram_109; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_638 = 10'h6e == _T_6[9:0] ? _ram_T_25[287:0] : ram_110; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_639 = 10'h6f == _T_6[9:0] ? _ram_T_25[287:0] : ram_111; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_640 = 10'h70 == _T_6[9:0] ? _ram_T_25[287:0] : ram_112; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_641 = 10'h71 == _T_6[9:0] ? _ram_T_25[287:0] : ram_113; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_642 = 10'h72 == _T_6[9:0] ? _ram_T_25[287:0] : ram_114; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_643 = 10'h73 == _T_6[9:0] ? _ram_T_25[287:0] : ram_115; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_644 = 10'h74 == _T_6[9:0] ? _ram_T_25[287:0] : ram_116; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_645 = 10'h75 == _T_6[9:0] ? _ram_T_25[287:0] : ram_117; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_646 = 10'h76 == _T_6[9:0] ? _ram_T_25[287:0] : ram_118; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_647 = 10'h77 == _T_6[9:0] ? _ram_T_25[287:0] : ram_119; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_648 = 10'h78 == _T_6[9:0] ? _ram_T_25[287:0] : ram_120; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_649 = 10'h79 == _T_6[9:0] ? _ram_T_25[287:0] : ram_121; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_650 = 10'h7a == _T_6[9:0] ? _ram_T_25[287:0] : ram_122; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_651 = 10'h7b == _T_6[9:0] ? _ram_T_25[287:0] : ram_123; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_652 = 10'h7c == _T_6[9:0] ? _ram_T_25[287:0] : ram_124; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_653 = 10'h7d == _T_6[9:0] ? _ram_T_25[287:0] : ram_125; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_654 = 10'h7e == _T_6[9:0] ? _ram_T_25[287:0] : ram_126; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_655 = 10'h7f == _T_6[9:0] ? _ram_T_25[287:0] : ram_127; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_656 = 10'h80 == _T_6[9:0] ? _ram_T_25[287:0] : ram_128; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_657 = 10'h81 == _T_6[9:0] ? _ram_T_25[287:0] : ram_129; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_658 = 10'h82 == _T_6[9:0] ? _ram_T_25[287:0] : ram_130; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_659 = 10'h83 == _T_6[9:0] ? _ram_T_25[287:0] : ram_131; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_660 = 10'h84 == _T_6[9:0] ? _ram_T_25[287:0] : ram_132; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_661 = 10'h85 == _T_6[9:0] ? _ram_T_25[287:0] : ram_133; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_662 = 10'h86 == _T_6[9:0] ? _ram_T_25[287:0] : ram_134; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_663 = 10'h87 == _T_6[9:0] ? _ram_T_25[287:0] : ram_135; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_664 = 10'h88 == _T_6[9:0] ? _ram_T_25[287:0] : ram_136; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_665 = 10'h89 == _T_6[9:0] ? _ram_T_25[287:0] : ram_137; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_666 = 10'h8a == _T_6[9:0] ? _ram_T_25[287:0] : ram_138; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_667 = 10'h8b == _T_6[9:0] ? _ram_T_25[287:0] : ram_139; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_668 = 10'h8c == _T_6[9:0] ? _ram_T_25[287:0] : ram_140; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_669 = 10'h8d == _T_6[9:0] ? _ram_T_25[287:0] : ram_141; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_670 = 10'h8e == _T_6[9:0] ? _ram_T_25[287:0] : ram_142; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_671 = 10'h8f == _T_6[9:0] ? _ram_T_25[287:0] : ram_143; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_672 = 10'h90 == _T_6[9:0] ? _ram_T_25[287:0] : ram_144; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_673 = 10'h91 == _T_6[9:0] ? _ram_T_25[287:0] : ram_145; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_674 = 10'h92 == _T_6[9:0] ? _ram_T_25[287:0] : ram_146; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_675 = 10'h93 == _T_6[9:0] ? _ram_T_25[287:0] : ram_147; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_676 = 10'h94 == _T_6[9:0] ? _ram_T_25[287:0] : ram_148; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_677 = 10'h95 == _T_6[9:0] ? _ram_T_25[287:0] : ram_149; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_678 = 10'h96 == _T_6[9:0] ? _ram_T_25[287:0] : ram_150; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_679 = 10'h97 == _T_6[9:0] ? _ram_T_25[287:0] : ram_151; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_680 = 10'h98 == _T_6[9:0] ? _ram_T_25[287:0] : ram_152; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_681 = 10'h99 == _T_6[9:0] ? _ram_T_25[287:0] : ram_153; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_682 = 10'h9a == _T_6[9:0] ? _ram_T_25[287:0] : ram_154; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_683 = 10'h9b == _T_6[9:0] ? _ram_T_25[287:0] : ram_155; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_684 = 10'h9c == _T_6[9:0] ? _ram_T_25[287:0] : ram_156; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_685 = 10'h9d == _T_6[9:0] ? _ram_T_25[287:0] : ram_157; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_686 = 10'h9e == _T_6[9:0] ? _ram_T_25[287:0] : ram_158; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_687 = 10'h9f == _T_6[9:0] ? _ram_T_25[287:0] : ram_159; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_688 = 10'ha0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_160; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_689 = 10'ha1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_161; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_690 = 10'ha2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_162; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_691 = 10'ha3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_163; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_692 = 10'ha4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_164; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_693 = 10'ha5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_165; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_694 = 10'ha6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_166; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_695 = 10'ha7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_167; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_696 = 10'ha8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_168; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_697 = 10'ha9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_169; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_698 = 10'haa == _T_6[9:0] ? _ram_T_25[287:0] : ram_170; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_699 = 10'hab == _T_6[9:0] ? _ram_T_25[287:0] : ram_171; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_700 = 10'hac == _T_6[9:0] ? _ram_T_25[287:0] : ram_172; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_701 = 10'had == _T_6[9:0] ? _ram_T_25[287:0] : ram_173; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_702 = 10'hae == _T_6[9:0] ? _ram_T_25[287:0] : ram_174; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_703 = 10'haf == _T_6[9:0] ? _ram_T_25[287:0] : ram_175; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_704 = 10'hb0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_176; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_705 = 10'hb1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_177; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_706 = 10'hb2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_178; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_707 = 10'hb3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_179; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_708 = 10'hb4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_180; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_709 = 10'hb5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_181; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_710 = 10'hb6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_182; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_711 = 10'hb7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_183; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_712 = 10'hb8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_184; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_713 = 10'hb9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_185; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_714 = 10'hba == _T_6[9:0] ? _ram_T_25[287:0] : ram_186; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_715 = 10'hbb == _T_6[9:0] ? _ram_T_25[287:0] : ram_187; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_716 = 10'hbc == _T_6[9:0] ? _ram_T_25[287:0] : ram_188; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_717 = 10'hbd == _T_6[9:0] ? _ram_T_25[287:0] : ram_189; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_718 = 10'hbe == _T_6[9:0] ? _ram_T_25[287:0] : ram_190; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_719 = 10'hbf == _T_6[9:0] ? _ram_T_25[287:0] : ram_191; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_720 = 10'hc0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_192; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_721 = 10'hc1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_193; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_722 = 10'hc2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_194; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_723 = 10'hc3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_195; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_724 = 10'hc4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_196; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_725 = 10'hc5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_197; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_726 = 10'hc6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_198; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_727 = 10'hc7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_199; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_728 = 10'hc8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_200; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_729 = 10'hc9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_201; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_730 = 10'hca == _T_6[9:0] ? _ram_T_25[287:0] : ram_202; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_731 = 10'hcb == _T_6[9:0] ? _ram_T_25[287:0] : ram_203; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_732 = 10'hcc == _T_6[9:0] ? _ram_T_25[287:0] : ram_204; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_733 = 10'hcd == _T_6[9:0] ? _ram_T_25[287:0] : ram_205; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_734 = 10'hce == _T_6[9:0] ? _ram_T_25[287:0] : ram_206; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_735 = 10'hcf == _T_6[9:0] ? _ram_T_25[287:0] : ram_207; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_736 = 10'hd0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_208; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_737 = 10'hd1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_209; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_738 = 10'hd2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_210; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_739 = 10'hd3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_211; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_740 = 10'hd4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_212; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_741 = 10'hd5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_213; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_742 = 10'hd6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_214; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_743 = 10'hd7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_215; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_744 = 10'hd8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_216; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_745 = 10'hd9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_217; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_746 = 10'hda == _T_6[9:0] ? _ram_T_25[287:0] : ram_218; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_747 = 10'hdb == _T_6[9:0] ? _ram_T_25[287:0] : ram_219; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_748 = 10'hdc == _T_6[9:0] ? _ram_T_25[287:0] : ram_220; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_749 = 10'hdd == _T_6[9:0] ? _ram_T_25[287:0] : ram_221; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_750 = 10'hde == _T_6[9:0] ? _ram_T_25[287:0] : ram_222; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_751 = 10'hdf == _T_6[9:0] ? _ram_T_25[287:0] : ram_223; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_752 = 10'he0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_224; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_753 = 10'he1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_225; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_754 = 10'he2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_226; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_755 = 10'he3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_227; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_756 = 10'he4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_228; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_757 = 10'he5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_229; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_758 = 10'he6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_230; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_759 = 10'he7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_231; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_760 = 10'he8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_232; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_761 = 10'he9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_233; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_762 = 10'hea == _T_6[9:0] ? _ram_T_25[287:0] : ram_234; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_763 = 10'heb == _T_6[9:0] ? _ram_T_25[287:0] : ram_235; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_764 = 10'hec == _T_6[9:0] ? _ram_T_25[287:0] : ram_236; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_765 = 10'hed == _T_6[9:0] ? _ram_T_25[287:0] : ram_237; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_766 = 10'hee == _T_6[9:0] ? _ram_T_25[287:0] : ram_238; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_767 = 10'hef == _T_6[9:0] ? _ram_T_25[287:0] : ram_239; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_768 = 10'hf0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_240; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_769 = 10'hf1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_241; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_770 = 10'hf2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_242; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_771 = 10'hf3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_243; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_772 = 10'hf4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_244; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_773 = 10'hf5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_245; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_774 = 10'hf6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_246; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_775 = 10'hf7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_247; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_776 = 10'hf8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_248; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_777 = 10'hf9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_249; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_778 = 10'hfa == _T_6[9:0] ? _ram_T_25[287:0] : ram_250; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_779 = 10'hfb == _T_6[9:0] ? _ram_T_25[287:0] : ram_251; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_780 = 10'hfc == _T_6[9:0] ? _ram_T_25[287:0] : ram_252; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_781 = 10'hfd == _T_6[9:0] ? _ram_T_25[287:0] : ram_253; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_782 = 10'hfe == _T_6[9:0] ? _ram_T_25[287:0] : ram_254; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_783 = 10'hff == _T_6[9:0] ? _ram_T_25[287:0] : ram_255; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_784 = 10'h100 == _T_6[9:0] ? _ram_T_25[287:0] : ram_256; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_785 = 10'h101 == _T_6[9:0] ? _ram_T_25[287:0] : ram_257; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_786 = 10'h102 == _T_6[9:0] ? _ram_T_25[287:0] : ram_258; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_787 = 10'h103 == _T_6[9:0] ? _ram_T_25[287:0] : ram_259; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_788 = 10'h104 == _T_6[9:0] ? _ram_T_25[287:0] : ram_260; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_789 = 10'h105 == _T_6[9:0] ? _ram_T_25[287:0] : ram_261; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_790 = 10'h106 == _T_6[9:0] ? _ram_T_25[287:0] : ram_262; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_791 = 10'h107 == _T_6[9:0] ? _ram_T_25[287:0] : ram_263; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_792 = 10'h108 == _T_6[9:0] ? _ram_T_25[287:0] : ram_264; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_793 = 10'h109 == _T_6[9:0] ? _ram_T_25[287:0] : ram_265; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_794 = 10'h10a == _T_6[9:0] ? _ram_T_25[287:0] : ram_266; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_795 = 10'h10b == _T_6[9:0] ? _ram_T_25[287:0] : ram_267; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_796 = 10'h10c == _T_6[9:0] ? _ram_T_25[287:0] : ram_268; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_797 = 10'h10d == _T_6[9:0] ? _ram_T_25[287:0] : ram_269; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_798 = 10'h10e == _T_6[9:0] ? _ram_T_25[287:0] : ram_270; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_799 = 10'h10f == _T_6[9:0] ? _ram_T_25[287:0] : ram_271; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_800 = 10'h110 == _T_6[9:0] ? _ram_T_25[287:0] : ram_272; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_801 = 10'h111 == _T_6[9:0] ? _ram_T_25[287:0] : ram_273; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_802 = 10'h112 == _T_6[9:0] ? _ram_T_25[287:0] : ram_274; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_803 = 10'h113 == _T_6[9:0] ? _ram_T_25[287:0] : ram_275; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_804 = 10'h114 == _T_6[9:0] ? _ram_T_25[287:0] : ram_276; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_805 = 10'h115 == _T_6[9:0] ? _ram_T_25[287:0] : ram_277; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_806 = 10'h116 == _T_6[9:0] ? _ram_T_25[287:0] : ram_278; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_807 = 10'h117 == _T_6[9:0] ? _ram_T_25[287:0] : ram_279; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_808 = 10'h118 == _T_6[9:0] ? _ram_T_25[287:0] : ram_280; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_809 = 10'h119 == _T_6[9:0] ? _ram_T_25[287:0] : ram_281; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_810 = 10'h11a == _T_6[9:0] ? _ram_T_25[287:0] : ram_282; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_811 = 10'h11b == _T_6[9:0] ? _ram_T_25[287:0] : ram_283; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_812 = 10'h11c == _T_6[9:0] ? _ram_T_25[287:0] : ram_284; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_813 = 10'h11d == _T_6[9:0] ? _ram_T_25[287:0] : ram_285; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_814 = 10'h11e == _T_6[9:0] ? _ram_T_25[287:0] : ram_286; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_815 = 10'h11f == _T_6[9:0] ? _ram_T_25[287:0] : ram_287; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_816 = 10'h120 == _T_6[9:0] ? _ram_T_25[287:0] : ram_288; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_817 = 10'h121 == _T_6[9:0] ? _ram_T_25[287:0] : ram_289; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_818 = 10'h122 == _T_6[9:0] ? _ram_T_25[287:0] : ram_290; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_819 = 10'h123 == _T_6[9:0] ? _ram_T_25[287:0] : ram_291; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_820 = 10'h124 == _T_6[9:0] ? _ram_T_25[287:0] : ram_292; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_821 = 10'h125 == _T_6[9:0] ? _ram_T_25[287:0] : ram_293; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_822 = 10'h126 == _T_6[9:0] ? _ram_T_25[287:0] : ram_294; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_823 = 10'h127 == _T_6[9:0] ? _ram_T_25[287:0] : ram_295; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_824 = 10'h128 == _T_6[9:0] ? _ram_T_25[287:0] : ram_296; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_825 = 10'h129 == _T_6[9:0] ? _ram_T_25[287:0] : ram_297; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_826 = 10'h12a == _T_6[9:0] ? _ram_T_25[287:0] : ram_298; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_827 = 10'h12b == _T_6[9:0] ? _ram_T_25[287:0] : ram_299; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_828 = 10'h12c == _T_6[9:0] ? _ram_T_25[287:0] : ram_300; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_829 = 10'h12d == _T_6[9:0] ? _ram_T_25[287:0] : ram_301; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_830 = 10'h12e == _T_6[9:0] ? _ram_T_25[287:0] : ram_302; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_831 = 10'h12f == _T_6[9:0] ? _ram_T_25[287:0] : ram_303; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_832 = 10'h130 == _T_6[9:0] ? _ram_T_25[287:0] : ram_304; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_833 = 10'h131 == _T_6[9:0] ? _ram_T_25[287:0] : ram_305; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_834 = 10'h132 == _T_6[9:0] ? _ram_T_25[287:0] : ram_306; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_835 = 10'h133 == _T_6[9:0] ? _ram_T_25[287:0] : ram_307; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_836 = 10'h134 == _T_6[9:0] ? _ram_T_25[287:0] : ram_308; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_837 = 10'h135 == _T_6[9:0] ? _ram_T_25[287:0] : ram_309; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_838 = 10'h136 == _T_6[9:0] ? _ram_T_25[287:0] : ram_310; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_839 = 10'h137 == _T_6[9:0] ? _ram_T_25[287:0] : ram_311; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_840 = 10'h138 == _T_6[9:0] ? _ram_T_25[287:0] : ram_312; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_841 = 10'h139 == _T_6[9:0] ? _ram_T_25[287:0] : ram_313; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_842 = 10'h13a == _T_6[9:0] ? _ram_T_25[287:0] : ram_314; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_843 = 10'h13b == _T_6[9:0] ? _ram_T_25[287:0] : ram_315; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_844 = 10'h13c == _T_6[9:0] ? _ram_T_25[287:0] : ram_316; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_845 = 10'h13d == _T_6[9:0] ? _ram_T_25[287:0] : ram_317; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_846 = 10'h13e == _T_6[9:0] ? _ram_T_25[287:0] : ram_318; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_847 = 10'h13f == _T_6[9:0] ? _ram_T_25[287:0] : ram_319; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_848 = 10'h140 == _T_6[9:0] ? _ram_T_25[287:0] : ram_320; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_849 = 10'h141 == _T_6[9:0] ? _ram_T_25[287:0] : ram_321; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_850 = 10'h142 == _T_6[9:0] ? _ram_T_25[287:0] : ram_322; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_851 = 10'h143 == _T_6[9:0] ? _ram_T_25[287:0] : ram_323; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_852 = 10'h144 == _T_6[9:0] ? _ram_T_25[287:0] : ram_324; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_853 = 10'h145 == _T_6[9:0] ? _ram_T_25[287:0] : ram_325; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_854 = 10'h146 == _T_6[9:0] ? _ram_T_25[287:0] : ram_326; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_855 = 10'h147 == _T_6[9:0] ? _ram_T_25[287:0] : ram_327; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_856 = 10'h148 == _T_6[9:0] ? _ram_T_25[287:0] : ram_328; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_857 = 10'h149 == _T_6[9:0] ? _ram_T_25[287:0] : ram_329; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_858 = 10'h14a == _T_6[9:0] ? _ram_T_25[287:0] : ram_330; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_859 = 10'h14b == _T_6[9:0] ? _ram_T_25[287:0] : ram_331; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_860 = 10'h14c == _T_6[9:0] ? _ram_T_25[287:0] : ram_332; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_861 = 10'h14d == _T_6[9:0] ? _ram_T_25[287:0] : ram_333; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_862 = 10'h14e == _T_6[9:0] ? _ram_T_25[287:0] : ram_334; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_863 = 10'h14f == _T_6[9:0] ? _ram_T_25[287:0] : ram_335; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_864 = 10'h150 == _T_6[9:0] ? _ram_T_25[287:0] : ram_336; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_865 = 10'h151 == _T_6[9:0] ? _ram_T_25[287:0] : ram_337; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_866 = 10'h152 == _T_6[9:0] ? _ram_T_25[287:0] : ram_338; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_867 = 10'h153 == _T_6[9:0] ? _ram_T_25[287:0] : ram_339; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_868 = 10'h154 == _T_6[9:0] ? _ram_T_25[287:0] : ram_340; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_869 = 10'h155 == _T_6[9:0] ? _ram_T_25[287:0] : ram_341; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_870 = 10'h156 == _T_6[9:0] ? _ram_T_25[287:0] : ram_342; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_871 = 10'h157 == _T_6[9:0] ? _ram_T_25[287:0] : ram_343; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_872 = 10'h158 == _T_6[9:0] ? _ram_T_25[287:0] : ram_344; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_873 = 10'h159 == _T_6[9:0] ? _ram_T_25[287:0] : ram_345; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_874 = 10'h15a == _T_6[9:0] ? _ram_T_25[287:0] : ram_346; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_875 = 10'h15b == _T_6[9:0] ? _ram_T_25[287:0] : ram_347; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_876 = 10'h15c == _T_6[9:0] ? _ram_T_25[287:0] : ram_348; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_877 = 10'h15d == _T_6[9:0] ? _ram_T_25[287:0] : ram_349; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_878 = 10'h15e == _T_6[9:0] ? _ram_T_25[287:0] : ram_350; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_879 = 10'h15f == _T_6[9:0] ? _ram_T_25[287:0] : ram_351; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_880 = 10'h160 == _T_6[9:0] ? _ram_T_25[287:0] : ram_352; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_881 = 10'h161 == _T_6[9:0] ? _ram_T_25[287:0] : ram_353; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_882 = 10'h162 == _T_6[9:0] ? _ram_T_25[287:0] : ram_354; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_883 = 10'h163 == _T_6[9:0] ? _ram_T_25[287:0] : ram_355; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_884 = 10'h164 == _T_6[9:0] ? _ram_T_25[287:0] : ram_356; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_885 = 10'h165 == _T_6[9:0] ? _ram_T_25[287:0] : ram_357; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_886 = 10'h166 == _T_6[9:0] ? _ram_T_25[287:0] : ram_358; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_887 = 10'h167 == _T_6[9:0] ? _ram_T_25[287:0] : ram_359; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_888 = 10'h168 == _T_6[9:0] ? _ram_T_25[287:0] : ram_360; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_889 = 10'h169 == _T_6[9:0] ? _ram_T_25[287:0] : ram_361; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_890 = 10'h16a == _T_6[9:0] ? _ram_T_25[287:0] : ram_362; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_891 = 10'h16b == _T_6[9:0] ? _ram_T_25[287:0] : ram_363; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_892 = 10'h16c == _T_6[9:0] ? _ram_T_25[287:0] : ram_364; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_893 = 10'h16d == _T_6[9:0] ? _ram_T_25[287:0] : ram_365; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_894 = 10'h16e == _T_6[9:0] ? _ram_T_25[287:0] : ram_366; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_895 = 10'h16f == _T_6[9:0] ? _ram_T_25[287:0] : ram_367; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_896 = 10'h170 == _T_6[9:0] ? _ram_T_25[287:0] : ram_368; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_897 = 10'h171 == _T_6[9:0] ? _ram_T_25[287:0] : ram_369; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_898 = 10'h172 == _T_6[9:0] ? _ram_T_25[287:0] : ram_370; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_899 = 10'h173 == _T_6[9:0] ? _ram_T_25[287:0] : ram_371; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_900 = 10'h174 == _T_6[9:0] ? _ram_T_25[287:0] : ram_372; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_901 = 10'h175 == _T_6[9:0] ? _ram_T_25[287:0] : ram_373; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_902 = 10'h176 == _T_6[9:0] ? _ram_T_25[287:0] : ram_374; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_903 = 10'h177 == _T_6[9:0] ? _ram_T_25[287:0] : ram_375; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_904 = 10'h178 == _T_6[9:0] ? _ram_T_25[287:0] : ram_376; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_905 = 10'h179 == _T_6[9:0] ? _ram_T_25[287:0] : ram_377; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_906 = 10'h17a == _T_6[9:0] ? _ram_T_25[287:0] : ram_378; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_907 = 10'h17b == _T_6[9:0] ? _ram_T_25[287:0] : ram_379; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_908 = 10'h17c == _T_6[9:0] ? _ram_T_25[287:0] : ram_380; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_909 = 10'h17d == _T_6[9:0] ? _ram_T_25[287:0] : ram_381; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_910 = 10'h17e == _T_6[9:0] ? _ram_T_25[287:0] : ram_382; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_911 = 10'h17f == _T_6[9:0] ? _ram_T_25[287:0] : ram_383; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_912 = 10'h180 == _T_6[9:0] ? _ram_T_25[287:0] : ram_384; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_913 = 10'h181 == _T_6[9:0] ? _ram_T_25[287:0] : ram_385; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_914 = 10'h182 == _T_6[9:0] ? _ram_T_25[287:0] : ram_386; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_915 = 10'h183 == _T_6[9:0] ? _ram_T_25[287:0] : ram_387; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_916 = 10'h184 == _T_6[9:0] ? _ram_T_25[287:0] : ram_388; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_917 = 10'h185 == _T_6[9:0] ? _ram_T_25[287:0] : ram_389; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_918 = 10'h186 == _T_6[9:0] ? _ram_T_25[287:0] : ram_390; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_919 = 10'h187 == _T_6[9:0] ? _ram_T_25[287:0] : ram_391; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_920 = 10'h188 == _T_6[9:0] ? _ram_T_25[287:0] : ram_392; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_921 = 10'h189 == _T_6[9:0] ? _ram_T_25[287:0] : ram_393; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_922 = 10'h18a == _T_6[9:0] ? _ram_T_25[287:0] : ram_394; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_923 = 10'h18b == _T_6[9:0] ? _ram_T_25[287:0] : ram_395; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_924 = 10'h18c == _T_6[9:0] ? _ram_T_25[287:0] : ram_396; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_925 = 10'h18d == _T_6[9:0] ? _ram_T_25[287:0] : ram_397; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_926 = 10'h18e == _T_6[9:0] ? _ram_T_25[287:0] : ram_398; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_927 = 10'h18f == _T_6[9:0] ? _ram_T_25[287:0] : ram_399; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_928 = 10'h190 == _T_6[9:0] ? _ram_T_25[287:0] : ram_400; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_929 = 10'h191 == _T_6[9:0] ? _ram_T_25[287:0] : ram_401; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_930 = 10'h192 == _T_6[9:0] ? _ram_T_25[287:0] : ram_402; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_931 = 10'h193 == _T_6[9:0] ? _ram_T_25[287:0] : ram_403; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_932 = 10'h194 == _T_6[9:0] ? _ram_T_25[287:0] : ram_404; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_933 = 10'h195 == _T_6[9:0] ? _ram_T_25[287:0] : ram_405; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_934 = 10'h196 == _T_6[9:0] ? _ram_T_25[287:0] : ram_406; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_935 = 10'h197 == _T_6[9:0] ? _ram_T_25[287:0] : ram_407; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_936 = 10'h198 == _T_6[9:0] ? _ram_T_25[287:0] : ram_408; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_937 = 10'h199 == _T_6[9:0] ? _ram_T_25[287:0] : ram_409; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_938 = 10'h19a == _T_6[9:0] ? _ram_T_25[287:0] : ram_410; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_939 = 10'h19b == _T_6[9:0] ? _ram_T_25[287:0] : ram_411; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_940 = 10'h19c == _T_6[9:0] ? _ram_T_25[287:0] : ram_412; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_941 = 10'h19d == _T_6[9:0] ? _ram_T_25[287:0] : ram_413; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_942 = 10'h19e == _T_6[9:0] ? _ram_T_25[287:0] : ram_414; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_943 = 10'h19f == _T_6[9:0] ? _ram_T_25[287:0] : ram_415; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_944 = 10'h1a0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_416; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_945 = 10'h1a1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_417; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_946 = 10'h1a2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_418; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_947 = 10'h1a3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_419; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_948 = 10'h1a4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_420; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_949 = 10'h1a5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_421; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_950 = 10'h1a6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_422; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_951 = 10'h1a7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_423; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_952 = 10'h1a8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_424; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_953 = 10'h1a9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_425; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_954 = 10'h1aa == _T_6[9:0] ? _ram_T_25[287:0] : ram_426; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_955 = 10'h1ab == _T_6[9:0] ? _ram_T_25[287:0] : ram_427; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_956 = 10'h1ac == _T_6[9:0] ? _ram_T_25[287:0] : ram_428; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_957 = 10'h1ad == _T_6[9:0] ? _ram_T_25[287:0] : ram_429; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_958 = 10'h1ae == _T_6[9:0] ? _ram_T_25[287:0] : ram_430; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_959 = 10'h1af == _T_6[9:0] ? _ram_T_25[287:0] : ram_431; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_960 = 10'h1b0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_432; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_961 = 10'h1b1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_433; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_962 = 10'h1b2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_434; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_963 = 10'h1b3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_435; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_964 = 10'h1b4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_436; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_965 = 10'h1b5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_437; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_966 = 10'h1b6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_438; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_967 = 10'h1b7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_439; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_968 = 10'h1b8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_440; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_969 = 10'h1b9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_441; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_970 = 10'h1ba == _T_6[9:0] ? _ram_T_25[287:0] : ram_442; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_971 = 10'h1bb == _T_6[9:0] ? _ram_T_25[287:0] : ram_443; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_972 = 10'h1bc == _T_6[9:0] ? _ram_T_25[287:0] : ram_444; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_973 = 10'h1bd == _T_6[9:0] ? _ram_T_25[287:0] : ram_445; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_974 = 10'h1be == _T_6[9:0] ? _ram_T_25[287:0] : ram_446; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_975 = 10'h1bf == _T_6[9:0] ? _ram_T_25[287:0] : ram_447; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_976 = 10'h1c0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_448; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_977 = 10'h1c1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_449; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_978 = 10'h1c2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_450; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_979 = 10'h1c3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_451; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_980 = 10'h1c4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_452; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_981 = 10'h1c5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_453; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_982 = 10'h1c6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_454; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_983 = 10'h1c7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_455; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_984 = 10'h1c8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_456; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_985 = 10'h1c9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_457; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_986 = 10'h1ca == _T_6[9:0] ? _ram_T_25[287:0] : ram_458; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_987 = 10'h1cb == _T_6[9:0] ? _ram_T_25[287:0] : ram_459; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_988 = 10'h1cc == _T_6[9:0] ? _ram_T_25[287:0] : ram_460; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_989 = 10'h1cd == _T_6[9:0] ? _ram_T_25[287:0] : ram_461; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_990 = 10'h1ce == _T_6[9:0] ? _ram_T_25[287:0] : ram_462; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_991 = 10'h1cf == _T_6[9:0] ? _ram_T_25[287:0] : ram_463; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_992 = 10'h1d0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_464; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_993 = 10'h1d1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_465; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_994 = 10'h1d2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_466; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_995 = 10'h1d3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_467; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_996 = 10'h1d4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_468; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_997 = 10'h1d5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_469; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_998 = 10'h1d6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_470; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_999 = 10'h1d7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_471; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1000 = 10'h1d8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_472; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1001 = 10'h1d9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_473; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1002 = 10'h1da == _T_6[9:0] ? _ram_T_25[287:0] : ram_474; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1003 = 10'h1db == _T_6[9:0] ? _ram_T_25[287:0] : ram_475; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1004 = 10'h1dc == _T_6[9:0] ? _ram_T_25[287:0] : ram_476; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1005 = 10'h1dd == _T_6[9:0] ? _ram_T_25[287:0] : ram_477; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1006 = 10'h1de == _T_6[9:0] ? _ram_T_25[287:0] : ram_478; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1007 = 10'h1df == _T_6[9:0] ? _ram_T_25[287:0] : ram_479; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1008 = 10'h1e0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_480; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1009 = 10'h1e1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_481; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1010 = 10'h1e2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_482; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1011 = 10'h1e3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_483; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1012 = 10'h1e4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_484; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1013 = 10'h1e5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_485; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1014 = 10'h1e6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_486; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1015 = 10'h1e7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_487; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1016 = 10'h1e8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_488; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1017 = 10'h1e9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_489; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1018 = 10'h1ea == _T_6[9:0] ? _ram_T_25[287:0] : ram_490; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1019 = 10'h1eb == _T_6[9:0] ? _ram_T_25[287:0] : ram_491; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1020 = 10'h1ec == _T_6[9:0] ? _ram_T_25[287:0] : ram_492; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1021 = 10'h1ed == _T_6[9:0] ? _ram_T_25[287:0] : ram_493; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1022 = 10'h1ee == _T_6[9:0] ? _ram_T_25[287:0] : ram_494; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1023 = 10'h1ef == _T_6[9:0] ? _ram_T_25[287:0] : ram_495; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1024 = 10'h1f0 == _T_6[9:0] ? _ram_T_25[287:0] : ram_496; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1025 = 10'h1f1 == _T_6[9:0] ? _ram_T_25[287:0] : ram_497; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1026 = 10'h1f2 == _T_6[9:0] ? _ram_T_25[287:0] : ram_498; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1027 = 10'h1f3 == _T_6[9:0] ? _ram_T_25[287:0] : ram_499; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1028 = 10'h1f4 == _T_6[9:0] ? _ram_T_25[287:0] : ram_500; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1029 = 10'h1f5 == _T_6[9:0] ? _ram_T_25[287:0] : ram_501; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1030 = 10'h1f6 == _T_6[9:0] ? _ram_T_25[287:0] : ram_502; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1031 = 10'h1f7 == _T_6[9:0] ? _ram_T_25[287:0] : ram_503; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1032 = 10'h1f8 == _T_6[9:0] ? _ram_T_25[287:0] : ram_504; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1033 = 10'h1f9 == _T_6[9:0] ? _ram_T_25[287:0] : ram_505; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1034 = 10'h1fa == _T_6[9:0] ? _ram_T_25[287:0] : ram_506; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1035 = 10'h1fb == _T_6[9:0] ? _ram_T_25[287:0] : ram_507; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1036 = 10'h1fc == _T_6[9:0] ? _ram_T_25[287:0] : ram_508; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1037 = 10'h1fd == _T_6[9:0] ? _ram_T_25[287:0] : ram_509; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1038 = 10'h1fe == _T_6[9:0] ? _ram_T_25[287:0] : ram_510; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1039 = 10'h1ff == _T_6[9:0] ? _ram_T_25[287:0] : ram_511; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1040 = 10'h200 == _T_6[9:0] ? _ram_T_25[287:0] : ram_512; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1041 = 10'h201 == _T_6[9:0] ? _ram_T_25[287:0] : ram_513; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1042 = 10'h202 == _T_6[9:0] ? _ram_T_25[287:0] : ram_514; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1043 = 10'h203 == _T_6[9:0] ? _ram_T_25[287:0] : ram_515; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1044 = 10'h204 == _T_6[9:0] ? _ram_T_25[287:0] : ram_516; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1045 = 10'h205 == _T_6[9:0] ? _ram_T_25[287:0] : ram_517; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1046 = 10'h206 == _T_6[9:0] ? _ram_T_25[287:0] : ram_518; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1047 = 10'h207 == _T_6[9:0] ? _ram_T_25[287:0] : ram_519; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1048 = 10'h208 == _T_6[9:0] ? _ram_T_25[287:0] : ram_520; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1049 = 10'h209 == _T_6[9:0] ? _ram_T_25[287:0] : ram_521; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1050 = 10'h20a == _T_6[9:0] ? _ram_T_25[287:0] : ram_522; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1051 = 10'h20b == _T_6[9:0] ? _ram_T_25[287:0] : ram_523; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [287:0] _GEN_1052 = 10'h20c == _T_6[9:0] ? _ram_T_25[287:0] : ram_524; // @[vga.scala 64:24 vga.scala 64:24 vga.scala 46:20]
  wire [9:0] _T_9 = h + 10'h1; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_1 = vga_mem_ram_MPORT_9_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_1 = vga_mem_ram_MPORT_10_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_1 = vga_mem_ram_MPORT_11_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_1 = vga_mem_ram_MPORT_12_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_1 = vga_mem_ram_MPORT_13_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_1 = vga_mem_ram_MPORT_14_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_1 = vga_mem_ram_MPORT_15_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_1 = vga_mem_ram_MPORT_16_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_1 = vga_mem_ram_MPORT_17_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_46 = {278'h0,ram_hi_hi_hi_lo_1,ram_hi_hi_lo_1,ram_hi_lo_hi_1,ram_hi_lo_lo_1,ram_lo_hi_hi_hi_1,
    ram_lo_hi_hi_lo_1,ram_lo_hi_lo_1,ram_lo_lo_hi_1,ram_lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19062 = {{8191'd0}, _ram_T_46}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_50 = _GEN_19062 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_1054 = 10'h1 == _T_9 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1055 = 10'h2 == _T_9 ? ram_2 : _GEN_1054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1056 = 10'h3 == _T_9 ? ram_3 : _GEN_1055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1057 = 10'h4 == _T_9 ? ram_4 : _GEN_1056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1058 = 10'h5 == _T_9 ? ram_5 : _GEN_1057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1059 = 10'h6 == _T_9 ? ram_6 : _GEN_1058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1060 = 10'h7 == _T_9 ? ram_7 : _GEN_1059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1061 = 10'h8 == _T_9 ? ram_8 : _GEN_1060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1062 = 10'h9 == _T_9 ? ram_9 : _GEN_1061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1063 = 10'ha == _T_9 ? ram_10 : _GEN_1062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1064 = 10'hb == _T_9 ? ram_11 : _GEN_1063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1065 = 10'hc == _T_9 ? ram_12 : _GEN_1064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1066 = 10'hd == _T_9 ? ram_13 : _GEN_1065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1067 = 10'he == _T_9 ? ram_14 : _GEN_1066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1068 = 10'hf == _T_9 ? ram_15 : _GEN_1067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1069 = 10'h10 == _T_9 ? ram_16 : _GEN_1068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1070 = 10'h11 == _T_9 ? ram_17 : _GEN_1069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1071 = 10'h12 == _T_9 ? ram_18 : _GEN_1070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1072 = 10'h13 == _T_9 ? ram_19 : _GEN_1071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1073 = 10'h14 == _T_9 ? ram_20 : _GEN_1072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1074 = 10'h15 == _T_9 ? ram_21 : _GEN_1073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1075 = 10'h16 == _T_9 ? ram_22 : _GEN_1074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1076 = 10'h17 == _T_9 ? ram_23 : _GEN_1075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1077 = 10'h18 == _T_9 ? ram_24 : _GEN_1076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1078 = 10'h19 == _T_9 ? ram_25 : _GEN_1077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1079 = 10'h1a == _T_9 ? ram_26 : _GEN_1078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1080 = 10'h1b == _T_9 ? ram_27 : _GEN_1079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1081 = 10'h1c == _T_9 ? ram_28 : _GEN_1080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1082 = 10'h1d == _T_9 ? ram_29 : _GEN_1081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1083 = 10'h1e == _T_9 ? ram_30 : _GEN_1082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1084 = 10'h1f == _T_9 ? ram_31 : _GEN_1083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1085 = 10'h20 == _T_9 ? ram_32 : _GEN_1084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1086 = 10'h21 == _T_9 ? ram_33 : _GEN_1085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1087 = 10'h22 == _T_9 ? ram_34 : _GEN_1086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1088 = 10'h23 == _T_9 ? ram_35 : _GEN_1087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1089 = 10'h24 == _T_9 ? ram_36 : _GEN_1088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1090 = 10'h25 == _T_9 ? ram_37 : _GEN_1089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1091 = 10'h26 == _T_9 ? ram_38 : _GEN_1090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1092 = 10'h27 == _T_9 ? ram_39 : _GEN_1091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1093 = 10'h28 == _T_9 ? ram_40 : _GEN_1092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1094 = 10'h29 == _T_9 ? ram_41 : _GEN_1093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1095 = 10'h2a == _T_9 ? ram_42 : _GEN_1094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1096 = 10'h2b == _T_9 ? ram_43 : _GEN_1095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1097 = 10'h2c == _T_9 ? ram_44 : _GEN_1096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1098 = 10'h2d == _T_9 ? ram_45 : _GEN_1097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1099 = 10'h2e == _T_9 ? ram_46 : _GEN_1098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1100 = 10'h2f == _T_9 ? ram_47 : _GEN_1099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1101 = 10'h30 == _T_9 ? ram_48 : _GEN_1100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1102 = 10'h31 == _T_9 ? ram_49 : _GEN_1101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1103 = 10'h32 == _T_9 ? ram_50 : _GEN_1102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1104 = 10'h33 == _T_9 ? ram_51 : _GEN_1103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1105 = 10'h34 == _T_9 ? ram_52 : _GEN_1104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1106 = 10'h35 == _T_9 ? ram_53 : _GEN_1105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1107 = 10'h36 == _T_9 ? ram_54 : _GEN_1106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1108 = 10'h37 == _T_9 ? ram_55 : _GEN_1107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1109 = 10'h38 == _T_9 ? ram_56 : _GEN_1108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1110 = 10'h39 == _T_9 ? ram_57 : _GEN_1109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1111 = 10'h3a == _T_9 ? ram_58 : _GEN_1110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1112 = 10'h3b == _T_9 ? ram_59 : _GEN_1111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1113 = 10'h3c == _T_9 ? ram_60 : _GEN_1112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1114 = 10'h3d == _T_9 ? ram_61 : _GEN_1113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1115 = 10'h3e == _T_9 ? ram_62 : _GEN_1114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1116 = 10'h3f == _T_9 ? ram_63 : _GEN_1115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1117 = 10'h40 == _T_9 ? ram_64 : _GEN_1116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1118 = 10'h41 == _T_9 ? ram_65 : _GEN_1117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1119 = 10'h42 == _T_9 ? ram_66 : _GEN_1118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1120 = 10'h43 == _T_9 ? ram_67 : _GEN_1119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1121 = 10'h44 == _T_9 ? ram_68 : _GEN_1120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1122 = 10'h45 == _T_9 ? ram_69 : _GEN_1121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1123 = 10'h46 == _T_9 ? ram_70 : _GEN_1122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1124 = 10'h47 == _T_9 ? ram_71 : _GEN_1123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1125 = 10'h48 == _T_9 ? ram_72 : _GEN_1124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1126 = 10'h49 == _T_9 ? ram_73 : _GEN_1125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1127 = 10'h4a == _T_9 ? ram_74 : _GEN_1126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1128 = 10'h4b == _T_9 ? ram_75 : _GEN_1127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1129 = 10'h4c == _T_9 ? ram_76 : _GEN_1128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1130 = 10'h4d == _T_9 ? ram_77 : _GEN_1129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1131 = 10'h4e == _T_9 ? ram_78 : _GEN_1130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1132 = 10'h4f == _T_9 ? ram_79 : _GEN_1131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1133 = 10'h50 == _T_9 ? ram_80 : _GEN_1132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1134 = 10'h51 == _T_9 ? ram_81 : _GEN_1133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1135 = 10'h52 == _T_9 ? ram_82 : _GEN_1134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1136 = 10'h53 == _T_9 ? ram_83 : _GEN_1135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1137 = 10'h54 == _T_9 ? ram_84 : _GEN_1136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1138 = 10'h55 == _T_9 ? ram_85 : _GEN_1137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1139 = 10'h56 == _T_9 ? ram_86 : _GEN_1138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1140 = 10'h57 == _T_9 ? ram_87 : _GEN_1139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1141 = 10'h58 == _T_9 ? ram_88 : _GEN_1140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1142 = 10'h59 == _T_9 ? ram_89 : _GEN_1141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1143 = 10'h5a == _T_9 ? ram_90 : _GEN_1142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1144 = 10'h5b == _T_9 ? ram_91 : _GEN_1143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1145 = 10'h5c == _T_9 ? ram_92 : _GEN_1144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1146 = 10'h5d == _T_9 ? ram_93 : _GEN_1145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1147 = 10'h5e == _T_9 ? ram_94 : _GEN_1146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1148 = 10'h5f == _T_9 ? ram_95 : _GEN_1147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1149 = 10'h60 == _T_9 ? ram_96 : _GEN_1148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1150 = 10'h61 == _T_9 ? ram_97 : _GEN_1149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1151 = 10'h62 == _T_9 ? ram_98 : _GEN_1150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1152 = 10'h63 == _T_9 ? ram_99 : _GEN_1151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1153 = 10'h64 == _T_9 ? ram_100 : _GEN_1152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1154 = 10'h65 == _T_9 ? ram_101 : _GEN_1153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1155 = 10'h66 == _T_9 ? ram_102 : _GEN_1154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1156 = 10'h67 == _T_9 ? ram_103 : _GEN_1155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1157 = 10'h68 == _T_9 ? ram_104 : _GEN_1156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1158 = 10'h69 == _T_9 ? ram_105 : _GEN_1157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1159 = 10'h6a == _T_9 ? ram_106 : _GEN_1158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1160 = 10'h6b == _T_9 ? ram_107 : _GEN_1159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1161 = 10'h6c == _T_9 ? ram_108 : _GEN_1160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1162 = 10'h6d == _T_9 ? ram_109 : _GEN_1161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1163 = 10'h6e == _T_9 ? ram_110 : _GEN_1162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1164 = 10'h6f == _T_9 ? ram_111 : _GEN_1163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1165 = 10'h70 == _T_9 ? ram_112 : _GEN_1164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1166 = 10'h71 == _T_9 ? ram_113 : _GEN_1165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1167 = 10'h72 == _T_9 ? ram_114 : _GEN_1166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1168 = 10'h73 == _T_9 ? ram_115 : _GEN_1167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1169 = 10'h74 == _T_9 ? ram_116 : _GEN_1168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1170 = 10'h75 == _T_9 ? ram_117 : _GEN_1169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1171 = 10'h76 == _T_9 ? ram_118 : _GEN_1170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1172 = 10'h77 == _T_9 ? ram_119 : _GEN_1171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1173 = 10'h78 == _T_9 ? ram_120 : _GEN_1172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1174 = 10'h79 == _T_9 ? ram_121 : _GEN_1173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1175 = 10'h7a == _T_9 ? ram_122 : _GEN_1174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1176 = 10'h7b == _T_9 ? ram_123 : _GEN_1175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1177 = 10'h7c == _T_9 ? ram_124 : _GEN_1176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1178 = 10'h7d == _T_9 ? ram_125 : _GEN_1177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1179 = 10'h7e == _T_9 ? ram_126 : _GEN_1178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1180 = 10'h7f == _T_9 ? ram_127 : _GEN_1179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1181 = 10'h80 == _T_9 ? ram_128 : _GEN_1180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1182 = 10'h81 == _T_9 ? ram_129 : _GEN_1181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1183 = 10'h82 == _T_9 ? ram_130 : _GEN_1182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1184 = 10'h83 == _T_9 ? ram_131 : _GEN_1183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1185 = 10'h84 == _T_9 ? ram_132 : _GEN_1184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1186 = 10'h85 == _T_9 ? ram_133 : _GEN_1185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1187 = 10'h86 == _T_9 ? ram_134 : _GEN_1186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1188 = 10'h87 == _T_9 ? ram_135 : _GEN_1187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1189 = 10'h88 == _T_9 ? ram_136 : _GEN_1188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1190 = 10'h89 == _T_9 ? ram_137 : _GEN_1189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1191 = 10'h8a == _T_9 ? ram_138 : _GEN_1190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1192 = 10'h8b == _T_9 ? ram_139 : _GEN_1191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1193 = 10'h8c == _T_9 ? ram_140 : _GEN_1192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1194 = 10'h8d == _T_9 ? ram_141 : _GEN_1193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1195 = 10'h8e == _T_9 ? ram_142 : _GEN_1194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1196 = 10'h8f == _T_9 ? ram_143 : _GEN_1195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1197 = 10'h90 == _T_9 ? ram_144 : _GEN_1196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1198 = 10'h91 == _T_9 ? ram_145 : _GEN_1197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1199 = 10'h92 == _T_9 ? ram_146 : _GEN_1198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1200 = 10'h93 == _T_9 ? ram_147 : _GEN_1199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1201 = 10'h94 == _T_9 ? ram_148 : _GEN_1200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1202 = 10'h95 == _T_9 ? ram_149 : _GEN_1201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1203 = 10'h96 == _T_9 ? ram_150 : _GEN_1202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1204 = 10'h97 == _T_9 ? ram_151 : _GEN_1203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1205 = 10'h98 == _T_9 ? ram_152 : _GEN_1204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1206 = 10'h99 == _T_9 ? ram_153 : _GEN_1205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1207 = 10'h9a == _T_9 ? ram_154 : _GEN_1206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1208 = 10'h9b == _T_9 ? ram_155 : _GEN_1207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1209 = 10'h9c == _T_9 ? ram_156 : _GEN_1208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1210 = 10'h9d == _T_9 ? ram_157 : _GEN_1209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1211 = 10'h9e == _T_9 ? ram_158 : _GEN_1210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1212 = 10'h9f == _T_9 ? ram_159 : _GEN_1211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1213 = 10'ha0 == _T_9 ? ram_160 : _GEN_1212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1214 = 10'ha1 == _T_9 ? ram_161 : _GEN_1213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1215 = 10'ha2 == _T_9 ? ram_162 : _GEN_1214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1216 = 10'ha3 == _T_9 ? ram_163 : _GEN_1215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1217 = 10'ha4 == _T_9 ? ram_164 : _GEN_1216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1218 = 10'ha5 == _T_9 ? ram_165 : _GEN_1217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1219 = 10'ha6 == _T_9 ? ram_166 : _GEN_1218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1220 = 10'ha7 == _T_9 ? ram_167 : _GEN_1219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1221 = 10'ha8 == _T_9 ? ram_168 : _GEN_1220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1222 = 10'ha9 == _T_9 ? ram_169 : _GEN_1221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1223 = 10'haa == _T_9 ? ram_170 : _GEN_1222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1224 = 10'hab == _T_9 ? ram_171 : _GEN_1223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1225 = 10'hac == _T_9 ? ram_172 : _GEN_1224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1226 = 10'had == _T_9 ? ram_173 : _GEN_1225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1227 = 10'hae == _T_9 ? ram_174 : _GEN_1226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1228 = 10'haf == _T_9 ? ram_175 : _GEN_1227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1229 = 10'hb0 == _T_9 ? ram_176 : _GEN_1228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1230 = 10'hb1 == _T_9 ? ram_177 : _GEN_1229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1231 = 10'hb2 == _T_9 ? ram_178 : _GEN_1230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1232 = 10'hb3 == _T_9 ? ram_179 : _GEN_1231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1233 = 10'hb4 == _T_9 ? ram_180 : _GEN_1232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1234 = 10'hb5 == _T_9 ? ram_181 : _GEN_1233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1235 = 10'hb6 == _T_9 ? ram_182 : _GEN_1234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1236 = 10'hb7 == _T_9 ? ram_183 : _GEN_1235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1237 = 10'hb8 == _T_9 ? ram_184 : _GEN_1236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1238 = 10'hb9 == _T_9 ? ram_185 : _GEN_1237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1239 = 10'hba == _T_9 ? ram_186 : _GEN_1238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1240 = 10'hbb == _T_9 ? ram_187 : _GEN_1239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1241 = 10'hbc == _T_9 ? ram_188 : _GEN_1240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1242 = 10'hbd == _T_9 ? ram_189 : _GEN_1241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1243 = 10'hbe == _T_9 ? ram_190 : _GEN_1242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1244 = 10'hbf == _T_9 ? ram_191 : _GEN_1243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1245 = 10'hc0 == _T_9 ? ram_192 : _GEN_1244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1246 = 10'hc1 == _T_9 ? ram_193 : _GEN_1245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1247 = 10'hc2 == _T_9 ? ram_194 : _GEN_1246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1248 = 10'hc3 == _T_9 ? ram_195 : _GEN_1247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1249 = 10'hc4 == _T_9 ? ram_196 : _GEN_1248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1250 = 10'hc5 == _T_9 ? ram_197 : _GEN_1249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1251 = 10'hc6 == _T_9 ? ram_198 : _GEN_1250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1252 = 10'hc7 == _T_9 ? ram_199 : _GEN_1251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1253 = 10'hc8 == _T_9 ? ram_200 : _GEN_1252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1254 = 10'hc9 == _T_9 ? ram_201 : _GEN_1253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1255 = 10'hca == _T_9 ? ram_202 : _GEN_1254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1256 = 10'hcb == _T_9 ? ram_203 : _GEN_1255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1257 = 10'hcc == _T_9 ? ram_204 : _GEN_1256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1258 = 10'hcd == _T_9 ? ram_205 : _GEN_1257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1259 = 10'hce == _T_9 ? ram_206 : _GEN_1258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1260 = 10'hcf == _T_9 ? ram_207 : _GEN_1259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1261 = 10'hd0 == _T_9 ? ram_208 : _GEN_1260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1262 = 10'hd1 == _T_9 ? ram_209 : _GEN_1261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1263 = 10'hd2 == _T_9 ? ram_210 : _GEN_1262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1264 = 10'hd3 == _T_9 ? ram_211 : _GEN_1263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1265 = 10'hd4 == _T_9 ? ram_212 : _GEN_1264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1266 = 10'hd5 == _T_9 ? ram_213 : _GEN_1265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1267 = 10'hd6 == _T_9 ? ram_214 : _GEN_1266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1268 = 10'hd7 == _T_9 ? ram_215 : _GEN_1267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1269 = 10'hd8 == _T_9 ? ram_216 : _GEN_1268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1270 = 10'hd9 == _T_9 ? ram_217 : _GEN_1269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1271 = 10'hda == _T_9 ? ram_218 : _GEN_1270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1272 = 10'hdb == _T_9 ? ram_219 : _GEN_1271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1273 = 10'hdc == _T_9 ? ram_220 : _GEN_1272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1274 = 10'hdd == _T_9 ? ram_221 : _GEN_1273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1275 = 10'hde == _T_9 ? ram_222 : _GEN_1274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1276 = 10'hdf == _T_9 ? ram_223 : _GEN_1275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1277 = 10'he0 == _T_9 ? ram_224 : _GEN_1276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1278 = 10'he1 == _T_9 ? ram_225 : _GEN_1277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1279 = 10'he2 == _T_9 ? ram_226 : _GEN_1278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1280 = 10'he3 == _T_9 ? ram_227 : _GEN_1279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1281 = 10'he4 == _T_9 ? ram_228 : _GEN_1280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1282 = 10'he5 == _T_9 ? ram_229 : _GEN_1281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1283 = 10'he6 == _T_9 ? ram_230 : _GEN_1282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1284 = 10'he7 == _T_9 ? ram_231 : _GEN_1283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1285 = 10'he8 == _T_9 ? ram_232 : _GEN_1284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1286 = 10'he9 == _T_9 ? ram_233 : _GEN_1285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1287 = 10'hea == _T_9 ? ram_234 : _GEN_1286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1288 = 10'heb == _T_9 ? ram_235 : _GEN_1287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1289 = 10'hec == _T_9 ? ram_236 : _GEN_1288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1290 = 10'hed == _T_9 ? ram_237 : _GEN_1289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1291 = 10'hee == _T_9 ? ram_238 : _GEN_1290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1292 = 10'hef == _T_9 ? ram_239 : _GEN_1291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1293 = 10'hf0 == _T_9 ? ram_240 : _GEN_1292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1294 = 10'hf1 == _T_9 ? ram_241 : _GEN_1293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1295 = 10'hf2 == _T_9 ? ram_242 : _GEN_1294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1296 = 10'hf3 == _T_9 ? ram_243 : _GEN_1295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1297 = 10'hf4 == _T_9 ? ram_244 : _GEN_1296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1298 = 10'hf5 == _T_9 ? ram_245 : _GEN_1297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1299 = 10'hf6 == _T_9 ? ram_246 : _GEN_1298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1300 = 10'hf7 == _T_9 ? ram_247 : _GEN_1299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1301 = 10'hf8 == _T_9 ? ram_248 : _GEN_1300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1302 = 10'hf9 == _T_9 ? ram_249 : _GEN_1301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1303 = 10'hfa == _T_9 ? ram_250 : _GEN_1302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1304 = 10'hfb == _T_9 ? ram_251 : _GEN_1303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1305 = 10'hfc == _T_9 ? ram_252 : _GEN_1304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1306 = 10'hfd == _T_9 ? ram_253 : _GEN_1305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1307 = 10'hfe == _T_9 ? ram_254 : _GEN_1306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1308 = 10'hff == _T_9 ? ram_255 : _GEN_1307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1309 = 10'h100 == _T_9 ? ram_256 : _GEN_1308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1310 = 10'h101 == _T_9 ? ram_257 : _GEN_1309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1311 = 10'h102 == _T_9 ? ram_258 : _GEN_1310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1312 = 10'h103 == _T_9 ? ram_259 : _GEN_1311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1313 = 10'h104 == _T_9 ? ram_260 : _GEN_1312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1314 = 10'h105 == _T_9 ? ram_261 : _GEN_1313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1315 = 10'h106 == _T_9 ? ram_262 : _GEN_1314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1316 = 10'h107 == _T_9 ? ram_263 : _GEN_1315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1317 = 10'h108 == _T_9 ? ram_264 : _GEN_1316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1318 = 10'h109 == _T_9 ? ram_265 : _GEN_1317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1319 = 10'h10a == _T_9 ? ram_266 : _GEN_1318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1320 = 10'h10b == _T_9 ? ram_267 : _GEN_1319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1321 = 10'h10c == _T_9 ? ram_268 : _GEN_1320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1322 = 10'h10d == _T_9 ? ram_269 : _GEN_1321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1323 = 10'h10e == _T_9 ? ram_270 : _GEN_1322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1324 = 10'h10f == _T_9 ? ram_271 : _GEN_1323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1325 = 10'h110 == _T_9 ? ram_272 : _GEN_1324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1326 = 10'h111 == _T_9 ? ram_273 : _GEN_1325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1327 = 10'h112 == _T_9 ? ram_274 : _GEN_1326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1328 = 10'h113 == _T_9 ? ram_275 : _GEN_1327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1329 = 10'h114 == _T_9 ? ram_276 : _GEN_1328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1330 = 10'h115 == _T_9 ? ram_277 : _GEN_1329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1331 = 10'h116 == _T_9 ? ram_278 : _GEN_1330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1332 = 10'h117 == _T_9 ? ram_279 : _GEN_1331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1333 = 10'h118 == _T_9 ? ram_280 : _GEN_1332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1334 = 10'h119 == _T_9 ? ram_281 : _GEN_1333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1335 = 10'h11a == _T_9 ? ram_282 : _GEN_1334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1336 = 10'h11b == _T_9 ? ram_283 : _GEN_1335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1337 = 10'h11c == _T_9 ? ram_284 : _GEN_1336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1338 = 10'h11d == _T_9 ? ram_285 : _GEN_1337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1339 = 10'h11e == _T_9 ? ram_286 : _GEN_1338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1340 = 10'h11f == _T_9 ? ram_287 : _GEN_1339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1341 = 10'h120 == _T_9 ? ram_288 : _GEN_1340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1342 = 10'h121 == _T_9 ? ram_289 : _GEN_1341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1343 = 10'h122 == _T_9 ? ram_290 : _GEN_1342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1344 = 10'h123 == _T_9 ? ram_291 : _GEN_1343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1345 = 10'h124 == _T_9 ? ram_292 : _GEN_1344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1346 = 10'h125 == _T_9 ? ram_293 : _GEN_1345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1347 = 10'h126 == _T_9 ? ram_294 : _GEN_1346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1348 = 10'h127 == _T_9 ? ram_295 : _GEN_1347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1349 = 10'h128 == _T_9 ? ram_296 : _GEN_1348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1350 = 10'h129 == _T_9 ? ram_297 : _GEN_1349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1351 = 10'h12a == _T_9 ? ram_298 : _GEN_1350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1352 = 10'h12b == _T_9 ? ram_299 : _GEN_1351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1353 = 10'h12c == _T_9 ? ram_300 : _GEN_1352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1354 = 10'h12d == _T_9 ? ram_301 : _GEN_1353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1355 = 10'h12e == _T_9 ? ram_302 : _GEN_1354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1356 = 10'h12f == _T_9 ? ram_303 : _GEN_1355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1357 = 10'h130 == _T_9 ? ram_304 : _GEN_1356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1358 = 10'h131 == _T_9 ? ram_305 : _GEN_1357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1359 = 10'h132 == _T_9 ? ram_306 : _GEN_1358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1360 = 10'h133 == _T_9 ? ram_307 : _GEN_1359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1361 = 10'h134 == _T_9 ? ram_308 : _GEN_1360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1362 = 10'h135 == _T_9 ? ram_309 : _GEN_1361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1363 = 10'h136 == _T_9 ? ram_310 : _GEN_1362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1364 = 10'h137 == _T_9 ? ram_311 : _GEN_1363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1365 = 10'h138 == _T_9 ? ram_312 : _GEN_1364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1366 = 10'h139 == _T_9 ? ram_313 : _GEN_1365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1367 = 10'h13a == _T_9 ? ram_314 : _GEN_1366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1368 = 10'h13b == _T_9 ? ram_315 : _GEN_1367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1369 = 10'h13c == _T_9 ? ram_316 : _GEN_1368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1370 = 10'h13d == _T_9 ? ram_317 : _GEN_1369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1371 = 10'h13e == _T_9 ? ram_318 : _GEN_1370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1372 = 10'h13f == _T_9 ? ram_319 : _GEN_1371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1373 = 10'h140 == _T_9 ? ram_320 : _GEN_1372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1374 = 10'h141 == _T_9 ? ram_321 : _GEN_1373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1375 = 10'h142 == _T_9 ? ram_322 : _GEN_1374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1376 = 10'h143 == _T_9 ? ram_323 : _GEN_1375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1377 = 10'h144 == _T_9 ? ram_324 : _GEN_1376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1378 = 10'h145 == _T_9 ? ram_325 : _GEN_1377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1379 = 10'h146 == _T_9 ? ram_326 : _GEN_1378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1380 = 10'h147 == _T_9 ? ram_327 : _GEN_1379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1381 = 10'h148 == _T_9 ? ram_328 : _GEN_1380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1382 = 10'h149 == _T_9 ? ram_329 : _GEN_1381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1383 = 10'h14a == _T_9 ? ram_330 : _GEN_1382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1384 = 10'h14b == _T_9 ? ram_331 : _GEN_1383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1385 = 10'h14c == _T_9 ? ram_332 : _GEN_1384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1386 = 10'h14d == _T_9 ? ram_333 : _GEN_1385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1387 = 10'h14e == _T_9 ? ram_334 : _GEN_1386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1388 = 10'h14f == _T_9 ? ram_335 : _GEN_1387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1389 = 10'h150 == _T_9 ? ram_336 : _GEN_1388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1390 = 10'h151 == _T_9 ? ram_337 : _GEN_1389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1391 = 10'h152 == _T_9 ? ram_338 : _GEN_1390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1392 = 10'h153 == _T_9 ? ram_339 : _GEN_1391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1393 = 10'h154 == _T_9 ? ram_340 : _GEN_1392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1394 = 10'h155 == _T_9 ? ram_341 : _GEN_1393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1395 = 10'h156 == _T_9 ? ram_342 : _GEN_1394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1396 = 10'h157 == _T_9 ? ram_343 : _GEN_1395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1397 = 10'h158 == _T_9 ? ram_344 : _GEN_1396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1398 = 10'h159 == _T_9 ? ram_345 : _GEN_1397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1399 = 10'h15a == _T_9 ? ram_346 : _GEN_1398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1400 = 10'h15b == _T_9 ? ram_347 : _GEN_1399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1401 = 10'h15c == _T_9 ? ram_348 : _GEN_1400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1402 = 10'h15d == _T_9 ? ram_349 : _GEN_1401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1403 = 10'h15e == _T_9 ? ram_350 : _GEN_1402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1404 = 10'h15f == _T_9 ? ram_351 : _GEN_1403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1405 = 10'h160 == _T_9 ? ram_352 : _GEN_1404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1406 = 10'h161 == _T_9 ? ram_353 : _GEN_1405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1407 = 10'h162 == _T_9 ? ram_354 : _GEN_1406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1408 = 10'h163 == _T_9 ? ram_355 : _GEN_1407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1409 = 10'h164 == _T_9 ? ram_356 : _GEN_1408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1410 = 10'h165 == _T_9 ? ram_357 : _GEN_1409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1411 = 10'h166 == _T_9 ? ram_358 : _GEN_1410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1412 = 10'h167 == _T_9 ? ram_359 : _GEN_1411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1413 = 10'h168 == _T_9 ? ram_360 : _GEN_1412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1414 = 10'h169 == _T_9 ? ram_361 : _GEN_1413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1415 = 10'h16a == _T_9 ? ram_362 : _GEN_1414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1416 = 10'h16b == _T_9 ? ram_363 : _GEN_1415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1417 = 10'h16c == _T_9 ? ram_364 : _GEN_1416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1418 = 10'h16d == _T_9 ? ram_365 : _GEN_1417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1419 = 10'h16e == _T_9 ? ram_366 : _GEN_1418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1420 = 10'h16f == _T_9 ? ram_367 : _GEN_1419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1421 = 10'h170 == _T_9 ? ram_368 : _GEN_1420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1422 = 10'h171 == _T_9 ? ram_369 : _GEN_1421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1423 = 10'h172 == _T_9 ? ram_370 : _GEN_1422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1424 = 10'h173 == _T_9 ? ram_371 : _GEN_1423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1425 = 10'h174 == _T_9 ? ram_372 : _GEN_1424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1426 = 10'h175 == _T_9 ? ram_373 : _GEN_1425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1427 = 10'h176 == _T_9 ? ram_374 : _GEN_1426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1428 = 10'h177 == _T_9 ? ram_375 : _GEN_1427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1429 = 10'h178 == _T_9 ? ram_376 : _GEN_1428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1430 = 10'h179 == _T_9 ? ram_377 : _GEN_1429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1431 = 10'h17a == _T_9 ? ram_378 : _GEN_1430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1432 = 10'h17b == _T_9 ? ram_379 : _GEN_1431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1433 = 10'h17c == _T_9 ? ram_380 : _GEN_1432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1434 = 10'h17d == _T_9 ? ram_381 : _GEN_1433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1435 = 10'h17e == _T_9 ? ram_382 : _GEN_1434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1436 = 10'h17f == _T_9 ? ram_383 : _GEN_1435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1437 = 10'h180 == _T_9 ? ram_384 : _GEN_1436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1438 = 10'h181 == _T_9 ? ram_385 : _GEN_1437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1439 = 10'h182 == _T_9 ? ram_386 : _GEN_1438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1440 = 10'h183 == _T_9 ? ram_387 : _GEN_1439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1441 = 10'h184 == _T_9 ? ram_388 : _GEN_1440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1442 = 10'h185 == _T_9 ? ram_389 : _GEN_1441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1443 = 10'h186 == _T_9 ? ram_390 : _GEN_1442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1444 = 10'h187 == _T_9 ? ram_391 : _GEN_1443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1445 = 10'h188 == _T_9 ? ram_392 : _GEN_1444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1446 = 10'h189 == _T_9 ? ram_393 : _GEN_1445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1447 = 10'h18a == _T_9 ? ram_394 : _GEN_1446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1448 = 10'h18b == _T_9 ? ram_395 : _GEN_1447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1449 = 10'h18c == _T_9 ? ram_396 : _GEN_1448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1450 = 10'h18d == _T_9 ? ram_397 : _GEN_1449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1451 = 10'h18e == _T_9 ? ram_398 : _GEN_1450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1452 = 10'h18f == _T_9 ? ram_399 : _GEN_1451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1453 = 10'h190 == _T_9 ? ram_400 : _GEN_1452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1454 = 10'h191 == _T_9 ? ram_401 : _GEN_1453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1455 = 10'h192 == _T_9 ? ram_402 : _GEN_1454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1456 = 10'h193 == _T_9 ? ram_403 : _GEN_1455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1457 = 10'h194 == _T_9 ? ram_404 : _GEN_1456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1458 = 10'h195 == _T_9 ? ram_405 : _GEN_1457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1459 = 10'h196 == _T_9 ? ram_406 : _GEN_1458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1460 = 10'h197 == _T_9 ? ram_407 : _GEN_1459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1461 = 10'h198 == _T_9 ? ram_408 : _GEN_1460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1462 = 10'h199 == _T_9 ? ram_409 : _GEN_1461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1463 = 10'h19a == _T_9 ? ram_410 : _GEN_1462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1464 = 10'h19b == _T_9 ? ram_411 : _GEN_1463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1465 = 10'h19c == _T_9 ? ram_412 : _GEN_1464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1466 = 10'h19d == _T_9 ? ram_413 : _GEN_1465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1467 = 10'h19e == _T_9 ? ram_414 : _GEN_1466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1468 = 10'h19f == _T_9 ? ram_415 : _GEN_1467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1469 = 10'h1a0 == _T_9 ? ram_416 : _GEN_1468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1470 = 10'h1a1 == _T_9 ? ram_417 : _GEN_1469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1471 = 10'h1a2 == _T_9 ? ram_418 : _GEN_1470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1472 = 10'h1a3 == _T_9 ? ram_419 : _GEN_1471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1473 = 10'h1a4 == _T_9 ? ram_420 : _GEN_1472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1474 = 10'h1a5 == _T_9 ? ram_421 : _GEN_1473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1475 = 10'h1a6 == _T_9 ? ram_422 : _GEN_1474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1476 = 10'h1a7 == _T_9 ? ram_423 : _GEN_1475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1477 = 10'h1a8 == _T_9 ? ram_424 : _GEN_1476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1478 = 10'h1a9 == _T_9 ? ram_425 : _GEN_1477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1479 = 10'h1aa == _T_9 ? ram_426 : _GEN_1478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1480 = 10'h1ab == _T_9 ? ram_427 : _GEN_1479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1481 = 10'h1ac == _T_9 ? ram_428 : _GEN_1480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1482 = 10'h1ad == _T_9 ? ram_429 : _GEN_1481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1483 = 10'h1ae == _T_9 ? ram_430 : _GEN_1482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1484 = 10'h1af == _T_9 ? ram_431 : _GEN_1483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1485 = 10'h1b0 == _T_9 ? ram_432 : _GEN_1484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1486 = 10'h1b1 == _T_9 ? ram_433 : _GEN_1485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1487 = 10'h1b2 == _T_9 ? ram_434 : _GEN_1486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1488 = 10'h1b3 == _T_9 ? ram_435 : _GEN_1487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1489 = 10'h1b4 == _T_9 ? ram_436 : _GEN_1488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1490 = 10'h1b5 == _T_9 ? ram_437 : _GEN_1489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1491 = 10'h1b6 == _T_9 ? ram_438 : _GEN_1490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1492 = 10'h1b7 == _T_9 ? ram_439 : _GEN_1491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1493 = 10'h1b8 == _T_9 ? ram_440 : _GEN_1492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1494 = 10'h1b9 == _T_9 ? ram_441 : _GEN_1493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1495 = 10'h1ba == _T_9 ? ram_442 : _GEN_1494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1496 = 10'h1bb == _T_9 ? ram_443 : _GEN_1495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1497 = 10'h1bc == _T_9 ? ram_444 : _GEN_1496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1498 = 10'h1bd == _T_9 ? ram_445 : _GEN_1497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1499 = 10'h1be == _T_9 ? ram_446 : _GEN_1498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1500 = 10'h1bf == _T_9 ? ram_447 : _GEN_1499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1501 = 10'h1c0 == _T_9 ? ram_448 : _GEN_1500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1502 = 10'h1c1 == _T_9 ? ram_449 : _GEN_1501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1503 = 10'h1c2 == _T_9 ? ram_450 : _GEN_1502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1504 = 10'h1c3 == _T_9 ? ram_451 : _GEN_1503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1505 = 10'h1c4 == _T_9 ? ram_452 : _GEN_1504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1506 = 10'h1c5 == _T_9 ? ram_453 : _GEN_1505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1507 = 10'h1c6 == _T_9 ? ram_454 : _GEN_1506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1508 = 10'h1c7 == _T_9 ? ram_455 : _GEN_1507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1509 = 10'h1c8 == _T_9 ? ram_456 : _GEN_1508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1510 = 10'h1c9 == _T_9 ? ram_457 : _GEN_1509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1511 = 10'h1ca == _T_9 ? ram_458 : _GEN_1510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1512 = 10'h1cb == _T_9 ? ram_459 : _GEN_1511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1513 = 10'h1cc == _T_9 ? ram_460 : _GEN_1512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1514 = 10'h1cd == _T_9 ? ram_461 : _GEN_1513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1515 = 10'h1ce == _T_9 ? ram_462 : _GEN_1514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1516 = 10'h1cf == _T_9 ? ram_463 : _GEN_1515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1517 = 10'h1d0 == _T_9 ? ram_464 : _GEN_1516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1518 = 10'h1d1 == _T_9 ? ram_465 : _GEN_1517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1519 = 10'h1d2 == _T_9 ? ram_466 : _GEN_1518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1520 = 10'h1d3 == _T_9 ? ram_467 : _GEN_1519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1521 = 10'h1d4 == _T_9 ? ram_468 : _GEN_1520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1522 = 10'h1d5 == _T_9 ? ram_469 : _GEN_1521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1523 = 10'h1d6 == _T_9 ? ram_470 : _GEN_1522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1524 = 10'h1d7 == _T_9 ? ram_471 : _GEN_1523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1525 = 10'h1d8 == _T_9 ? ram_472 : _GEN_1524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1526 = 10'h1d9 == _T_9 ? ram_473 : _GEN_1525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1527 = 10'h1da == _T_9 ? ram_474 : _GEN_1526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1528 = 10'h1db == _T_9 ? ram_475 : _GEN_1527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1529 = 10'h1dc == _T_9 ? ram_476 : _GEN_1528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1530 = 10'h1dd == _T_9 ? ram_477 : _GEN_1529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1531 = 10'h1de == _T_9 ? ram_478 : _GEN_1530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1532 = 10'h1df == _T_9 ? ram_479 : _GEN_1531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1533 = 10'h1e0 == _T_9 ? ram_480 : _GEN_1532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1534 = 10'h1e1 == _T_9 ? ram_481 : _GEN_1533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1535 = 10'h1e2 == _T_9 ? ram_482 : _GEN_1534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1536 = 10'h1e3 == _T_9 ? ram_483 : _GEN_1535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1537 = 10'h1e4 == _T_9 ? ram_484 : _GEN_1536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1538 = 10'h1e5 == _T_9 ? ram_485 : _GEN_1537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1539 = 10'h1e6 == _T_9 ? ram_486 : _GEN_1538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1540 = 10'h1e7 == _T_9 ? ram_487 : _GEN_1539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1541 = 10'h1e8 == _T_9 ? ram_488 : _GEN_1540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1542 = 10'h1e9 == _T_9 ? ram_489 : _GEN_1541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1543 = 10'h1ea == _T_9 ? ram_490 : _GEN_1542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1544 = 10'h1eb == _T_9 ? ram_491 : _GEN_1543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1545 = 10'h1ec == _T_9 ? ram_492 : _GEN_1544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1546 = 10'h1ed == _T_9 ? ram_493 : _GEN_1545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1547 = 10'h1ee == _T_9 ? ram_494 : _GEN_1546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1548 = 10'h1ef == _T_9 ? ram_495 : _GEN_1547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1549 = 10'h1f0 == _T_9 ? ram_496 : _GEN_1548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1550 = 10'h1f1 == _T_9 ? ram_497 : _GEN_1549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1551 = 10'h1f2 == _T_9 ? ram_498 : _GEN_1550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1552 = 10'h1f3 == _T_9 ? ram_499 : _GEN_1551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1553 = 10'h1f4 == _T_9 ? ram_500 : _GEN_1552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1554 = 10'h1f5 == _T_9 ? ram_501 : _GEN_1553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1555 = 10'h1f6 == _T_9 ? ram_502 : _GEN_1554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1556 = 10'h1f7 == _T_9 ? ram_503 : _GEN_1555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1557 = 10'h1f8 == _T_9 ? ram_504 : _GEN_1556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1558 = 10'h1f9 == _T_9 ? ram_505 : _GEN_1557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1559 = 10'h1fa == _T_9 ? ram_506 : _GEN_1558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1560 = 10'h1fb == _T_9 ? ram_507 : _GEN_1559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1561 = 10'h1fc == _T_9 ? ram_508 : _GEN_1560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1562 = 10'h1fd == _T_9 ? ram_509 : _GEN_1561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1563 = 10'h1fe == _T_9 ? ram_510 : _GEN_1562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1564 = 10'h1ff == _T_9 ? ram_511 : _GEN_1563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1565 = 10'h200 == _T_9 ? ram_512 : _GEN_1564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1566 = 10'h201 == _T_9 ? ram_513 : _GEN_1565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1567 = 10'h202 == _T_9 ? ram_514 : _GEN_1566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1568 = 10'h203 == _T_9 ? ram_515 : _GEN_1567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1569 = 10'h204 == _T_9 ? ram_516 : _GEN_1568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1570 = 10'h205 == _T_9 ? ram_517 : _GEN_1569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1571 = 10'h206 == _T_9 ? ram_518 : _GEN_1570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1572 = 10'h207 == _T_9 ? ram_519 : _GEN_1571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1573 = 10'h208 == _T_9 ? ram_520 : _GEN_1572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1574 = 10'h209 == _T_9 ? ram_521 : _GEN_1573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1575 = 10'h20a == _T_9 ? ram_522 : _GEN_1574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1576 = 10'h20b == _T_9 ? ram_523 : _GEN_1575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_1577 = 10'h20c == _T_9 ? ram_524 : _GEN_1576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19063 = {{8190'd0}, _GEN_1577}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_51 = _GEN_19063 ^ _ram_T_50; // @[vga.scala 64:41]
  wire [287:0] _GEN_1578 = 10'h0 == _T_9 ? _ram_T_51[287:0] : _GEN_528; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1579 = 10'h1 == _T_9 ? _ram_T_51[287:0] : _GEN_529; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1580 = 10'h2 == _T_9 ? _ram_T_51[287:0] : _GEN_530; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1581 = 10'h3 == _T_9 ? _ram_T_51[287:0] : _GEN_531; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1582 = 10'h4 == _T_9 ? _ram_T_51[287:0] : _GEN_532; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1583 = 10'h5 == _T_9 ? _ram_T_51[287:0] : _GEN_533; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1584 = 10'h6 == _T_9 ? _ram_T_51[287:0] : _GEN_534; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1585 = 10'h7 == _T_9 ? _ram_T_51[287:0] : _GEN_535; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1586 = 10'h8 == _T_9 ? _ram_T_51[287:0] : _GEN_536; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1587 = 10'h9 == _T_9 ? _ram_T_51[287:0] : _GEN_537; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1588 = 10'ha == _T_9 ? _ram_T_51[287:0] : _GEN_538; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1589 = 10'hb == _T_9 ? _ram_T_51[287:0] : _GEN_539; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1590 = 10'hc == _T_9 ? _ram_T_51[287:0] : _GEN_540; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1591 = 10'hd == _T_9 ? _ram_T_51[287:0] : _GEN_541; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1592 = 10'he == _T_9 ? _ram_T_51[287:0] : _GEN_542; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1593 = 10'hf == _T_9 ? _ram_T_51[287:0] : _GEN_543; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1594 = 10'h10 == _T_9 ? _ram_T_51[287:0] : _GEN_544; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1595 = 10'h11 == _T_9 ? _ram_T_51[287:0] : _GEN_545; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1596 = 10'h12 == _T_9 ? _ram_T_51[287:0] : _GEN_546; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1597 = 10'h13 == _T_9 ? _ram_T_51[287:0] : _GEN_547; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1598 = 10'h14 == _T_9 ? _ram_T_51[287:0] : _GEN_548; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1599 = 10'h15 == _T_9 ? _ram_T_51[287:0] : _GEN_549; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1600 = 10'h16 == _T_9 ? _ram_T_51[287:0] : _GEN_550; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1601 = 10'h17 == _T_9 ? _ram_T_51[287:0] : _GEN_551; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1602 = 10'h18 == _T_9 ? _ram_T_51[287:0] : _GEN_552; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1603 = 10'h19 == _T_9 ? _ram_T_51[287:0] : _GEN_553; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1604 = 10'h1a == _T_9 ? _ram_T_51[287:0] : _GEN_554; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1605 = 10'h1b == _T_9 ? _ram_T_51[287:0] : _GEN_555; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1606 = 10'h1c == _T_9 ? _ram_T_51[287:0] : _GEN_556; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1607 = 10'h1d == _T_9 ? _ram_T_51[287:0] : _GEN_557; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1608 = 10'h1e == _T_9 ? _ram_T_51[287:0] : _GEN_558; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1609 = 10'h1f == _T_9 ? _ram_T_51[287:0] : _GEN_559; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1610 = 10'h20 == _T_9 ? _ram_T_51[287:0] : _GEN_560; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1611 = 10'h21 == _T_9 ? _ram_T_51[287:0] : _GEN_561; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1612 = 10'h22 == _T_9 ? _ram_T_51[287:0] : _GEN_562; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1613 = 10'h23 == _T_9 ? _ram_T_51[287:0] : _GEN_563; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1614 = 10'h24 == _T_9 ? _ram_T_51[287:0] : _GEN_564; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1615 = 10'h25 == _T_9 ? _ram_T_51[287:0] : _GEN_565; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1616 = 10'h26 == _T_9 ? _ram_T_51[287:0] : _GEN_566; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1617 = 10'h27 == _T_9 ? _ram_T_51[287:0] : _GEN_567; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1618 = 10'h28 == _T_9 ? _ram_T_51[287:0] : _GEN_568; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1619 = 10'h29 == _T_9 ? _ram_T_51[287:0] : _GEN_569; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1620 = 10'h2a == _T_9 ? _ram_T_51[287:0] : _GEN_570; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1621 = 10'h2b == _T_9 ? _ram_T_51[287:0] : _GEN_571; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1622 = 10'h2c == _T_9 ? _ram_T_51[287:0] : _GEN_572; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1623 = 10'h2d == _T_9 ? _ram_T_51[287:0] : _GEN_573; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1624 = 10'h2e == _T_9 ? _ram_T_51[287:0] : _GEN_574; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1625 = 10'h2f == _T_9 ? _ram_T_51[287:0] : _GEN_575; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1626 = 10'h30 == _T_9 ? _ram_T_51[287:0] : _GEN_576; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1627 = 10'h31 == _T_9 ? _ram_T_51[287:0] : _GEN_577; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1628 = 10'h32 == _T_9 ? _ram_T_51[287:0] : _GEN_578; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1629 = 10'h33 == _T_9 ? _ram_T_51[287:0] : _GEN_579; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1630 = 10'h34 == _T_9 ? _ram_T_51[287:0] : _GEN_580; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1631 = 10'h35 == _T_9 ? _ram_T_51[287:0] : _GEN_581; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1632 = 10'h36 == _T_9 ? _ram_T_51[287:0] : _GEN_582; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1633 = 10'h37 == _T_9 ? _ram_T_51[287:0] : _GEN_583; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1634 = 10'h38 == _T_9 ? _ram_T_51[287:0] : _GEN_584; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1635 = 10'h39 == _T_9 ? _ram_T_51[287:0] : _GEN_585; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1636 = 10'h3a == _T_9 ? _ram_T_51[287:0] : _GEN_586; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1637 = 10'h3b == _T_9 ? _ram_T_51[287:0] : _GEN_587; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1638 = 10'h3c == _T_9 ? _ram_T_51[287:0] : _GEN_588; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1639 = 10'h3d == _T_9 ? _ram_T_51[287:0] : _GEN_589; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1640 = 10'h3e == _T_9 ? _ram_T_51[287:0] : _GEN_590; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1641 = 10'h3f == _T_9 ? _ram_T_51[287:0] : _GEN_591; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1642 = 10'h40 == _T_9 ? _ram_T_51[287:0] : _GEN_592; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1643 = 10'h41 == _T_9 ? _ram_T_51[287:0] : _GEN_593; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1644 = 10'h42 == _T_9 ? _ram_T_51[287:0] : _GEN_594; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1645 = 10'h43 == _T_9 ? _ram_T_51[287:0] : _GEN_595; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1646 = 10'h44 == _T_9 ? _ram_T_51[287:0] : _GEN_596; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1647 = 10'h45 == _T_9 ? _ram_T_51[287:0] : _GEN_597; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1648 = 10'h46 == _T_9 ? _ram_T_51[287:0] : _GEN_598; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1649 = 10'h47 == _T_9 ? _ram_T_51[287:0] : _GEN_599; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1650 = 10'h48 == _T_9 ? _ram_T_51[287:0] : _GEN_600; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1651 = 10'h49 == _T_9 ? _ram_T_51[287:0] : _GEN_601; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1652 = 10'h4a == _T_9 ? _ram_T_51[287:0] : _GEN_602; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1653 = 10'h4b == _T_9 ? _ram_T_51[287:0] : _GEN_603; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1654 = 10'h4c == _T_9 ? _ram_T_51[287:0] : _GEN_604; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1655 = 10'h4d == _T_9 ? _ram_T_51[287:0] : _GEN_605; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1656 = 10'h4e == _T_9 ? _ram_T_51[287:0] : _GEN_606; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1657 = 10'h4f == _T_9 ? _ram_T_51[287:0] : _GEN_607; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1658 = 10'h50 == _T_9 ? _ram_T_51[287:0] : _GEN_608; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1659 = 10'h51 == _T_9 ? _ram_T_51[287:0] : _GEN_609; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1660 = 10'h52 == _T_9 ? _ram_T_51[287:0] : _GEN_610; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1661 = 10'h53 == _T_9 ? _ram_T_51[287:0] : _GEN_611; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1662 = 10'h54 == _T_9 ? _ram_T_51[287:0] : _GEN_612; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1663 = 10'h55 == _T_9 ? _ram_T_51[287:0] : _GEN_613; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1664 = 10'h56 == _T_9 ? _ram_T_51[287:0] : _GEN_614; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1665 = 10'h57 == _T_9 ? _ram_T_51[287:0] : _GEN_615; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1666 = 10'h58 == _T_9 ? _ram_T_51[287:0] : _GEN_616; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1667 = 10'h59 == _T_9 ? _ram_T_51[287:0] : _GEN_617; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1668 = 10'h5a == _T_9 ? _ram_T_51[287:0] : _GEN_618; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1669 = 10'h5b == _T_9 ? _ram_T_51[287:0] : _GEN_619; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1670 = 10'h5c == _T_9 ? _ram_T_51[287:0] : _GEN_620; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1671 = 10'h5d == _T_9 ? _ram_T_51[287:0] : _GEN_621; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1672 = 10'h5e == _T_9 ? _ram_T_51[287:0] : _GEN_622; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1673 = 10'h5f == _T_9 ? _ram_T_51[287:0] : _GEN_623; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1674 = 10'h60 == _T_9 ? _ram_T_51[287:0] : _GEN_624; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1675 = 10'h61 == _T_9 ? _ram_T_51[287:0] : _GEN_625; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1676 = 10'h62 == _T_9 ? _ram_T_51[287:0] : _GEN_626; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1677 = 10'h63 == _T_9 ? _ram_T_51[287:0] : _GEN_627; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1678 = 10'h64 == _T_9 ? _ram_T_51[287:0] : _GEN_628; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1679 = 10'h65 == _T_9 ? _ram_T_51[287:0] : _GEN_629; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1680 = 10'h66 == _T_9 ? _ram_T_51[287:0] : _GEN_630; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1681 = 10'h67 == _T_9 ? _ram_T_51[287:0] : _GEN_631; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1682 = 10'h68 == _T_9 ? _ram_T_51[287:0] : _GEN_632; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1683 = 10'h69 == _T_9 ? _ram_T_51[287:0] : _GEN_633; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1684 = 10'h6a == _T_9 ? _ram_T_51[287:0] : _GEN_634; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1685 = 10'h6b == _T_9 ? _ram_T_51[287:0] : _GEN_635; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1686 = 10'h6c == _T_9 ? _ram_T_51[287:0] : _GEN_636; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1687 = 10'h6d == _T_9 ? _ram_T_51[287:0] : _GEN_637; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1688 = 10'h6e == _T_9 ? _ram_T_51[287:0] : _GEN_638; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1689 = 10'h6f == _T_9 ? _ram_T_51[287:0] : _GEN_639; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1690 = 10'h70 == _T_9 ? _ram_T_51[287:0] : _GEN_640; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1691 = 10'h71 == _T_9 ? _ram_T_51[287:0] : _GEN_641; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1692 = 10'h72 == _T_9 ? _ram_T_51[287:0] : _GEN_642; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1693 = 10'h73 == _T_9 ? _ram_T_51[287:0] : _GEN_643; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1694 = 10'h74 == _T_9 ? _ram_T_51[287:0] : _GEN_644; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1695 = 10'h75 == _T_9 ? _ram_T_51[287:0] : _GEN_645; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1696 = 10'h76 == _T_9 ? _ram_T_51[287:0] : _GEN_646; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1697 = 10'h77 == _T_9 ? _ram_T_51[287:0] : _GEN_647; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1698 = 10'h78 == _T_9 ? _ram_T_51[287:0] : _GEN_648; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1699 = 10'h79 == _T_9 ? _ram_T_51[287:0] : _GEN_649; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1700 = 10'h7a == _T_9 ? _ram_T_51[287:0] : _GEN_650; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1701 = 10'h7b == _T_9 ? _ram_T_51[287:0] : _GEN_651; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1702 = 10'h7c == _T_9 ? _ram_T_51[287:0] : _GEN_652; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1703 = 10'h7d == _T_9 ? _ram_T_51[287:0] : _GEN_653; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1704 = 10'h7e == _T_9 ? _ram_T_51[287:0] : _GEN_654; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1705 = 10'h7f == _T_9 ? _ram_T_51[287:0] : _GEN_655; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1706 = 10'h80 == _T_9 ? _ram_T_51[287:0] : _GEN_656; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1707 = 10'h81 == _T_9 ? _ram_T_51[287:0] : _GEN_657; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1708 = 10'h82 == _T_9 ? _ram_T_51[287:0] : _GEN_658; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1709 = 10'h83 == _T_9 ? _ram_T_51[287:0] : _GEN_659; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1710 = 10'h84 == _T_9 ? _ram_T_51[287:0] : _GEN_660; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1711 = 10'h85 == _T_9 ? _ram_T_51[287:0] : _GEN_661; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1712 = 10'h86 == _T_9 ? _ram_T_51[287:0] : _GEN_662; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1713 = 10'h87 == _T_9 ? _ram_T_51[287:0] : _GEN_663; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1714 = 10'h88 == _T_9 ? _ram_T_51[287:0] : _GEN_664; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1715 = 10'h89 == _T_9 ? _ram_T_51[287:0] : _GEN_665; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1716 = 10'h8a == _T_9 ? _ram_T_51[287:0] : _GEN_666; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1717 = 10'h8b == _T_9 ? _ram_T_51[287:0] : _GEN_667; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1718 = 10'h8c == _T_9 ? _ram_T_51[287:0] : _GEN_668; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1719 = 10'h8d == _T_9 ? _ram_T_51[287:0] : _GEN_669; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1720 = 10'h8e == _T_9 ? _ram_T_51[287:0] : _GEN_670; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1721 = 10'h8f == _T_9 ? _ram_T_51[287:0] : _GEN_671; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1722 = 10'h90 == _T_9 ? _ram_T_51[287:0] : _GEN_672; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1723 = 10'h91 == _T_9 ? _ram_T_51[287:0] : _GEN_673; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1724 = 10'h92 == _T_9 ? _ram_T_51[287:0] : _GEN_674; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1725 = 10'h93 == _T_9 ? _ram_T_51[287:0] : _GEN_675; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1726 = 10'h94 == _T_9 ? _ram_T_51[287:0] : _GEN_676; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1727 = 10'h95 == _T_9 ? _ram_T_51[287:0] : _GEN_677; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1728 = 10'h96 == _T_9 ? _ram_T_51[287:0] : _GEN_678; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1729 = 10'h97 == _T_9 ? _ram_T_51[287:0] : _GEN_679; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1730 = 10'h98 == _T_9 ? _ram_T_51[287:0] : _GEN_680; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1731 = 10'h99 == _T_9 ? _ram_T_51[287:0] : _GEN_681; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1732 = 10'h9a == _T_9 ? _ram_T_51[287:0] : _GEN_682; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1733 = 10'h9b == _T_9 ? _ram_T_51[287:0] : _GEN_683; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1734 = 10'h9c == _T_9 ? _ram_T_51[287:0] : _GEN_684; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1735 = 10'h9d == _T_9 ? _ram_T_51[287:0] : _GEN_685; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1736 = 10'h9e == _T_9 ? _ram_T_51[287:0] : _GEN_686; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1737 = 10'h9f == _T_9 ? _ram_T_51[287:0] : _GEN_687; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1738 = 10'ha0 == _T_9 ? _ram_T_51[287:0] : _GEN_688; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1739 = 10'ha1 == _T_9 ? _ram_T_51[287:0] : _GEN_689; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1740 = 10'ha2 == _T_9 ? _ram_T_51[287:0] : _GEN_690; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1741 = 10'ha3 == _T_9 ? _ram_T_51[287:0] : _GEN_691; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1742 = 10'ha4 == _T_9 ? _ram_T_51[287:0] : _GEN_692; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1743 = 10'ha5 == _T_9 ? _ram_T_51[287:0] : _GEN_693; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1744 = 10'ha6 == _T_9 ? _ram_T_51[287:0] : _GEN_694; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1745 = 10'ha7 == _T_9 ? _ram_T_51[287:0] : _GEN_695; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1746 = 10'ha8 == _T_9 ? _ram_T_51[287:0] : _GEN_696; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1747 = 10'ha9 == _T_9 ? _ram_T_51[287:0] : _GEN_697; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1748 = 10'haa == _T_9 ? _ram_T_51[287:0] : _GEN_698; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1749 = 10'hab == _T_9 ? _ram_T_51[287:0] : _GEN_699; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1750 = 10'hac == _T_9 ? _ram_T_51[287:0] : _GEN_700; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1751 = 10'had == _T_9 ? _ram_T_51[287:0] : _GEN_701; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1752 = 10'hae == _T_9 ? _ram_T_51[287:0] : _GEN_702; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1753 = 10'haf == _T_9 ? _ram_T_51[287:0] : _GEN_703; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1754 = 10'hb0 == _T_9 ? _ram_T_51[287:0] : _GEN_704; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1755 = 10'hb1 == _T_9 ? _ram_T_51[287:0] : _GEN_705; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1756 = 10'hb2 == _T_9 ? _ram_T_51[287:0] : _GEN_706; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1757 = 10'hb3 == _T_9 ? _ram_T_51[287:0] : _GEN_707; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1758 = 10'hb4 == _T_9 ? _ram_T_51[287:0] : _GEN_708; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1759 = 10'hb5 == _T_9 ? _ram_T_51[287:0] : _GEN_709; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1760 = 10'hb6 == _T_9 ? _ram_T_51[287:0] : _GEN_710; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1761 = 10'hb7 == _T_9 ? _ram_T_51[287:0] : _GEN_711; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1762 = 10'hb8 == _T_9 ? _ram_T_51[287:0] : _GEN_712; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1763 = 10'hb9 == _T_9 ? _ram_T_51[287:0] : _GEN_713; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1764 = 10'hba == _T_9 ? _ram_T_51[287:0] : _GEN_714; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1765 = 10'hbb == _T_9 ? _ram_T_51[287:0] : _GEN_715; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1766 = 10'hbc == _T_9 ? _ram_T_51[287:0] : _GEN_716; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1767 = 10'hbd == _T_9 ? _ram_T_51[287:0] : _GEN_717; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1768 = 10'hbe == _T_9 ? _ram_T_51[287:0] : _GEN_718; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1769 = 10'hbf == _T_9 ? _ram_T_51[287:0] : _GEN_719; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1770 = 10'hc0 == _T_9 ? _ram_T_51[287:0] : _GEN_720; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1771 = 10'hc1 == _T_9 ? _ram_T_51[287:0] : _GEN_721; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1772 = 10'hc2 == _T_9 ? _ram_T_51[287:0] : _GEN_722; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1773 = 10'hc3 == _T_9 ? _ram_T_51[287:0] : _GEN_723; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1774 = 10'hc4 == _T_9 ? _ram_T_51[287:0] : _GEN_724; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1775 = 10'hc5 == _T_9 ? _ram_T_51[287:0] : _GEN_725; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1776 = 10'hc6 == _T_9 ? _ram_T_51[287:0] : _GEN_726; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1777 = 10'hc7 == _T_9 ? _ram_T_51[287:0] : _GEN_727; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1778 = 10'hc8 == _T_9 ? _ram_T_51[287:0] : _GEN_728; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1779 = 10'hc9 == _T_9 ? _ram_T_51[287:0] : _GEN_729; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1780 = 10'hca == _T_9 ? _ram_T_51[287:0] : _GEN_730; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1781 = 10'hcb == _T_9 ? _ram_T_51[287:0] : _GEN_731; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1782 = 10'hcc == _T_9 ? _ram_T_51[287:0] : _GEN_732; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1783 = 10'hcd == _T_9 ? _ram_T_51[287:0] : _GEN_733; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1784 = 10'hce == _T_9 ? _ram_T_51[287:0] : _GEN_734; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1785 = 10'hcf == _T_9 ? _ram_T_51[287:0] : _GEN_735; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1786 = 10'hd0 == _T_9 ? _ram_T_51[287:0] : _GEN_736; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1787 = 10'hd1 == _T_9 ? _ram_T_51[287:0] : _GEN_737; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1788 = 10'hd2 == _T_9 ? _ram_T_51[287:0] : _GEN_738; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1789 = 10'hd3 == _T_9 ? _ram_T_51[287:0] : _GEN_739; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1790 = 10'hd4 == _T_9 ? _ram_T_51[287:0] : _GEN_740; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1791 = 10'hd5 == _T_9 ? _ram_T_51[287:0] : _GEN_741; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1792 = 10'hd6 == _T_9 ? _ram_T_51[287:0] : _GEN_742; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1793 = 10'hd7 == _T_9 ? _ram_T_51[287:0] : _GEN_743; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1794 = 10'hd8 == _T_9 ? _ram_T_51[287:0] : _GEN_744; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1795 = 10'hd9 == _T_9 ? _ram_T_51[287:0] : _GEN_745; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1796 = 10'hda == _T_9 ? _ram_T_51[287:0] : _GEN_746; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1797 = 10'hdb == _T_9 ? _ram_T_51[287:0] : _GEN_747; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1798 = 10'hdc == _T_9 ? _ram_T_51[287:0] : _GEN_748; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1799 = 10'hdd == _T_9 ? _ram_T_51[287:0] : _GEN_749; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1800 = 10'hde == _T_9 ? _ram_T_51[287:0] : _GEN_750; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1801 = 10'hdf == _T_9 ? _ram_T_51[287:0] : _GEN_751; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1802 = 10'he0 == _T_9 ? _ram_T_51[287:0] : _GEN_752; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1803 = 10'he1 == _T_9 ? _ram_T_51[287:0] : _GEN_753; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1804 = 10'he2 == _T_9 ? _ram_T_51[287:0] : _GEN_754; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1805 = 10'he3 == _T_9 ? _ram_T_51[287:0] : _GEN_755; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1806 = 10'he4 == _T_9 ? _ram_T_51[287:0] : _GEN_756; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1807 = 10'he5 == _T_9 ? _ram_T_51[287:0] : _GEN_757; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1808 = 10'he6 == _T_9 ? _ram_T_51[287:0] : _GEN_758; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1809 = 10'he7 == _T_9 ? _ram_T_51[287:0] : _GEN_759; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1810 = 10'he8 == _T_9 ? _ram_T_51[287:0] : _GEN_760; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1811 = 10'he9 == _T_9 ? _ram_T_51[287:0] : _GEN_761; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1812 = 10'hea == _T_9 ? _ram_T_51[287:0] : _GEN_762; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1813 = 10'heb == _T_9 ? _ram_T_51[287:0] : _GEN_763; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1814 = 10'hec == _T_9 ? _ram_T_51[287:0] : _GEN_764; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1815 = 10'hed == _T_9 ? _ram_T_51[287:0] : _GEN_765; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1816 = 10'hee == _T_9 ? _ram_T_51[287:0] : _GEN_766; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1817 = 10'hef == _T_9 ? _ram_T_51[287:0] : _GEN_767; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1818 = 10'hf0 == _T_9 ? _ram_T_51[287:0] : _GEN_768; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1819 = 10'hf1 == _T_9 ? _ram_T_51[287:0] : _GEN_769; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1820 = 10'hf2 == _T_9 ? _ram_T_51[287:0] : _GEN_770; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1821 = 10'hf3 == _T_9 ? _ram_T_51[287:0] : _GEN_771; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1822 = 10'hf4 == _T_9 ? _ram_T_51[287:0] : _GEN_772; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1823 = 10'hf5 == _T_9 ? _ram_T_51[287:0] : _GEN_773; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1824 = 10'hf6 == _T_9 ? _ram_T_51[287:0] : _GEN_774; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1825 = 10'hf7 == _T_9 ? _ram_T_51[287:0] : _GEN_775; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1826 = 10'hf8 == _T_9 ? _ram_T_51[287:0] : _GEN_776; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1827 = 10'hf9 == _T_9 ? _ram_T_51[287:0] : _GEN_777; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1828 = 10'hfa == _T_9 ? _ram_T_51[287:0] : _GEN_778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1829 = 10'hfb == _T_9 ? _ram_T_51[287:0] : _GEN_779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1830 = 10'hfc == _T_9 ? _ram_T_51[287:0] : _GEN_780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1831 = 10'hfd == _T_9 ? _ram_T_51[287:0] : _GEN_781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1832 = 10'hfe == _T_9 ? _ram_T_51[287:0] : _GEN_782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1833 = 10'hff == _T_9 ? _ram_T_51[287:0] : _GEN_783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1834 = 10'h100 == _T_9 ? _ram_T_51[287:0] : _GEN_784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1835 = 10'h101 == _T_9 ? _ram_T_51[287:0] : _GEN_785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1836 = 10'h102 == _T_9 ? _ram_T_51[287:0] : _GEN_786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1837 = 10'h103 == _T_9 ? _ram_T_51[287:0] : _GEN_787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1838 = 10'h104 == _T_9 ? _ram_T_51[287:0] : _GEN_788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1839 = 10'h105 == _T_9 ? _ram_T_51[287:0] : _GEN_789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1840 = 10'h106 == _T_9 ? _ram_T_51[287:0] : _GEN_790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1841 = 10'h107 == _T_9 ? _ram_T_51[287:0] : _GEN_791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1842 = 10'h108 == _T_9 ? _ram_T_51[287:0] : _GEN_792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1843 = 10'h109 == _T_9 ? _ram_T_51[287:0] : _GEN_793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1844 = 10'h10a == _T_9 ? _ram_T_51[287:0] : _GEN_794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1845 = 10'h10b == _T_9 ? _ram_T_51[287:0] : _GEN_795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1846 = 10'h10c == _T_9 ? _ram_T_51[287:0] : _GEN_796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1847 = 10'h10d == _T_9 ? _ram_T_51[287:0] : _GEN_797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1848 = 10'h10e == _T_9 ? _ram_T_51[287:0] : _GEN_798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1849 = 10'h10f == _T_9 ? _ram_T_51[287:0] : _GEN_799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1850 = 10'h110 == _T_9 ? _ram_T_51[287:0] : _GEN_800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1851 = 10'h111 == _T_9 ? _ram_T_51[287:0] : _GEN_801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1852 = 10'h112 == _T_9 ? _ram_T_51[287:0] : _GEN_802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1853 = 10'h113 == _T_9 ? _ram_T_51[287:0] : _GEN_803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1854 = 10'h114 == _T_9 ? _ram_T_51[287:0] : _GEN_804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1855 = 10'h115 == _T_9 ? _ram_T_51[287:0] : _GEN_805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1856 = 10'h116 == _T_9 ? _ram_T_51[287:0] : _GEN_806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1857 = 10'h117 == _T_9 ? _ram_T_51[287:0] : _GEN_807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1858 = 10'h118 == _T_9 ? _ram_T_51[287:0] : _GEN_808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1859 = 10'h119 == _T_9 ? _ram_T_51[287:0] : _GEN_809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1860 = 10'h11a == _T_9 ? _ram_T_51[287:0] : _GEN_810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1861 = 10'h11b == _T_9 ? _ram_T_51[287:0] : _GEN_811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1862 = 10'h11c == _T_9 ? _ram_T_51[287:0] : _GEN_812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1863 = 10'h11d == _T_9 ? _ram_T_51[287:0] : _GEN_813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1864 = 10'h11e == _T_9 ? _ram_T_51[287:0] : _GEN_814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1865 = 10'h11f == _T_9 ? _ram_T_51[287:0] : _GEN_815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1866 = 10'h120 == _T_9 ? _ram_T_51[287:0] : _GEN_816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1867 = 10'h121 == _T_9 ? _ram_T_51[287:0] : _GEN_817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1868 = 10'h122 == _T_9 ? _ram_T_51[287:0] : _GEN_818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1869 = 10'h123 == _T_9 ? _ram_T_51[287:0] : _GEN_819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1870 = 10'h124 == _T_9 ? _ram_T_51[287:0] : _GEN_820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1871 = 10'h125 == _T_9 ? _ram_T_51[287:0] : _GEN_821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1872 = 10'h126 == _T_9 ? _ram_T_51[287:0] : _GEN_822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1873 = 10'h127 == _T_9 ? _ram_T_51[287:0] : _GEN_823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1874 = 10'h128 == _T_9 ? _ram_T_51[287:0] : _GEN_824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1875 = 10'h129 == _T_9 ? _ram_T_51[287:0] : _GEN_825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1876 = 10'h12a == _T_9 ? _ram_T_51[287:0] : _GEN_826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1877 = 10'h12b == _T_9 ? _ram_T_51[287:0] : _GEN_827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1878 = 10'h12c == _T_9 ? _ram_T_51[287:0] : _GEN_828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1879 = 10'h12d == _T_9 ? _ram_T_51[287:0] : _GEN_829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1880 = 10'h12e == _T_9 ? _ram_T_51[287:0] : _GEN_830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1881 = 10'h12f == _T_9 ? _ram_T_51[287:0] : _GEN_831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1882 = 10'h130 == _T_9 ? _ram_T_51[287:0] : _GEN_832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1883 = 10'h131 == _T_9 ? _ram_T_51[287:0] : _GEN_833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1884 = 10'h132 == _T_9 ? _ram_T_51[287:0] : _GEN_834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1885 = 10'h133 == _T_9 ? _ram_T_51[287:0] : _GEN_835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1886 = 10'h134 == _T_9 ? _ram_T_51[287:0] : _GEN_836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1887 = 10'h135 == _T_9 ? _ram_T_51[287:0] : _GEN_837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1888 = 10'h136 == _T_9 ? _ram_T_51[287:0] : _GEN_838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1889 = 10'h137 == _T_9 ? _ram_T_51[287:0] : _GEN_839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1890 = 10'h138 == _T_9 ? _ram_T_51[287:0] : _GEN_840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1891 = 10'h139 == _T_9 ? _ram_T_51[287:0] : _GEN_841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1892 = 10'h13a == _T_9 ? _ram_T_51[287:0] : _GEN_842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1893 = 10'h13b == _T_9 ? _ram_T_51[287:0] : _GEN_843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1894 = 10'h13c == _T_9 ? _ram_T_51[287:0] : _GEN_844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1895 = 10'h13d == _T_9 ? _ram_T_51[287:0] : _GEN_845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1896 = 10'h13e == _T_9 ? _ram_T_51[287:0] : _GEN_846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1897 = 10'h13f == _T_9 ? _ram_T_51[287:0] : _GEN_847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1898 = 10'h140 == _T_9 ? _ram_T_51[287:0] : _GEN_848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1899 = 10'h141 == _T_9 ? _ram_T_51[287:0] : _GEN_849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1900 = 10'h142 == _T_9 ? _ram_T_51[287:0] : _GEN_850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1901 = 10'h143 == _T_9 ? _ram_T_51[287:0] : _GEN_851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1902 = 10'h144 == _T_9 ? _ram_T_51[287:0] : _GEN_852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1903 = 10'h145 == _T_9 ? _ram_T_51[287:0] : _GEN_853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1904 = 10'h146 == _T_9 ? _ram_T_51[287:0] : _GEN_854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1905 = 10'h147 == _T_9 ? _ram_T_51[287:0] : _GEN_855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1906 = 10'h148 == _T_9 ? _ram_T_51[287:0] : _GEN_856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1907 = 10'h149 == _T_9 ? _ram_T_51[287:0] : _GEN_857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1908 = 10'h14a == _T_9 ? _ram_T_51[287:0] : _GEN_858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1909 = 10'h14b == _T_9 ? _ram_T_51[287:0] : _GEN_859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1910 = 10'h14c == _T_9 ? _ram_T_51[287:0] : _GEN_860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1911 = 10'h14d == _T_9 ? _ram_T_51[287:0] : _GEN_861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1912 = 10'h14e == _T_9 ? _ram_T_51[287:0] : _GEN_862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1913 = 10'h14f == _T_9 ? _ram_T_51[287:0] : _GEN_863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1914 = 10'h150 == _T_9 ? _ram_T_51[287:0] : _GEN_864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1915 = 10'h151 == _T_9 ? _ram_T_51[287:0] : _GEN_865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1916 = 10'h152 == _T_9 ? _ram_T_51[287:0] : _GEN_866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1917 = 10'h153 == _T_9 ? _ram_T_51[287:0] : _GEN_867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1918 = 10'h154 == _T_9 ? _ram_T_51[287:0] : _GEN_868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1919 = 10'h155 == _T_9 ? _ram_T_51[287:0] : _GEN_869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1920 = 10'h156 == _T_9 ? _ram_T_51[287:0] : _GEN_870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1921 = 10'h157 == _T_9 ? _ram_T_51[287:0] : _GEN_871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1922 = 10'h158 == _T_9 ? _ram_T_51[287:0] : _GEN_872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1923 = 10'h159 == _T_9 ? _ram_T_51[287:0] : _GEN_873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1924 = 10'h15a == _T_9 ? _ram_T_51[287:0] : _GEN_874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1925 = 10'h15b == _T_9 ? _ram_T_51[287:0] : _GEN_875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1926 = 10'h15c == _T_9 ? _ram_T_51[287:0] : _GEN_876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1927 = 10'h15d == _T_9 ? _ram_T_51[287:0] : _GEN_877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1928 = 10'h15e == _T_9 ? _ram_T_51[287:0] : _GEN_878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1929 = 10'h15f == _T_9 ? _ram_T_51[287:0] : _GEN_879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1930 = 10'h160 == _T_9 ? _ram_T_51[287:0] : _GEN_880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1931 = 10'h161 == _T_9 ? _ram_T_51[287:0] : _GEN_881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1932 = 10'h162 == _T_9 ? _ram_T_51[287:0] : _GEN_882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1933 = 10'h163 == _T_9 ? _ram_T_51[287:0] : _GEN_883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1934 = 10'h164 == _T_9 ? _ram_T_51[287:0] : _GEN_884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1935 = 10'h165 == _T_9 ? _ram_T_51[287:0] : _GEN_885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1936 = 10'h166 == _T_9 ? _ram_T_51[287:0] : _GEN_886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1937 = 10'h167 == _T_9 ? _ram_T_51[287:0] : _GEN_887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1938 = 10'h168 == _T_9 ? _ram_T_51[287:0] : _GEN_888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1939 = 10'h169 == _T_9 ? _ram_T_51[287:0] : _GEN_889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1940 = 10'h16a == _T_9 ? _ram_T_51[287:0] : _GEN_890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1941 = 10'h16b == _T_9 ? _ram_T_51[287:0] : _GEN_891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1942 = 10'h16c == _T_9 ? _ram_T_51[287:0] : _GEN_892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1943 = 10'h16d == _T_9 ? _ram_T_51[287:0] : _GEN_893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1944 = 10'h16e == _T_9 ? _ram_T_51[287:0] : _GEN_894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1945 = 10'h16f == _T_9 ? _ram_T_51[287:0] : _GEN_895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1946 = 10'h170 == _T_9 ? _ram_T_51[287:0] : _GEN_896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1947 = 10'h171 == _T_9 ? _ram_T_51[287:0] : _GEN_897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1948 = 10'h172 == _T_9 ? _ram_T_51[287:0] : _GEN_898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1949 = 10'h173 == _T_9 ? _ram_T_51[287:0] : _GEN_899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1950 = 10'h174 == _T_9 ? _ram_T_51[287:0] : _GEN_900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1951 = 10'h175 == _T_9 ? _ram_T_51[287:0] : _GEN_901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1952 = 10'h176 == _T_9 ? _ram_T_51[287:0] : _GEN_902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1953 = 10'h177 == _T_9 ? _ram_T_51[287:0] : _GEN_903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1954 = 10'h178 == _T_9 ? _ram_T_51[287:0] : _GEN_904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1955 = 10'h179 == _T_9 ? _ram_T_51[287:0] : _GEN_905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1956 = 10'h17a == _T_9 ? _ram_T_51[287:0] : _GEN_906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1957 = 10'h17b == _T_9 ? _ram_T_51[287:0] : _GEN_907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1958 = 10'h17c == _T_9 ? _ram_T_51[287:0] : _GEN_908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1959 = 10'h17d == _T_9 ? _ram_T_51[287:0] : _GEN_909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1960 = 10'h17e == _T_9 ? _ram_T_51[287:0] : _GEN_910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1961 = 10'h17f == _T_9 ? _ram_T_51[287:0] : _GEN_911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1962 = 10'h180 == _T_9 ? _ram_T_51[287:0] : _GEN_912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1963 = 10'h181 == _T_9 ? _ram_T_51[287:0] : _GEN_913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1964 = 10'h182 == _T_9 ? _ram_T_51[287:0] : _GEN_914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1965 = 10'h183 == _T_9 ? _ram_T_51[287:0] : _GEN_915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1966 = 10'h184 == _T_9 ? _ram_T_51[287:0] : _GEN_916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1967 = 10'h185 == _T_9 ? _ram_T_51[287:0] : _GEN_917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1968 = 10'h186 == _T_9 ? _ram_T_51[287:0] : _GEN_918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1969 = 10'h187 == _T_9 ? _ram_T_51[287:0] : _GEN_919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1970 = 10'h188 == _T_9 ? _ram_T_51[287:0] : _GEN_920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1971 = 10'h189 == _T_9 ? _ram_T_51[287:0] : _GEN_921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1972 = 10'h18a == _T_9 ? _ram_T_51[287:0] : _GEN_922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1973 = 10'h18b == _T_9 ? _ram_T_51[287:0] : _GEN_923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1974 = 10'h18c == _T_9 ? _ram_T_51[287:0] : _GEN_924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1975 = 10'h18d == _T_9 ? _ram_T_51[287:0] : _GEN_925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1976 = 10'h18e == _T_9 ? _ram_T_51[287:0] : _GEN_926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1977 = 10'h18f == _T_9 ? _ram_T_51[287:0] : _GEN_927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1978 = 10'h190 == _T_9 ? _ram_T_51[287:0] : _GEN_928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1979 = 10'h191 == _T_9 ? _ram_T_51[287:0] : _GEN_929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1980 = 10'h192 == _T_9 ? _ram_T_51[287:0] : _GEN_930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1981 = 10'h193 == _T_9 ? _ram_T_51[287:0] : _GEN_931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1982 = 10'h194 == _T_9 ? _ram_T_51[287:0] : _GEN_932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1983 = 10'h195 == _T_9 ? _ram_T_51[287:0] : _GEN_933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1984 = 10'h196 == _T_9 ? _ram_T_51[287:0] : _GEN_934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1985 = 10'h197 == _T_9 ? _ram_T_51[287:0] : _GEN_935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1986 = 10'h198 == _T_9 ? _ram_T_51[287:0] : _GEN_936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1987 = 10'h199 == _T_9 ? _ram_T_51[287:0] : _GEN_937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1988 = 10'h19a == _T_9 ? _ram_T_51[287:0] : _GEN_938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1989 = 10'h19b == _T_9 ? _ram_T_51[287:0] : _GEN_939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1990 = 10'h19c == _T_9 ? _ram_T_51[287:0] : _GEN_940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1991 = 10'h19d == _T_9 ? _ram_T_51[287:0] : _GEN_941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1992 = 10'h19e == _T_9 ? _ram_T_51[287:0] : _GEN_942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1993 = 10'h19f == _T_9 ? _ram_T_51[287:0] : _GEN_943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1994 = 10'h1a0 == _T_9 ? _ram_T_51[287:0] : _GEN_944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1995 = 10'h1a1 == _T_9 ? _ram_T_51[287:0] : _GEN_945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1996 = 10'h1a2 == _T_9 ? _ram_T_51[287:0] : _GEN_946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1997 = 10'h1a3 == _T_9 ? _ram_T_51[287:0] : _GEN_947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1998 = 10'h1a4 == _T_9 ? _ram_T_51[287:0] : _GEN_948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_1999 = 10'h1a5 == _T_9 ? _ram_T_51[287:0] : _GEN_949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2000 = 10'h1a6 == _T_9 ? _ram_T_51[287:0] : _GEN_950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2001 = 10'h1a7 == _T_9 ? _ram_T_51[287:0] : _GEN_951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2002 = 10'h1a8 == _T_9 ? _ram_T_51[287:0] : _GEN_952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2003 = 10'h1a9 == _T_9 ? _ram_T_51[287:0] : _GEN_953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2004 = 10'h1aa == _T_9 ? _ram_T_51[287:0] : _GEN_954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2005 = 10'h1ab == _T_9 ? _ram_T_51[287:0] : _GEN_955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2006 = 10'h1ac == _T_9 ? _ram_T_51[287:0] : _GEN_956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2007 = 10'h1ad == _T_9 ? _ram_T_51[287:0] : _GEN_957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2008 = 10'h1ae == _T_9 ? _ram_T_51[287:0] : _GEN_958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2009 = 10'h1af == _T_9 ? _ram_T_51[287:0] : _GEN_959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2010 = 10'h1b0 == _T_9 ? _ram_T_51[287:0] : _GEN_960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2011 = 10'h1b1 == _T_9 ? _ram_T_51[287:0] : _GEN_961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2012 = 10'h1b2 == _T_9 ? _ram_T_51[287:0] : _GEN_962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2013 = 10'h1b3 == _T_9 ? _ram_T_51[287:0] : _GEN_963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2014 = 10'h1b4 == _T_9 ? _ram_T_51[287:0] : _GEN_964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2015 = 10'h1b5 == _T_9 ? _ram_T_51[287:0] : _GEN_965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2016 = 10'h1b6 == _T_9 ? _ram_T_51[287:0] : _GEN_966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2017 = 10'h1b7 == _T_9 ? _ram_T_51[287:0] : _GEN_967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2018 = 10'h1b8 == _T_9 ? _ram_T_51[287:0] : _GEN_968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2019 = 10'h1b9 == _T_9 ? _ram_T_51[287:0] : _GEN_969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2020 = 10'h1ba == _T_9 ? _ram_T_51[287:0] : _GEN_970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2021 = 10'h1bb == _T_9 ? _ram_T_51[287:0] : _GEN_971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2022 = 10'h1bc == _T_9 ? _ram_T_51[287:0] : _GEN_972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2023 = 10'h1bd == _T_9 ? _ram_T_51[287:0] : _GEN_973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2024 = 10'h1be == _T_9 ? _ram_T_51[287:0] : _GEN_974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2025 = 10'h1bf == _T_9 ? _ram_T_51[287:0] : _GEN_975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2026 = 10'h1c0 == _T_9 ? _ram_T_51[287:0] : _GEN_976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2027 = 10'h1c1 == _T_9 ? _ram_T_51[287:0] : _GEN_977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2028 = 10'h1c2 == _T_9 ? _ram_T_51[287:0] : _GEN_978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2029 = 10'h1c3 == _T_9 ? _ram_T_51[287:0] : _GEN_979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2030 = 10'h1c4 == _T_9 ? _ram_T_51[287:0] : _GEN_980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2031 = 10'h1c5 == _T_9 ? _ram_T_51[287:0] : _GEN_981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2032 = 10'h1c6 == _T_9 ? _ram_T_51[287:0] : _GEN_982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2033 = 10'h1c7 == _T_9 ? _ram_T_51[287:0] : _GEN_983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2034 = 10'h1c8 == _T_9 ? _ram_T_51[287:0] : _GEN_984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2035 = 10'h1c9 == _T_9 ? _ram_T_51[287:0] : _GEN_985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2036 = 10'h1ca == _T_9 ? _ram_T_51[287:0] : _GEN_986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2037 = 10'h1cb == _T_9 ? _ram_T_51[287:0] : _GEN_987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2038 = 10'h1cc == _T_9 ? _ram_T_51[287:0] : _GEN_988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2039 = 10'h1cd == _T_9 ? _ram_T_51[287:0] : _GEN_989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2040 = 10'h1ce == _T_9 ? _ram_T_51[287:0] : _GEN_990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2041 = 10'h1cf == _T_9 ? _ram_T_51[287:0] : _GEN_991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2042 = 10'h1d0 == _T_9 ? _ram_T_51[287:0] : _GEN_992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2043 = 10'h1d1 == _T_9 ? _ram_T_51[287:0] : _GEN_993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2044 = 10'h1d2 == _T_9 ? _ram_T_51[287:0] : _GEN_994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2045 = 10'h1d3 == _T_9 ? _ram_T_51[287:0] : _GEN_995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2046 = 10'h1d4 == _T_9 ? _ram_T_51[287:0] : _GEN_996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2047 = 10'h1d5 == _T_9 ? _ram_T_51[287:0] : _GEN_997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2048 = 10'h1d6 == _T_9 ? _ram_T_51[287:0] : _GEN_998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2049 = 10'h1d7 == _T_9 ? _ram_T_51[287:0] : _GEN_999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2050 = 10'h1d8 == _T_9 ? _ram_T_51[287:0] : _GEN_1000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2051 = 10'h1d9 == _T_9 ? _ram_T_51[287:0] : _GEN_1001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2052 = 10'h1da == _T_9 ? _ram_T_51[287:0] : _GEN_1002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2053 = 10'h1db == _T_9 ? _ram_T_51[287:0] : _GEN_1003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2054 = 10'h1dc == _T_9 ? _ram_T_51[287:0] : _GEN_1004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2055 = 10'h1dd == _T_9 ? _ram_T_51[287:0] : _GEN_1005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2056 = 10'h1de == _T_9 ? _ram_T_51[287:0] : _GEN_1006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2057 = 10'h1df == _T_9 ? _ram_T_51[287:0] : _GEN_1007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2058 = 10'h1e0 == _T_9 ? _ram_T_51[287:0] : _GEN_1008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2059 = 10'h1e1 == _T_9 ? _ram_T_51[287:0] : _GEN_1009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2060 = 10'h1e2 == _T_9 ? _ram_T_51[287:0] : _GEN_1010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2061 = 10'h1e3 == _T_9 ? _ram_T_51[287:0] : _GEN_1011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2062 = 10'h1e4 == _T_9 ? _ram_T_51[287:0] : _GEN_1012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2063 = 10'h1e5 == _T_9 ? _ram_T_51[287:0] : _GEN_1013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2064 = 10'h1e6 == _T_9 ? _ram_T_51[287:0] : _GEN_1014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2065 = 10'h1e7 == _T_9 ? _ram_T_51[287:0] : _GEN_1015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2066 = 10'h1e8 == _T_9 ? _ram_T_51[287:0] : _GEN_1016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2067 = 10'h1e9 == _T_9 ? _ram_T_51[287:0] : _GEN_1017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2068 = 10'h1ea == _T_9 ? _ram_T_51[287:0] : _GEN_1018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2069 = 10'h1eb == _T_9 ? _ram_T_51[287:0] : _GEN_1019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2070 = 10'h1ec == _T_9 ? _ram_T_51[287:0] : _GEN_1020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2071 = 10'h1ed == _T_9 ? _ram_T_51[287:0] : _GEN_1021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2072 = 10'h1ee == _T_9 ? _ram_T_51[287:0] : _GEN_1022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2073 = 10'h1ef == _T_9 ? _ram_T_51[287:0] : _GEN_1023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2074 = 10'h1f0 == _T_9 ? _ram_T_51[287:0] : _GEN_1024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2075 = 10'h1f1 == _T_9 ? _ram_T_51[287:0] : _GEN_1025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2076 = 10'h1f2 == _T_9 ? _ram_T_51[287:0] : _GEN_1026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2077 = 10'h1f3 == _T_9 ? _ram_T_51[287:0] : _GEN_1027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2078 = 10'h1f4 == _T_9 ? _ram_T_51[287:0] : _GEN_1028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2079 = 10'h1f5 == _T_9 ? _ram_T_51[287:0] : _GEN_1029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2080 = 10'h1f6 == _T_9 ? _ram_T_51[287:0] : _GEN_1030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2081 = 10'h1f7 == _T_9 ? _ram_T_51[287:0] : _GEN_1031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2082 = 10'h1f8 == _T_9 ? _ram_T_51[287:0] : _GEN_1032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2083 = 10'h1f9 == _T_9 ? _ram_T_51[287:0] : _GEN_1033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2084 = 10'h1fa == _T_9 ? _ram_T_51[287:0] : _GEN_1034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2085 = 10'h1fb == _T_9 ? _ram_T_51[287:0] : _GEN_1035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2086 = 10'h1fc == _T_9 ? _ram_T_51[287:0] : _GEN_1036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2087 = 10'h1fd == _T_9 ? _ram_T_51[287:0] : _GEN_1037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2088 = 10'h1fe == _T_9 ? _ram_T_51[287:0] : _GEN_1038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2089 = 10'h1ff == _T_9 ? _ram_T_51[287:0] : _GEN_1039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2090 = 10'h200 == _T_9 ? _ram_T_51[287:0] : _GEN_1040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2091 = 10'h201 == _T_9 ? _ram_T_51[287:0] : _GEN_1041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2092 = 10'h202 == _T_9 ? _ram_T_51[287:0] : _GEN_1042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2093 = 10'h203 == _T_9 ? _ram_T_51[287:0] : _GEN_1043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2094 = 10'h204 == _T_9 ? _ram_T_51[287:0] : _GEN_1044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2095 = 10'h205 == _T_9 ? _ram_T_51[287:0] : _GEN_1045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2096 = 10'h206 == _T_9 ? _ram_T_51[287:0] : _GEN_1046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2097 = 10'h207 == _T_9 ? _ram_T_51[287:0] : _GEN_1047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2098 = 10'h208 == _T_9 ? _ram_T_51[287:0] : _GEN_1048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2099 = 10'h209 == _T_9 ? _ram_T_51[287:0] : _GEN_1049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2100 = 10'h20a == _T_9 ? _ram_T_51[287:0] : _GEN_1050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2101 = 10'h20b == _T_9 ? _ram_T_51[287:0] : _GEN_1051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2102 = 10'h20c == _T_9 ? _ram_T_51[287:0] : _GEN_1052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_11 = h + 10'h2; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_2 = vga_mem_ram_MPORT_18_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_2 = vga_mem_ram_MPORT_19_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_2 = vga_mem_ram_MPORT_20_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_2 = vga_mem_ram_MPORT_21_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_2 = vga_mem_ram_MPORT_22_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_2 = vga_mem_ram_MPORT_23_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_2 = vga_mem_ram_MPORT_24_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_2 = vga_mem_ram_MPORT_25_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_2 = vga_mem_ram_MPORT_26_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_72 = {278'h0,ram_hi_hi_hi_lo_2,ram_hi_hi_lo_2,ram_hi_lo_hi_2,ram_hi_lo_lo_2,ram_lo_hi_hi_hi_2,
    ram_lo_hi_hi_lo_2,ram_lo_hi_lo_2,ram_lo_lo_hi_2,ram_lo_lo_lo_2}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19064 = {{8191'd0}, _ram_T_72}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_76 = _GEN_19064 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_2104 = 10'h1 == _T_11 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2105 = 10'h2 == _T_11 ? ram_2 : _GEN_2104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2106 = 10'h3 == _T_11 ? ram_3 : _GEN_2105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2107 = 10'h4 == _T_11 ? ram_4 : _GEN_2106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2108 = 10'h5 == _T_11 ? ram_5 : _GEN_2107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2109 = 10'h6 == _T_11 ? ram_6 : _GEN_2108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2110 = 10'h7 == _T_11 ? ram_7 : _GEN_2109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2111 = 10'h8 == _T_11 ? ram_8 : _GEN_2110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2112 = 10'h9 == _T_11 ? ram_9 : _GEN_2111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2113 = 10'ha == _T_11 ? ram_10 : _GEN_2112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2114 = 10'hb == _T_11 ? ram_11 : _GEN_2113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2115 = 10'hc == _T_11 ? ram_12 : _GEN_2114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2116 = 10'hd == _T_11 ? ram_13 : _GEN_2115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2117 = 10'he == _T_11 ? ram_14 : _GEN_2116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2118 = 10'hf == _T_11 ? ram_15 : _GEN_2117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2119 = 10'h10 == _T_11 ? ram_16 : _GEN_2118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2120 = 10'h11 == _T_11 ? ram_17 : _GEN_2119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2121 = 10'h12 == _T_11 ? ram_18 : _GEN_2120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2122 = 10'h13 == _T_11 ? ram_19 : _GEN_2121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2123 = 10'h14 == _T_11 ? ram_20 : _GEN_2122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2124 = 10'h15 == _T_11 ? ram_21 : _GEN_2123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2125 = 10'h16 == _T_11 ? ram_22 : _GEN_2124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2126 = 10'h17 == _T_11 ? ram_23 : _GEN_2125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2127 = 10'h18 == _T_11 ? ram_24 : _GEN_2126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2128 = 10'h19 == _T_11 ? ram_25 : _GEN_2127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2129 = 10'h1a == _T_11 ? ram_26 : _GEN_2128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2130 = 10'h1b == _T_11 ? ram_27 : _GEN_2129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2131 = 10'h1c == _T_11 ? ram_28 : _GEN_2130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2132 = 10'h1d == _T_11 ? ram_29 : _GEN_2131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2133 = 10'h1e == _T_11 ? ram_30 : _GEN_2132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2134 = 10'h1f == _T_11 ? ram_31 : _GEN_2133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2135 = 10'h20 == _T_11 ? ram_32 : _GEN_2134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2136 = 10'h21 == _T_11 ? ram_33 : _GEN_2135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2137 = 10'h22 == _T_11 ? ram_34 : _GEN_2136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2138 = 10'h23 == _T_11 ? ram_35 : _GEN_2137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2139 = 10'h24 == _T_11 ? ram_36 : _GEN_2138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2140 = 10'h25 == _T_11 ? ram_37 : _GEN_2139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2141 = 10'h26 == _T_11 ? ram_38 : _GEN_2140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2142 = 10'h27 == _T_11 ? ram_39 : _GEN_2141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2143 = 10'h28 == _T_11 ? ram_40 : _GEN_2142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2144 = 10'h29 == _T_11 ? ram_41 : _GEN_2143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2145 = 10'h2a == _T_11 ? ram_42 : _GEN_2144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2146 = 10'h2b == _T_11 ? ram_43 : _GEN_2145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2147 = 10'h2c == _T_11 ? ram_44 : _GEN_2146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2148 = 10'h2d == _T_11 ? ram_45 : _GEN_2147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2149 = 10'h2e == _T_11 ? ram_46 : _GEN_2148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2150 = 10'h2f == _T_11 ? ram_47 : _GEN_2149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2151 = 10'h30 == _T_11 ? ram_48 : _GEN_2150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2152 = 10'h31 == _T_11 ? ram_49 : _GEN_2151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2153 = 10'h32 == _T_11 ? ram_50 : _GEN_2152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2154 = 10'h33 == _T_11 ? ram_51 : _GEN_2153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2155 = 10'h34 == _T_11 ? ram_52 : _GEN_2154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2156 = 10'h35 == _T_11 ? ram_53 : _GEN_2155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2157 = 10'h36 == _T_11 ? ram_54 : _GEN_2156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2158 = 10'h37 == _T_11 ? ram_55 : _GEN_2157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2159 = 10'h38 == _T_11 ? ram_56 : _GEN_2158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2160 = 10'h39 == _T_11 ? ram_57 : _GEN_2159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2161 = 10'h3a == _T_11 ? ram_58 : _GEN_2160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2162 = 10'h3b == _T_11 ? ram_59 : _GEN_2161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2163 = 10'h3c == _T_11 ? ram_60 : _GEN_2162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2164 = 10'h3d == _T_11 ? ram_61 : _GEN_2163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2165 = 10'h3e == _T_11 ? ram_62 : _GEN_2164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2166 = 10'h3f == _T_11 ? ram_63 : _GEN_2165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2167 = 10'h40 == _T_11 ? ram_64 : _GEN_2166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2168 = 10'h41 == _T_11 ? ram_65 : _GEN_2167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2169 = 10'h42 == _T_11 ? ram_66 : _GEN_2168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2170 = 10'h43 == _T_11 ? ram_67 : _GEN_2169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2171 = 10'h44 == _T_11 ? ram_68 : _GEN_2170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2172 = 10'h45 == _T_11 ? ram_69 : _GEN_2171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2173 = 10'h46 == _T_11 ? ram_70 : _GEN_2172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2174 = 10'h47 == _T_11 ? ram_71 : _GEN_2173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2175 = 10'h48 == _T_11 ? ram_72 : _GEN_2174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2176 = 10'h49 == _T_11 ? ram_73 : _GEN_2175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2177 = 10'h4a == _T_11 ? ram_74 : _GEN_2176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2178 = 10'h4b == _T_11 ? ram_75 : _GEN_2177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2179 = 10'h4c == _T_11 ? ram_76 : _GEN_2178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2180 = 10'h4d == _T_11 ? ram_77 : _GEN_2179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2181 = 10'h4e == _T_11 ? ram_78 : _GEN_2180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2182 = 10'h4f == _T_11 ? ram_79 : _GEN_2181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2183 = 10'h50 == _T_11 ? ram_80 : _GEN_2182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2184 = 10'h51 == _T_11 ? ram_81 : _GEN_2183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2185 = 10'h52 == _T_11 ? ram_82 : _GEN_2184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2186 = 10'h53 == _T_11 ? ram_83 : _GEN_2185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2187 = 10'h54 == _T_11 ? ram_84 : _GEN_2186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2188 = 10'h55 == _T_11 ? ram_85 : _GEN_2187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2189 = 10'h56 == _T_11 ? ram_86 : _GEN_2188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2190 = 10'h57 == _T_11 ? ram_87 : _GEN_2189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2191 = 10'h58 == _T_11 ? ram_88 : _GEN_2190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2192 = 10'h59 == _T_11 ? ram_89 : _GEN_2191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2193 = 10'h5a == _T_11 ? ram_90 : _GEN_2192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2194 = 10'h5b == _T_11 ? ram_91 : _GEN_2193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2195 = 10'h5c == _T_11 ? ram_92 : _GEN_2194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2196 = 10'h5d == _T_11 ? ram_93 : _GEN_2195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2197 = 10'h5e == _T_11 ? ram_94 : _GEN_2196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2198 = 10'h5f == _T_11 ? ram_95 : _GEN_2197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2199 = 10'h60 == _T_11 ? ram_96 : _GEN_2198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2200 = 10'h61 == _T_11 ? ram_97 : _GEN_2199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2201 = 10'h62 == _T_11 ? ram_98 : _GEN_2200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2202 = 10'h63 == _T_11 ? ram_99 : _GEN_2201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2203 = 10'h64 == _T_11 ? ram_100 : _GEN_2202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2204 = 10'h65 == _T_11 ? ram_101 : _GEN_2203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2205 = 10'h66 == _T_11 ? ram_102 : _GEN_2204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2206 = 10'h67 == _T_11 ? ram_103 : _GEN_2205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2207 = 10'h68 == _T_11 ? ram_104 : _GEN_2206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2208 = 10'h69 == _T_11 ? ram_105 : _GEN_2207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2209 = 10'h6a == _T_11 ? ram_106 : _GEN_2208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2210 = 10'h6b == _T_11 ? ram_107 : _GEN_2209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2211 = 10'h6c == _T_11 ? ram_108 : _GEN_2210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2212 = 10'h6d == _T_11 ? ram_109 : _GEN_2211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2213 = 10'h6e == _T_11 ? ram_110 : _GEN_2212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2214 = 10'h6f == _T_11 ? ram_111 : _GEN_2213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2215 = 10'h70 == _T_11 ? ram_112 : _GEN_2214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2216 = 10'h71 == _T_11 ? ram_113 : _GEN_2215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2217 = 10'h72 == _T_11 ? ram_114 : _GEN_2216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2218 = 10'h73 == _T_11 ? ram_115 : _GEN_2217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2219 = 10'h74 == _T_11 ? ram_116 : _GEN_2218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2220 = 10'h75 == _T_11 ? ram_117 : _GEN_2219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2221 = 10'h76 == _T_11 ? ram_118 : _GEN_2220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2222 = 10'h77 == _T_11 ? ram_119 : _GEN_2221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2223 = 10'h78 == _T_11 ? ram_120 : _GEN_2222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2224 = 10'h79 == _T_11 ? ram_121 : _GEN_2223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2225 = 10'h7a == _T_11 ? ram_122 : _GEN_2224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2226 = 10'h7b == _T_11 ? ram_123 : _GEN_2225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2227 = 10'h7c == _T_11 ? ram_124 : _GEN_2226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2228 = 10'h7d == _T_11 ? ram_125 : _GEN_2227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2229 = 10'h7e == _T_11 ? ram_126 : _GEN_2228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2230 = 10'h7f == _T_11 ? ram_127 : _GEN_2229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2231 = 10'h80 == _T_11 ? ram_128 : _GEN_2230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2232 = 10'h81 == _T_11 ? ram_129 : _GEN_2231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2233 = 10'h82 == _T_11 ? ram_130 : _GEN_2232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2234 = 10'h83 == _T_11 ? ram_131 : _GEN_2233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2235 = 10'h84 == _T_11 ? ram_132 : _GEN_2234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2236 = 10'h85 == _T_11 ? ram_133 : _GEN_2235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2237 = 10'h86 == _T_11 ? ram_134 : _GEN_2236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2238 = 10'h87 == _T_11 ? ram_135 : _GEN_2237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2239 = 10'h88 == _T_11 ? ram_136 : _GEN_2238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2240 = 10'h89 == _T_11 ? ram_137 : _GEN_2239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2241 = 10'h8a == _T_11 ? ram_138 : _GEN_2240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2242 = 10'h8b == _T_11 ? ram_139 : _GEN_2241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2243 = 10'h8c == _T_11 ? ram_140 : _GEN_2242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2244 = 10'h8d == _T_11 ? ram_141 : _GEN_2243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2245 = 10'h8e == _T_11 ? ram_142 : _GEN_2244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2246 = 10'h8f == _T_11 ? ram_143 : _GEN_2245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2247 = 10'h90 == _T_11 ? ram_144 : _GEN_2246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2248 = 10'h91 == _T_11 ? ram_145 : _GEN_2247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2249 = 10'h92 == _T_11 ? ram_146 : _GEN_2248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2250 = 10'h93 == _T_11 ? ram_147 : _GEN_2249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2251 = 10'h94 == _T_11 ? ram_148 : _GEN_2250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2252 = 10'h95 == _T_11 ? ram_149 : _GEN_2251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2253 = 10'h96 == _T_11 ? ram_150 : _GEN_2252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2254 = 10'h97 == _T_11 ? ram_151 : _GEN_2253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2255 = 10'h98 == _T_11 ? ram_152 : _GEN_2254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2256 = 10'h99 == _T_11 ? ram_153 : _GEN_2255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2257 = 10'h9a == _T_11 ? ram_154 : _GEN_2256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2258 = 10'h9b == _T_11 ? ram_155 : _GEN_2257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2259 = 10'h9c == _T_11 ? ram_156 : _GEN_2258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2260 = 10'h9d == _T_11 ? ram_157 : _GEN_2259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2261 = 10'h9e == _T_11 ? ram_158 : _GEN_2260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2262 = 10'h9f == _T_11 ? ram_159 : _GEN_2261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2263 = 10'ha0 == _T_11 ? ram_160 : _GEN_2262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2264 = 10'ha1 == _T_11 ? ram_161 : _GEN_2263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2265 = 10'ha2 == _T_11 ? ram_162 : _GEN_2264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2266 = 10'ha3 == _T_11 ? ram_163 : _GEN_2265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2267 = 10'ha4 == _T_11 ? ram_164 : _GEN_2266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2268 = 10'ha5 == _T_11 ? ram_165 : _GEN_2267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2269 = 10'ha6 == _T_11 ? ram_166 : _GEN_2268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2270 = 10'ha7 == _T_11 ? ram_167 : _GEN_2269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2271 = 10'ha8 == _T_11 ? ram_168 : _GEN_2270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2272 = 10'ha9 == _T_11 ? ram_169 : _GEN_2271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2273 = 10'haa == _T_11 ? ram_170 : _GEN_2272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2274 = 10'hab == _T_11 ? ram_171 : _GEN_2273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2275 = 10'hac == _T_11 ? ram_172 : _GEN_2274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2276 = 10'had == _T_11 ? ram_173 : _GEN_2275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2277 = 10'hae == _T_11 ? ram_174 : _GEN_2276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2278 = 10'haf == _T_11 ? ram_175 : _GEN_2277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2279 = 10'hb0 == _T_11 ? ram_176 : _GEN_2278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2280 = 10'hb1 == _T_11 ? ram_177 : _GEN_2279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2281 = 10'hb2 == _T_11 ? ram_178 : _GEN_2280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2282 = 10'hb3 == _T_11 ? ram_179 : _GEN_2281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2283 = 10'hb4 == _T_11 ? ram_180 : _GEN_2282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2284 = 10'hb5 == _T_11 ? ram_181 : _GEN_2283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2285 = 10'hb6 == _T_11 ? ram_182 : _GEN_2284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2286 = 10'hb7 == _T_11 ? ram_183 : _GEN_2285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2287 = 10'hb8 == _T_11 ? ram_184 : _GEN_2286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2288 = 10'hb9 == _T_11 ? ram_185 : _GEN_2287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2289 = 10'hba == _T_11 ? ram_186 : _GEN_2288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2290 = 10'hbb == _T_11 ? ram_187 : _GEN_2289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2291 = 10'hbc == _T_11 ? ram_188 : _GEN_2290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2292 = 10'hbd == _T_11 ? ram_189 : _GEN_2291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2293 = 10'hbe == _T_11 ? ram_190 : _GEN_2292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2294 = 10'hbf == _T_11 ? ram_191 : _GEN_2293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2295 = 10'hc0 == _T_11 ? ram_192 : _GEN_2294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2296 = 10'hc1 == _T_11 ? ram_193 : _GEN_2295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2297 = 10'hc2 == _T_11 ? ram_194 : _GEN_2296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2298 = 10'hc3 == _T_11 ? ram_195 : _GEN_2297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2299 = 10'hc4 == _T_11 ? ram_196 : _GEN_2298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2300 = 10'hc5 == _T_11 ? ram_197 : _GEN_2299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2301 = 10'hc6 == _T_11 ? ram_198 : _GEN_2300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2302 = 10'hc7 == _T_11 ? ram_199 : _GEN_2301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2303 = 10'hc8 == _T_11 ? ram_200 : _GEN_2302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2304 = 10'hc9 == _T_11 ? ram_201 : _GEN_2303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2305 = 10'hca == _T_11 ? ram_202 : _GEN_2304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2306 = 10'hcb == _T_11 ? ram_203 : _GEN_2305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2307 = 10'hcc == _T_11 ? ram_204 : _GEN_2306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2308 = 10'hcd == _T_11 ? ram_205 : _GEN_2307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2309 = 10'hce == _T_11 ? ram_206 : _GEN_2308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2310 = 10'hcf == _T_11 ? ram_207 : _GEN_2309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2311 = 10'hd0 == _T_11 ? ram_208 : _GEN_2310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2312 = 10'hd1 == _T_11 ? ram_209 : _GEN_2311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2313 = 10'hd2 == _T_11 ? ram_210 : _GEN_2312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2314 = 10'hd3 == _T_11 ? ram_211 : _GEN_2313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2315 = 10'hd4 == _T_11 ? ram_212 : _GEN_2314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2316 = 10'hd5 == _T_11 ? ram_213 : _GEN_2315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2317 = 10'hd6 == _T_11 ? ram_214 : _GEN_2316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2318 = 10'hd7 == _T_11 ? ram_215 : _GEN_2317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2319 = 10'hd8 == _T_11 ? ram_216 : _GEN_2318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2320 = 10'hd9 == _T_11 ? ram_217 : _GEN_2319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2321 = 10'hda == _T_11 ? ram_218 : _GEN_2320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2322 = 10'hdb == _T_11 ? ram_219 : _GEN_2321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2323 = 10'hdc == _T_11 ? ram_220 : _GEN_2322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2324 = 10'hdd == _T_11 ? ram_221 : _GEN_2323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2325 = 10'hde == _T_11 ? ram_222 : _GEN_2324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2326 = 10'hdf == _T_11 ? ram_223 : _GEN_2325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2327 = 10'he0 == _T_11 ? ram_224 : _GEN_2326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2328 = 10'he1 == _T_11 ? ram_225 : _GEN_2327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2329 = 10'he2 == _T_11 ? ram_226 : _GEN_2328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2330 = 10'he3 == _T_11 ? ram_227 : _GEN_2329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2331 = 10'he4 == _T_11 ? ram_228 : _GEN_2330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2332 = 10'he5 == _T_11 ? ram_229 : _GEN_2331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2333 = 10'he6 == _T_11 ? ram_230 : _GEN_2332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2334 = 10'he7 == _T_11 ? ram_231 : _GEN_2333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2335 = 10'he8 == _T_11 ? ram_232 : _GEN_2334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2336 = 10'he9 == _T_11 ? ram_233 : _GEN_2335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2337 = 10'hea == _T_11 ? ram_234 : _GEN_2336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2338 = 10'heb == _T_11 ? ram_235 : _GEN_2337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2339 = 10'hec == _T_11 ? ram_236 : _GEN_2338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2340 = 10'hed == _T_11 ? ram_237 : _GEN_2339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2341 = 10'hee == _T_11 ? ram_238 : _GEN_2340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2342 = 10'hef == _T_11 ? ram_239 : _GEN_2341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2343 = 10'hf0 == _T_11 ? ram_240 : _GEN_2342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2344 = 10'hf1 == _T_11 ? ram_241 : _GEN_2343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2345 = 10'hf2 == _T_11 ? ram_242 : _GEN_2344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2346 = 10'hf3 == _T_11 ? ram_243 : _GEN_2345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2347 = 10'hf4 == _T_11 ? ram_244 : _GEN_2346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2348 = 10'hf5 == _T_11 ? ram_245 : _GEN_2347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2349 = 10'hf6 == _T_11 ? ram_246 : _GEN_2348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2350 = 10'hf7 == _T_11 ? ram_247 : _GEN_2349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2351 = 10'hf8 == _T_11 ? ram_248 : _GEN_2350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2352 = 10'hf9 == _T_11 ? ram_249 : _GEN_2351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2353 = 10'hfa == _T_11 ? ram_250 : _GEN_2352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2354 = 10'hfb == _T_11 ? ram_251 : _GEN_2353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2355 = 10'hfc == _T_11 ? ram_252 : _GEN_2354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2356 = 10'hfd == _T_11 ? ram_253 : _GEN_2355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2357 = 10'hfe == _T_11 ? ram_254 : _GEN_2356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2358 = 10'hff == _T_11 ? ram_255 : _GEN_2357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2359 = 10'h100 == _T_11 ? ram_256 : _GEN_2358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2360 = 10'h101 == _T_11 ? ram_257 : _GEN_2359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2361 = 10'h102 == _T_11 ? ram_258 : _GEN_2360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2362 = 10'h103 == _T_11 ? ram_259 : _GEN_2361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2363 = 10'h104 == _T_11 ? ram_260 : _GEN_2362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2364 = 10'h105 == _T_11 ? ram_261 : _GEN_2363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2365 = 10'h106 == _T_11 ? ram_262 : _GEN_2364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2366 = 10'h107 == _T_11 ? ram_263 : _GEN_2365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2367 = 10'h108 == _T_11 ? ram_264 : _GEN_2366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2368 = 10'h109 == _T_11 ? ram_265 : _GEN_2367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2369 = 10'h10a == _T_11 ? ram_266 : _GEN_2368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2370 = 10'h10b == _T_11 ? ram_267 : _GEN_2369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2371 = 10'h10c == _T_11 ? ram_268 : _GEN_2370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2372 = 10'h10d == _T_11 ? ram_269 : _GEN_2371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2373 = 10'h10e == _T_11 ? ram_270 : _GEN_2372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2374 = 10'h10f == _T_11 ? ram_271 : _GEN_2373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2375 = 10'h110 == _T_11 ? ram_272 : _GEN_2374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2376 = 10'h111 == _T_11 ? ram_273 : _GEN_2375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2377 = 10'h112 == _T_11 ? ram_274 : _GEN_2376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2378 = 10'h113 == _T_11 ? ram_275 : _GEN_2377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2379 = 10'h114 == _T_11 ? ram_276 : _GEN_2378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2380 = 10'h115 == _T_11 ? ram_277 : _GEN_2379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2381 = 10'h116 == _T_11 ? ram_278 : _GEN_2380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2382 = 10'h117 == _T_11 ? ram_279 : _GEN_2381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2383 = 10'h118 == _T_11 ? ram_280 : _GEN_2382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2384 = 10'h119 == _T_11 ? ram_281 : _GEN_2383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2385 = 10'h11a == _T_11 ? ram_282 : _GEN_2384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2386 = 10'h11b == _T_11 ? ram_283 : _GEN_2385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2387 = 10'h11c == _T_11 ? ram_284 : _GEN_2386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2388 = 10'h11d == _T_11 ? ram_285 : _GEN_2387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2389 = 10'h11e == _T_11 ? ram_286 : _GEN_2388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2390 = 10'h11f == _T_11 ? ram_287 : _GEN_2389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2391 = 10'h120 == _T_11 ? ram_288 : _GEN_2390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2392 = 10'h121 == _T_11 ? ram_289 : _GEN_2391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2393 = 10'h122 == _T_11 ? ram_290 : _GEN_2392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2394 = 10'h123 == _T_11 ? ram_291 : _GEN_2393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2395 = 10'h124 == _T_11 ? ram_292 : _GEN_2394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2396 = 10'h125 == _T_11 ? ram_293 : _GEN_2395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2397 = 10'h126 == _T_11 ? ram_294 : _GEN_2396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2398 = 10'h127 == _T_11 ? ram_295 : _GEN_2397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2399 = 10'h128 == _T_11 ? ram_296 : _GEN_2398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2400 = 10'h129 == _T_11 ? ram_297 : _GEN_2399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2401 = 10'h12a == _T_11 ? ram_298 : _GEN_2400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2402 = 10'h12b == _T_11 ? ram_299 : _GEN_2401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2403 = 10'h12c == _T_11 ? ram_300 : _GEN_2402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2404 = 10'h12d == _T_11 ? ram_301 : _GEN_2403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2405 = 10'h12e == _T_11 ? ram_302 : _GEN_2404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2406 = 10'h12f == _T_11 ? ram_303 : _GEN_2405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2407 = 10'h130 == _T_11 ? ram_304 : _GEN_2406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2408 = 10'h131 == _T_11 ? ram_305 : _GEN_2407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2409 = 10'h132 == _T_11 ? ram_306 : _GEN_2408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2410 = 10'h133 == _T_11 ? ram_307 : _GEN_2409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2411 = 10'h134 == _T_11 ? ram_308 : _GEN_2410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2412 = 10'h135 == _T_11 ? ram_309 : _GEN_2411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2413 = 10'h136 == _T_11 ? ram_310 : _GEN_2412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2414 = 10'h137 == _T_11 ? ram_311 : _GEN_2413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2415 = 10'h138 == _T_11 ? ram_312 : _GEN_2414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2416 = 10'h139 == _T_11 ? ram_313 : _GEN_2415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2417 = 10'h13a == _T_11 ? ram_314 : _GEN_2416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2418 = 10'h13b == _T_11 ? ram_315 : _GEN_2417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2419 = 10'h13c == _T_11 ? ram_316 : _GEN_2418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2420 = 10'h13d == _T_11 ? ram_317 : _GEN_2419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2421 = 10'h13e == _T_11 ? ram_318 : _GEN_2420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2422 = 10'h13f == _T_11 ? ram_319 : _GEN_2421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2423 = 10'h140 == _T_11 ? ram_320 : _GEN_2422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2424 = 10'h141 == _T_11 ? ram_321 : _GEN_2423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2425 = 10'h142 == _T_11 ? ram_322 : _GEN_2424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2426 = 10'h143 == _T_11 ? ram_323 : _GEN_2425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2427 = 10'h144 == _T_11 ? ram_324 : _GEN_2426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2428 = 10'h145 == _T_11 ? ram_325 : _GEN_2427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2429 = 10'h146 == _T_11 ? ram_326 : _GEN_2428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2430 = 10'h147 == _T_11 ? ram_327 : _GEN_2429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2431 = 10'h148 == _T_11 ? ram_328 : _GEN_2430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2432 = 10'h149 == _T_11 ? ram_329 : _GEN_2431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2433 = 10'h14a == _T_11 ? ram_330 : _GEN_2432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2434 = 10'h14b == _T_11 ? ram_331 : _GEN_2433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2435 = 10'h14c == _T_11 ? ram_332 : _GEN_2434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2436 = 10'h14d == _T_11 ? ram_333 : _GEN_2435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2437 = 10'h14e == _T_11 ? ram_334 : _GEN_2436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2438 = 10'h14f == _T_11 ? ram_335 : _GEN_2437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2439 = 10'h150 == _T_11 ? ram_336 : _GEN_2438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2440 = 10'h151 == _T_11 ? ram_337 : _GEN_2439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2441 = 10'h152 == _T_11 ? ram_338 : _GEN_2440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2442 = 10'h153 == _T_11 ? ram_339 : _GEN_2441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2443 = 10'h154 == _T_11 ? ram_340 : _GEN_2442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2444 = 10'h155 == _T_11 ? ram_341 : _GEN_2443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2445 = 10'h156 == _T_11 ? ram_342 : _GEN_2444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2446 = 10'h157 == _T_11 ? ram_343 : _GEN_2445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2447 = 10'h158 == _T_11 ? ram_344 : _GEN_2446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2448 = 10'h159 == _T_11 ? ram_345 : _GEN_2447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2449 = 10'h15a == _T_11 ? ram_346 : _GEN_2448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2450 = 10'h15b == _T_11 ? ram_347 : _GEN_2449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2451 = 10'h15c == _T_11 ? ram_348 : _GEN_2450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2452 = 10'h15d == _T_11 ? ram_349 : _GEN_2451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2453 = 10'h15e == _T_11 ? ram_350 : _GEN_2452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2454 = 10'h15f == _T_11 ? ram_351 : _GEN_2453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2455 = 10'h160 == _T_11 ? ram_352 : _GEN_2454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2456 = 10'h161 == _T_11 ? ram_353 : _GEN_2455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2457 = 10'h162 == _T_11 ? ram_354 : _GEN_2456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2458 = 10'h163 == _T_11 ? ram_355 : _GEN_2457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2459 = 10'h164 == _T_11 ? ram_356 : _GEN_2458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2460 = 10'h165 == _T_11 ? ram_357 : _GEN_2459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2461 = 10'h166 == _T_11 ? ram_358 : _GEN_2460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2462 = 10'h167 == _T_11 ? ram_359 : _GEN_2461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2463 = 10'h168 == _T_11 ? ram_360 : _GEN_2462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2464 = 10'h169 == _T_11 ? ram_361 : _GEN_2463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2465 = 10'h16a == _T_11 ? ram_362 : _GEN_2464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2466 = 10'h16b == _T_11 ? ram_363 : _GEN_2465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2467 = 10'h16c == _T_11 ? ram_364 : _GEN_2466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2468 = 10'h16d == _T_11 ? ram_365 : _GEN_2467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2469 = 10'h16e == _T_11 ? ram_366 : _GEN_2468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2470 = 10'h16f == _T_11 ? ram_367 : _GEN_2469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2471 = 10'h170 == _T_11 ? ram_368 : _GEN_2470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2472 = 10'h171 == _T_11 ? ram_369 : _GEN_2471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2473 = 10'h172 == _T_11 ? ram_370 : _GEN_2472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2474 = 10'h173 == _T_11 ? ram_371 : _GEN_2473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2475 = 10'h174 == _T_11 ? ram_372 : _GEN_2474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2476 = 10'h175 == _T_11 ? ram_373 : _GEN_2475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2477 = 10'h176 == _T_11 ? ram_374 : _GEN_2476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2478 = 10'h177 == _T_11 ? ram_375 : _GEN_2477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2479 = 10'h178 == _T_11 ? ram_376 : _GEN_2478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2480 = 10'h179 == _T_11 ? ram_377 : _GEN_2479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2481 = 10'h17a == _T_11 ? ram_378 : _GEN_2480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2482 = 10'h17b == _T_11 ? ram_379 : _GEN_2481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2483 = 10'h17c == _T_11 ? ram_380 : _GEN_2482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2484 = 10'h17d == _T_11 ? ram_381 : _GEN_2483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2485 = 10'h17e == _T_11 ? ram_382 : _GEN_2484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2486 = 10'h17f == _T_11 ? ram_383 : _GEN_2485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2487 = 10'h180 == _T_11 ? ram_384 : _GEN_2486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2488 = 10'h181 == _T_11 ? ram_385 : _GEN_2487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2489 = 10'h182 == _T_11 ? ram_386 : _GEN_2488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2490 = 10'h183 == _T_11 ? ram_387 : _GEN_2489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2491 = 10'h184 == _T_11 ? ram_388 : _GEN_2490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2492 = 10'h185 == _T_11 ? ram_389 : _GEN_2491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2493 = 10'h186 == _T_11 ? ram_390 : _GEN_2492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2494 = 10'h187 == _T_11 ? ram_391 : _GEN_2493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2495 = 10'h188 == _T_11 ? ram_392 : _GEN_2494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2496 = 10'h189 == _T_11 ? ram_393 : _GEN_2495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2497 = 10'h18a == _T_11 ? ram_394 : _GEN_2496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2498 = 10'h18b == _T_11 ? ram_395 : _GEN_2497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2499 = 10'h18c == _T_11 ? ram_396 : _GEN_2498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2500 = 10'h18d == _T_11 ? ram_397 : _GEN_2499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2501 = 10'h18e == _T_11 ? ram_398 : _GEN_2500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2502 = 10'h18f == _T_11 ? ram_399 : _GEN_2501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2503 = 10'h190 == _T_11 ? ram_400 : _GEN_2502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2504 = 10'h191 == _T_11 ? ram_401 : _GEN_2503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2505 = 10'h192 == _T_11 ? ram_402 : _GEN_2504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2506 = 10'h193 == _T_11 ? ram_403 : _GEN_2505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2507 = 10'h194 == _T_11 ? ram_404 : _GEN_2506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2508 = 10'h195 == _T_11 ? ram_405 : _GEN_2507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2509 = 10'h196 == _T_11 ? ram_406 : _GEN_2508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2510 = 10'h197 == _T_11 ? ram_407 : _GEN_2509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2511 = 10'h198 == _T_11 ? ram_408 : _GEN_2510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2512 = 10'h199 == _T_11 ? ram_409 : _GEN_2511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2513 = 10'h19a == _T_11 ? ram_410 : _GEN_2512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2514 = 10'h19b == _T_11 ? ram_411 : _GEN_2513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2515 = 10'h19c == _T_11 ? ram_412 : _GEN_2514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2516 = 10'h19d == _T_11 ? ram_413 : _GEN_2515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2517 = 10'h19e == _T_11 ? ram_414 : _GEN_2516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2518 = 10'h19f == _T_11 ? ram_415 : _GEN_2517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2519 = 10'h1a0 == _T_11 ? ram_416 : _GEN_2518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2520 = 10'h1a1 == _T_11 ? ram_417 : _GEN_2519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2521 = 10'h1a2 == _T_11 ? ram_418 : _GEN_2520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2522 = 10'h1a3 == _T_11 ? ram_419 : _GEN_2521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2523 = 10'h1a4 == _T_11 ? ram_420 : _GEN_2522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2524 = 10'h1a5 == _T_11 ? ram_421 : _GEN_2523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2525 = 10'h1a6 == _T_11 ? ram_422 : _GEN_2524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2526 = 10'h1a7 == _T_11 ? ram_423 : _GEN_2525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2527 = 10'h1a8 == _T_11 ? ram_424 : _GEN_2526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2528 = 10'h1a9 == _T_11 ? ram_425 : _GEN_2527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2529 = 10'h1aa == _T_11 ? ram_426 : _GEN_2528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2530 = 10'h1ab == _T_11 ? ram_427 : _GEN_2529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2531 = 10'h1ac == _T_11 ? ram_428 : _GEN_2530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2532 = 10'h1ad == _T_11 ? ram_429 : _GEN_2531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2533 = 10'h1ae == _T_11 ? ram_430 : _GEN_2532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2534 = 10'h1af == _T_11 ? ram_431 : _GEN_2533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2535 = 10'h1b0 == _T_11 ? ram_432 : _GEN_2534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2536 = 10'h1b1 == _T_11 ? ram_433 : _GEN_2535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2537 = 10'h1b2 == _T_11 ? ram_434 : _GEN_2536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2538 = 10'h1b3 == _T_11 ? ram_435 : _GEN_2537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2539 = 10'h1b4 == _T_11 ? ram_436 : _GEN_2538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2540 = 10'h1b5 == _T_11 ? ram_437 : _GEN_2539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2541 = 10'h1b6 == _T_11 ? ram_438 : _GEN_2540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2542 = 10'h1b7 == _T_11 ? ram_439 : _GEN_2541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2543 = 10'h1b8 == _T_11 ? ram_440 : _GEN_2542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2544 = 10'h1b9 == _T_11 ? ram_441 : _GEN_2543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2545 = 10'h1ba == _T_11 ? ram_442 : _GEN_2544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2546 = 10'h1bb == _T_11 ? ram_443 : _GEN_2545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2547 = 10'h1bc == _T_11 ? ram_444 : _GEN_2546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2548 = 10'h1bd == _T_11 ? ram_445 : _GEN_2547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2549 = 10'h1be == _T_11 ? ram_446 : _GEN_2548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2550 = 10'h1bf == _T_11 ? ram_447 : _GEN_2549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2551 = 10'h1c0 == _T_11 ? ram_448 : _GEN_2550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2552 = 10'h1c1 == _T_11 ? ram_449 : _GEN_2551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2553 = 10'h1c2 == _T_11 ? ram_450 : _GEN_2552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2554 = 10'h1c3 == _T_11 ? ram_451 : _GEN_2553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2555 = 10'h1c4 == _T_11 ? ram_452 : _GEN_2554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2556 = 10'h1c5 == _T_11 ? ram_453 : _GEN_2555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2557 = 10'h1c6 == _T_11 ? ram_454 : _GEN_2556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2558 = 10'h1c7 == _T_11 ? ram_455 : _GEN_2557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2559 = 10'h1c8 == _T_11 ? ram_456 : _GEN_2558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2560 = 10'h1c9 == _T_11 ? ram_457 : _GEN_2559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2561 = 10'h1ca == _T_11 ? ram_458 : _GEN_2560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2562 = 10'h1cb == _T_11 ? ram_459 : _GEN_2561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2563 = 10'h1cc == _T_11 ? ram_460 : _GEN_2562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2564 = 10'h1cd == _T_11 ? ram_461 : _GEN_2563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2565 = 10'h1ce == _T_11 ? ram_462 : _GEN_2564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2566 = 10'h1cf == _T_11 ? ram_463 : _GEN_2565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2567 = 10'h1d0 == _T_11 ? ram_464 : _GEN_2566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2568 = 10'h1d1 == _T_11 ? ram_465 : _GEN_2567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2569 = 10'h1d2 == _T_11 ? ram_466 : _GEN_2568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2570 = 10'h1d3 == _T_11 ? ram_467 : _GEN_2569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2571 = 10'h1d4 == _T_11 ? ram_468 : _GEN_2570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2572 = 10'h1d5 == _T_11 ? ram_469 : _GEN_2571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2573 = 10'h1d6 == _T_11 ? ram_470 : _GEN_2572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2574 = 10'h1d7 == _T_11 ? ram_471 : _GEN_2573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2575 = 10'h1d8 == _T_11 ? ram_472 : _GEN_2574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2576 = 10'h1d9 == _T_11 ? ram_473 : _GEN_2575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2577 = 10'h1da == _T_11 ? ram_474 : _GEN_2576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2578 = 10'h1db == _T_11 ? ram_475 : _GEN_2577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2579 = 10'h1dc == _T_11 ? ram_476 : _GEN_2578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2580 = 10'h1dd == _T_11 ? ram_477 : _GEN_2579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2581 = 10'h1de == _T_11 ? ram_478 : _GEN_2580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2582 = 10'h1df == _T_11 ? ram_479 : _GEN_2581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2583 = 10'h1e0 == _T_11 ? ram_480 : _GEN_2582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2584 = 10'h1e1 == _T_11 ? ram_481 : _GEN_2583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2585 = 10'h1e2 == _T_11 ? ram_482 : _GEN_2584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2586 = 10'h1e3 == _T_11 ? ram_483 : _GEN_2585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2587 = 10'h1e4 == _T_11 ? ram_484 : _GEN_2586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2588 = 10'h1e5 == _T_11 ? ram_485 : _GEN_2587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2589 = 10'h1e6 == _T_11 ? ram_486 : _GEN_2588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2590 = 10'h1e7 == _T_11 ? ram_487 : _GEN_2589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2591 = 10'h1e8 == _T_11 ? ram_488 : _GEN_2590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2592 = 10'h1e9 == _T_11 ? ram_489 : _GEN_2591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2593 = 10'h1ea == _T_11 ? ram_490 : _GEN_2592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2594 = 10'h1eb == _T_11 ? ram_491 : _GEN_2593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2595 = 10'h1ec == _T_11 ? ram_492 : _GEN_2594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2596 = 10'h1ed == _T_11 ? ram_493 : _GEN_2595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2597 = 10'h1ee == _T_11 ? ram_494 : _GEN_2596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2598 = 10'h1ef == _T_11 ? ram_495 : _GEN_2597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2599 = 10'h1f0 == _T_11 ? ram_496 : _GEN_2598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2600 = 10'h1f1 == _T_11 ? ram_497 : _GEN_2599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2601 = 10'h1f2 == _T_11 ? ram_498 : _GEN_2600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2602 = 10'h1f3 == _T_11 ? ram_499 : _GEN_2601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2603 = 10'h1f4 == _T_11 ? ram_500 : _GEN_2602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2604 = 10'h1f5 == _T_11 ? ram_501 : _GEN_2603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2605 = 10'h1f6 == _T_11 ? ram_502 : _GEN_2604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2606 = 10'h1f7 == _T_11 ? ram_503 : _GEN_2605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2607 = 10'h1f8 == _T_11 ? ram_504 : _GEN_2606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2608 = 10'h1f9 == _T_11 ? ram_505 : _GEN_2607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2609 = 10'h1fa == _T_11 ? ram_506 : _GEN_2608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2610 = 10'h1fb == _T_11 ? ram_507 : _GEN_2609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2611 = 10'h1fc == _T_11 ? ram_508 : _GEN_2610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2612 = 10'h1fd == _T_11 ? ram_509 : _GEN_2611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2613 = 10'h1fe == _T_11 ? ram_510 : _GEN_2612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2614 = 10'h1ff == _T_11 ? ram_511 : _GEN_2613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2615 = 10'h200 == _T_11 ? ram_512 : _GEN_2614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2616 = 10'h201 == _T_11 ? ram_513 : _GEN_2615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2617 = 10'h202 == _T_11 ? ram_514 : _GEN_2616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2618 = 10'h203 == _T_11 ? ram_515 : _GEN_2617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2619 = 10'h204 == _T_11 ? ram_516 : _GEN_2618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2620 = 10'h205 == _T_11 ? ram_517 : _GEN_2619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2621 = 10'h206 == _T_11 ? ram_518 : _GEN_2620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2622 = 10'h207 == _T_11 ? ram_519 : _GEN_2621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2623 = 10'h208 == _T_11 ? ram_520 : _GEN_2622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2624 = 10'h209 == _T_11 ? ram_521 : _GEN_2623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2625 = 10'h20a == _T_11 ? ram_522 : _GEN_2624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2626 = 10'h20b == _T_11 ? ram_523 : _GEN_2625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_2627 = 10'h20c == _T_11 ? ram_524 : _GEN_2626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19065 = {{8190'd0}, _GEN_2627}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_77 = _GEN_19065 ^ _ram_T_76; // @[vga.scala 64:41]
  wire [287:0] _GEN_2628 = 10'h0 == _T_11 ? _ram_T_77[287:0] : _GEN_1578; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2629 = 10'h1 == _T_11 ? _ram_T_77[287:0] : _GEN_1579; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2630 = 10'h2 == _T_11 ? _ram_T_77[287:0] : _GEN_1580; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2631 = 10'h3 == _T_11 ? _ram_T_77[287:0] : _GEN_1581; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2632 = 10'h4 == _T_11 ? _ram_T_77[287:0] : _GEN_1582; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2633 = 10'h5 == _T_11 ? _ram_T_77[287:0] : _GEN_1583; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2634 = 10'h6 == _T_11 ? _ram_T_77[287:0] : _GEN_1584; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2635 = 10'h7 == _T_11 ? _ram_T_77[287:0] : _GEN_1585; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2636 = 10'h8 == _T_11 ? _ram_T_77[287:0] : _GEN_1586; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2637 = 10'h9 == _T_11 ? _ram_T_77[287:0] : _GEN_1587; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2638 = 10'ha == _T_11 ? _ram_T_77[287:0] : _GEN_1588; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2639 = 10'hb == _T_11 ? _ram_T_77[287:0] : _GEN_1589; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2640 = 10'hc == _T_11 ? _ram_T_77[287:0] : _GEN_1590; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2641 = 10'hd == _T_11 ? _ram_T_77[287:0] : _GEN_1591; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2642 = 10'he == _T_11 ? _ram_T_77[287:0] : _GEN_1592; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2643 = 10'hf == _T_11 ? _ram_T_77[287:0] : _GEN_1593; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2644 = 10'h10 == _T_11 ? _ram_T_77[287:0] : _GEN_1594; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2645 = 10'h11 == _T_11 ? _ram_T_77[287:0] : _GEN_1595; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2646 = 10'h12 == _T_11 ? _ram_T_77[287:0] : _GEN_1596; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2647 = 10'h13 == _T_11 ? _ram_T_77[287:0] : _GEN_1597; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2648 = 10'h14 == _T_11 ? _ram_T_77[287:0] : _GEN_1598; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2649 = 10'h15 == _T_11 ? _ram_T_77[287:0] : _GEN_1599; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2650 = 10'h16 == _T_11 ? _ram_T_77[287:0] : _GEN_1600; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2651 = 10'h17 == _T_11 ? _ram_T_77[287:0] : _GEN_1601; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2652 = 10'h18 == _T_11 ? _ram_T_77[287:0] : _GEN_1602; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2653 = 10'h19 == _T_11 ? _ram_T_77[287:0] : _GEN_1603; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2654 = 10'h1a == _T_11 ? _ram_T_77[287:0] : _GEN_1604; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2655 = 10'h1b == _T_11 ? _ram_T_77[287:0] : _GEN_1605; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2656 = 10'h1c == _T_11 ? _ram_T_77[287:0] : _GEN_1606; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2657 = 10'h1d == _T_11 ? _ram_T_77[287:0] : _GEN_1607; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2658 = 10'h1e == _T_11 ? _ram_T_77[287:0] : _GEN_1608; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2659 = 10'h1f == _T_11 ? _ram_T_77[287:0] : _GEN_1609; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2660 = 10'h20 == _T_11 ? _ram_T_77[287:0] : _GEN_1610; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2661 = 10'h21 == _T_11 ? _ram_T_77[287:0] : _GEN_1611; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2662 = 10'h22 == _T_11 ? _ram_T_77[287:0] : _GEN_1612; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2663 = 10'h23 == _T_11 ? _ram_T_77[287:0] : _GEN_1613; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2664 = 10'h24 == _T_11 ? _ram_T_77[287:0] : _GEN_1614; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2665 = 10'h25 == _T_11 ? _ram_T_77[287:0] : _GEN_1615; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2666 = 10'h26 == _T_11 ? _ram_T_77[287:0] : _GEN_1616; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2667 = 10'h27 == _T_11 ? _ram_T_77[287:0] : _GEN_1617; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2668 = 10'h28 == _T_11 ? _ram_T_77[287:0] : _GEN_1618; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2669 = 10'h29 == _T_11 ? _ram_T_77[287:0] : _GEN_1619; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2670 = 10'h2a == _T_11 ? _ram_T_77[287:0] : _GEN_1620; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2671 = 10'h2b == _T_11 ? _ram_T_77[287:0] : _GEN_1621; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2672 = 10'h2c == _T_11 ? _ram_T_77[287:0] : _GEN_1622; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2673 = 10'h2d == _T_11 ? _ram_T_77[287:0] : _GEN_1623; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2674 = 10'h2e == _T_11 ? _ram_T_77[287:0] : _GEN_1624; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2675 = 10'h2f == _T_11 ? _ram_T_77[287:0] : _GEN_1625; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2676 = 10'h30 == _T_11 ? _ram_T_77[287:0] : _GEN_1626; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2677 = 10'h31 == _T_11 ? _ram_T_77[287:0] : _GEN_1627; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2678 = 10'h32 == _T_11 ? _ram_T_77[287:0] : _GEN_1628; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2679 = 10'h33 == _T_11 ? _ram_T_77[287:0] : _GEN_1629; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2680 = 10'h34 == _T_11 ? _ram_T_77[287:0] : _GEN_1630; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2681 = 10'h35 == _T_11 ? _ram_T_77[287:0] : _GEN_1631; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2682 = 10'h36 == _T_11 ? _ram_T_77[287:0] : _GEN_1632; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2683 = 10'h37 == _T_11 ? _ram_T_77[287:0] : _GEN_1633; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2684 = 10'h38 == _T_11 ? _ram_T_77[287:0] : _GEN_1634; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2685 = 10'h39 == _T_11 ? _ram_T_77[287:0] : _GEN_1635; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2686 = 10'h3a == _T_11 ? _ram_T_77[287:0] : _GEN_1636; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2687 = 10'h3b == _T_11 ? _ram_T_77[287:0] : _GEN_1637; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2688 = 10'h3c == _T_11 ? _ram_T_77[287:0] : _GEN_1638; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2689 = 10'h3d == _T_11 ? _ram_T_77[287:0] : _GEN_1639; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2690 = 10'h3e == _T_11 ? _ram_T_77[287:0] : _GEN_1640; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2691 = 10'h3f == _T_11 ? _ram_T_77[287:0] : _GEN_1641; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2692 = 10'h40 == _T_11 ? _ram_T_77[287:0] : _GEN_1642; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2693 = 10'h41 == _T_11 ? _ram_T_77[287:0] : _GEN_1643; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2694 = 10'h42 == _T_11 ? _ram_T_77[287:0] : _GEN_1644; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2695 = 10'h43 == _T_11 ? _ram_T_77[287:0] : _GEN_1645; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2696 = 10'h44 == _T_11 ? _ram_T_77[287:0] : _GEN_1646; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2697 = 10'h45 == _T_11 ? _ram_T_77[287:0] : _GEN_1647; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2698 = 10'h46 == _T_11 ? _ram_T_77[287:0] : _GEN_1648; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2699 = 10'h47 == _T_11 ? _ram_T_77[287:0] : _GEN_1649; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2700 = 10'h48 == _T_11 ? _ram_T_77[287:0] : _GEN_1650; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2701 = 10'h49 == _T_11 ? _ram_T_77[287:0] : _GEN_1651; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2702 = 10'h4a == _T_11 ? _ram_T_77[287:0] : _GEN_1652; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2703 = 10'h4b == _T_11 ? _ram_T_77[287:0] : _GEN_1653; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2704 = 10'h4c == _T_11 ? _ram_T_77[287:0] : _GEN_1654; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2705 = 10'h4d == _T_11 ? _ram_T_77[287:0] : _GEN_1655; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2706 = 10'h4e == _T_11 ? _ram_T_77[287:0] : _GEN_1656; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2707 = 10'h4f == _T_11 ? _ram_T_77[287:0] : _GEN_1657; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2708 = 10'h50 == _T_11 ? _ram_T_77[287:0] : _GEN_1658; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2709 = 10'h51 == _T_11 ? _ram_T_77[287:0] : _GEN_1659; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2710 = 10'h52 == _T_11 ? _ram_T_77[287:0] : _GEN_1660; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2711 = 10'h53 == _T_11 ? _ram_T_77[287:0] : _GEN_1661; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2712 = 10'h54 == _T_11 ? _ram_T_77[287:0] : _GEN_1662; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2713 = 10'h55 == _T_11 ? _ram_T_77[287:0] : _GEN_1663; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2714 = 10'h56 == _T_11 ? _ram_T_77[287:0] : _GEN_1664; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2715 = 10'h57 == _T_11 ? _ram_T_77[287:0] : _GEN_1665; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2716 = 10'h58 == _T_11 ? _ram_T_77[287:0] : _GEN_1666; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2717 = 10'h59 == _T_11 ? _ram_T_77[287:0] : _GEN_1667; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2718 = 10'h5a == _T_11 ? _ram_T_77[287:0] : _GEN_1668; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2719 = 10'h5b == _T_11 ? _ram_T_77[287:0] : _GEN_1669; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2720 = 10'h5c == _T_11 ? _ram_T_77[287:0] : _GEN_1670; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2721 = 10'h5d == _T_11 ? _ram_T_77[287:0] : _GEN_1671; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2722 = 10'h5e == _T_11 ? _ram_T_77[287:0] : _GEN_1672; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2723 = 10'h5f == _T_11 ? _ram_T_77[287:0] : _GEN_1673; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2724 = 10'h60 == _T_11 ? _ram_T_77[287:0] : _GEN_1674; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2725 = 10'h61 == _T_11 ? _ram_T_77[287:0] : _GEN_1675; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2726 = 10'h62 == _T_11 ? _ram_T_77[287:0] : _GEN_1676; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2727 = 10'h63 == _T_11 ? _ram_T_77[287:0] : _GEN_1677; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2728 = 10'h64 == _T_11 ? _ram_T_77[287:0] : _GEN_1678; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2729 = 10'h65 == _T_11 ? _ram_T_77[287:0] : _GEN_1679; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2730 = 10'h66 == _T_11 ? _ram_T_77[287:0] : _GEN_1680; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2731 = 10'h67 == _T_11 ? _ram_T_77[287:0] : _GEN_1681; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2732 = 10'h68 == _T_11 ? _ram_T_77[287:0] : _GEN_1682; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2733 = 10'h69 == _T_11 ? _ram_T_77[287:0] : _GEN_1683; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2734 = 10'h6a == _T_11 ? _ram_T_77[287:0] : _GEN_1684; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2735 = 10'h6b == _T_11 ? _ram_T_77[287:0] : _GEN_1685; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2736 = 10'h6c == _T_11 ? _ram_T_77[287:0] : _GEN_1686; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2737 = 10'h6d == _T_11 ? _ram_T_77[287:0] : _GEN_1687; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2738 = 10'h6e == _T_11 ? _ram_T_77[287:0] : _GEN_1688; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2739 = 10'h6f == _T_11 ? _ram_T_77[287:0] : _GEN_1689; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2740 = 10'h70 == _T_11 ? _ram_T_77[287:0] : _GEN_1690; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2741 = 10'h71 == _T_11 ? _ram_T_77[287:0] : _GEN_1691; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2742 = 10'h72 == _T_11 ? _ram_T_77[287:0] : _GEN_1692; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2743 = 10'h73 == _T_11 ? _ram_T_77[287:0] : _GEN_1693; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2744 = 10'h74 == _T_11 ? _ram_T_77[287:0] : _GEN_1694; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2745 = 10'h75 == _T_11 ? _ram_T_77[287:0] : _GEN_1695; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2746 = 10'h76 == _T_11 ? _ram_T_77[287:0] : _GEN_1696; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2747 = 10'h77 == _T_11 ? _ram_T_77[287:0] : _GEN_1697; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2748 = 10'h78 == _T_11 ? _ram_T_77[287:0] : _GEN_1698; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2749 = 10'h79 == _T_11 ? _ram_T_77[287:0] : _GEN_1699; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2750 = 10'h7a == _T_11 ? _ram_T_77[287:0] : _GEN_1700; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2751 = 10'h7b == _T_11 ? _ram_T_77[287:0] : _GEN_1701; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2752 = 10'h7c == _T_11 ? _ram_T_77[287:0] : _GEN_1702; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2753 = 10'h7d == _T_11 ? _ram_T_77[287:0] : _GEN_1703; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2754 = 10'h7e == _T_11 ? _ram_T_77[287:0] : _GEN_1704; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2755 = 10'h7f == _T_11 ? _ram_T_77[287:0] : _GEN_1705; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2756 = 10'h80 == _T_11 ? _ram_T_77[287:0] : _GEN_1706; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2757 = 10'h81 == _T_11 ? _ram_T_77[287:0] : _GEN_1707; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2758 = 10'h82 == _T_11 ? _ram_T_77[287:0] : _GEN_1708; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2759 = 10'h83 == _T_11 ? _ram_T_77[287:0] : _GEN_1709; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2760 = 10'h84 == _T_11 ? _ram_T_77[287:0] : _GEN_1710; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2761 = 10'h85 == _T_11 ? _ram_T_77[287:0] : _GEN_1711; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2762 = 10'h86 == _T_11 ? _ram_T_77[287:0] : _GEN_1712; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2763 = 10'h87 == _T_11 ? _ram_T_77[287:0] : _GEN_1713; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2764 = 10'h88 == _T_11 ? _ram_T_77[287:0] : _GEN_1714; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2765 = 10'h89 == _T_11 ? _ram_T_77[287:0] : _GEN_1715; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2766 = 10'h8a == _T_11 ? _ram_T_77[287:0] : _GEN_1716; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2767 = 10'h8b == _T_11 ? _ram_T_77[287:0] : _GEN_1717; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2768 = 10'h8c == _T_11 ? _ram_T_77[287:0] : _GEN_1718; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2769 = 10'h8d == _T_11 ? _ram_T_77[287:0] : _GEN_1719; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2770 = 10'h8e == _T_11 ? _ram_T_77[287:0] : _GEN_1720; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2771 = 10'h8f == _T_11 ? _ram_T_77[287:0] : _GEN_1721; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2772 = 10'h90 == _T_11 ? _ram_T_77[287:0] : _GEN_1722; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2773 = 10'h91 == _T_11 ? _ram_T_77[287:0] : _GEN_1723; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2774 = 10'h92 == _T_11 ? _ram_T_77[287:0] : _GEN_1724; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2775 = 10'h93 == _T_11 ? _ram_T_77[287:0] : _GEN_1725; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2776 = 10'h94 == _T_11 ? _ram_T_77[287:0] : _GEN_1726; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2777 = 10'h95 == _T_11 ? _ram_T_77[287:0] : _GEN_1727; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2778 = 10'h96 == _T_11 ? _ram_T_77[287:0] : _GEN_1728; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2779 = 10'h97 == _T_11 ? _ram_T_77[287:0] : _GEN_1729; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2780 = 10'h98 == _T_11 ? _ram_T_77[287:0] : _GEN_1730; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2781 = 10'h99 == _T_11 ? _ram_T_77[287:0] : _GEN_1731; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2782 = 10'h9a == _T_11 ? _ram_T_77[287:0] : _GEN_1732; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2783 = 10'h9b == _T_11 ? _ram_T_77[287:0] : _GEN_1733; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2784 = 10'h9c == _T_11 ? _ram_T_77[287:0] : _GEN_1734; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2785 = 10'h9d == _T_11 ? _ram_T_77[287:0] : _GEN_1735; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2786 = 10'h9e == _T_11 ? _ram_T_77[287:0] : _GEN_1736; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2787 = 10'h9f == _T_11 ? _ram_T_77[287:0] : _GEN_1737; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2788 = 10'ha0 == _T_11 ? _ram_T_77[287:0] : _GEN_1738; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2789 = 10'ha1 == _T_11 ? _ram_T_77[287:0] : _GEN_1739; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2790 = 10'ha2 == _T_11 ? _ram_T_77[287:0] : _GEN_1740; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2791 = 10'ha3 == _T_11 ? _ram_T_77[287:0] : _GEN_1741; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2792 = 10'ha4 == _T_11 ? _ram_T_77[287:0] : _GEN_1742; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2793 = 10'ha5 == _T_11 ? _ram_T_77[287:0] : _GEN_1743; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2794 = 10'ha6 == _T_11 ? _ram_T_77[287:0] : _GEN_1744; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2795 = 10'ha7 == _T_11 ? _ram_T_77[287:0] : _GEN_1745; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2796 = 10'ha8 == _T_11 ? _ram_T_77[287:0] : _GEN_1746; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2797 = 10'ha9 == _T_11 ? _ram_T_77[287:0] : _GEN_1747; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2798 = 10'haa == _T_11 ? _ram_T_77[287:0] : _GEN_1748; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2799 = 10'hab == _T_11 ? _ram_T_77[287:0] : _GEN_1749; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2800 = 10'hac == _T_11 ? _ram_T_77[287:0] : _GEN_1750; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2801 = 10'had == _T_11 ? _ram_T_77[287:0] : _GEN_1751; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2802 = 10'hae == _T_11 ? _ram_T_77[287:0] : _GEN_1752; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2803 = 10'haf == _T_11 ? _ram_T_77[287:0] : _GEN_1753; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2804 = 10'hb0 == _T_11 ? _ram_T_77[287:0] : _GEN_1754; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2805 = 10'hb1 == _T_11 ? _ram_T_77[287:0] : _GEN_1755; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2806 = 10'hb2 == _T_11 ? _ram_T_77[287:0] : _GEN_1756; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2807 = 10'hb3 == _T_11 ? _ram_T_77[287:0] : _GEN_1757; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2808 = 10'hb4 == _T_11 ? _ram_T_77[287:0] : _GEN_1758; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2809 = 10'hb5 == _T_11 ? _ram_T_77[287:0] : _GEN_1759; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2810 = 10'hb6 == _T_11 ? _ram_T_77[287:0] : _GEN_1760; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2811 = 10'hb7 == _T_11 ? _ram_T_77[287:0] : _GEN_1761; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2812 = 10'hb8 == _T_11 ? _ram_T_77[287:0] : _GEN_1762; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2813 = 10'hb9 == _T_11 ? _ram_T_77[287:0] : _GEN_1763; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2814 = 10'hba == _T_11 ? _ram_T_77[287:0] : _GEN_1764; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2815 = 10'hbb == _T_11 ? _ram_T_77[287:0] : _GEN_1765; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2816 = 10'hbc == _T_11 ? _ram_T_77[287:0] : _GEN_1766; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2817 = 10'hbd == _T_11 ? _ram_T_77[287:0] : _GEN_1767; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2818 = 10'hbe == _T_11 ? _ram_T_77[287:0] : _GEN_1768; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2819 = 10'hbf == _T_11 ? _ram_T_77[287:0] : _GEN_1769; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2820 = 10'hc0 == _T_11 ? _ram_T_77[287:0] : _GEN_1770; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2821 = 10'hc1 == _T_11 ? _ram_T_77[287:0] : _GEN_1771; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2822 = 10'hc2 == _T_11 ? _ram_T_77[287:0] : _GEN_1772; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2823 = 10'hc3 == _T_11 ? _ram_T_77[287:0] : _GEN_1773; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2824 = 10'hc4 == _T_11 ? _ram_T_77[287:0] : _GEN_1774; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2825 = 10'hc5 == _T_11 ? _ram_T_77[287:0] : _GEN_1775; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2826 = 10'hc6 == _T_11 ? _ram_T_77[287:0] : _GEN_1776; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2827 = 10'hc7 == _T_11 ? _ram_T_77[287:0] : _GEN_1777; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2828 = 10'hc8 == _T_11 ? _ram_T_77[287:0] : _GEN_1778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2829 = 10'hc9 == _T_11 ? _ram_T_77[287:0] : _GEN_1779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2830 = 10'hca == _T_11 ? _ram_T_77[287:0] : _GEN_1780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2831 = 10'hcb == _T_11 ? _ram_T_77[287:0] : _GEN_1781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2832 = 10'hcc == _T_11 ? _ram_T_77[287:0] : _GEN_1782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2833 = 10'hcd == _T_11 ? _ram_T_77[287:0] : _GEN_1783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2834 = 10'hce == _T_11 ? _ram_T_77[287:0] : _GEN_1784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2835 = 10'hcf == _T_11 ? _ram_T_77[287:0] : _GEN_1785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2836 = 10'hd0 == _T_11 ? _ram_T_77[287:0] : _GEN_1786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2837 = 10'hd1 == _T_11 ? _ram_T_77[287:0] : _GEN_1787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2838 = 10'hd2 == _T_11 ? _ram_T_77[287:0] : _GEN_1788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2839 = 10'hd3 == _T_11 ? _ram_T_77[287:0] : _GEN_1789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2840 = 10'hd4 == _T_11 ? _ram_T_77[287:0] : _GEN_1790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2841 = 10'hd5 == _T_11 ? _ram_T_77[287:0] : _GEN_1791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2842 = 10'hd6 == _T_11 ? _ram_T_77[287:0] : _GEN_1792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2843 = 10'hd7 == _T_11 ? _ram_T_77[287:0] : _GEN_1793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2844 = 10'hd8 == _T_11 ? _ram_T_77[287:0] : _GEN_1794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2845 = 10'hd9 == _T_11 ? _ram_T_77[287:0] : _GEN_1795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2846 = 10'hda == _T_11 ? _ram_T_77[287:0] : _GEN_1796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2847 = 10'hdb == _T_11 ? _ram_T_77[287:0] : _GEN_1797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2848 = 10'hdc == _T_11 ? _ram_T_77[287:0] : _GEN_1798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2849 = 10'hdd == _T_11 ? _ram_T_77[287:0] : _GEN_1799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2850 = 10'hde == _T_11 ? _ram_T_77[287:0] : _GEN_1800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2851 = 10'hdf == _T_11 ? _ram_T_77[287:0] : _GEN_1801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2852 = 10'he0 == _T_11 ? _ram_T_77[287:0] : _GEN_1802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2853 = 10'he1 == _T_11 ? _ram_T_77[287:0] : _GEN_1803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2854 = 10'he2 == _T_11 ? _ram_T_77[287:0] : _GEN_1804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2855 = 10'he3 == _T_11 ? _ram_T_77[287:0] : _GEN_1805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2856 = 10'he4 == _T_11 ? _ram_T_77[287:0] : _GEN_1806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2857 = 10'he5 == _T_11 ? _ram_T_77[287:0] : _GEN_1807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2858 = 10'he6 == _T_11 ? _ram_T_77[287:0] : _GEN_1808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2859 = 10'he7 == _T_11 ? _ram_T_77[287:0] : _GEN_1809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2860 = 10'he8 == _T_11 ? _ram_T_77[287:0] : _GEN_1810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2861 = 10'he9 == _T_11 ? _ram_T_77[287:0] : _GEN_1811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2862 = 10'hea == _T_11 ? _ram_T_77[287:0] : _GEN_1812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2863 = 10'heb == _T_11 ? _ram_T_77[287:0] : _GEN_1813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2864 = 10'hec == _T_11 ? _ram_T_77[287:0] : _GEN_1814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2865 = 10'hed == _T_11 ? _ram_T_77[287:0] : _GEN_1815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2866 = 10'hee == _T_11 ? _ram_T_77[287:0] : _GEN_1816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2867 = 10'hef == _T_11 ? _ram_T_77[287:0] : _GEN_1817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2868 = 10'hf0 == _T_11 ? _ram_T_77[287:0] : _GEN_1818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2869 = 10'hf1 == _T_11 ? _ram_T_77[287:0] : _GEN_1819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2870 = 10'hf2 == _T_11 ? _ram_T_77[287:0] : _GEN_1820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2871 = 10'hf3 == _T_11 ? _ram_T_77[287:0] : _GEN_1821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2872 = 10'hf4 == _T_11 ? _ram_T_77[287:0] : _GEN_1822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2873 = 10'hf5 == _T_11 ? _ram_T_77[287:0] : _GEN_1823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2874 = 10'hf6 == _T_11 ? _ram_T_77[287:0] : _GEN_1824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2875 = 10'hf7 == _T_11 ? _ram_T_77[287:0] : _GEN_1825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2876 = 10'hf8 == _T_11 ? _ram_T_77[287:0] : _GEN_1826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2877 = 10'hf9 == _T_11 ? _ram_T_77[287:0] : _GEN_1827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2878 = 10'hfa == _T_11 ? _ram_T_77[287:0] : _GEN_1828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2879 = 10'hfb == _T_11 ? _ram_T_77[287:0] : _GEN_1829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2880 = 10'hfc == _T_11 ? _ram_T_77[287:0] : _GEN_1830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2881 = 10'hfd == _T_11 ? _ram_T_77[287:0] : _GEN_1831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2882 = 10'hfe == _T_11 ? _ram_T_77[287:0] : _GEN_1832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2883 = 10'hff == _T_11 ? _ram_T_77[287:0] : _GEN_1833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2884 = 10'h100 == _T_11 ? _ram_T_77[287:0] : _GEN_1834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2885 = 10'h101 == _T_11 ? _ram_T_77[287:0] : _GEN_1835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2886 = 10'h102 == _T_11 ? _ram_T_77[287:0] : _GEN_1836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2887 = 10'h103 == _T_11 ? _ram_T_77[287:0] : _GEN_1837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2888 = 10'h104 == _T_11 ? _ram_T_77[287:0] : _GEN_1838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2889 = 10'h105 == _T_11 ? _ram_T_77[287:0] : _GEN_1839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2890 = 10'h106 == _T_11 ? _ram_T_77[287:0] : _GEN_1840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2891 = 10'h107 == _T_11 ? _ram_T_77[287:0] : _GEN_1841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2892 = 10'h108 == _T_11 ? _ram_T_77[287:0] : _GEN_1842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2893 = 10'h109 == _T_11 ? _ram_T_77[287:0] : _GEN_1843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2894 = 10'h10a == _T_11 ? _ram_T_77[287:0] : _GEN_1844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2895 = 10'h10b == _T_11 ? _ram_T_77[287:0] : _GEN_1845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2896 = 10'h10c == _T_11 ? _ram_T_77[287:0] : _GEN_1846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2897 = 10'h10d == _T_11 ? _ram_T_77[287:0] : _GEN_1847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2898 = 10'h10e == _T_11 ? _ram_T_77[287:0] : _GEN_1848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2899 = 10'h10f == _T_11 ? _ram_T_77[287:0] : _GEN_1849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2900 = 10'h110 == _T_11 ? _ram_T_77[287:0] : _GEN_1850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2901 = 10'h111 == _T_11 ? _ram_T_77[287:0] : _GEN_1851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2902 = 10'h112 == _T_11 ? _ram_T_77[287:0] : _GEN_1852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2903 = 10'h113 == _T_11 ? _ram_T_77[287:0] : _GEN_1853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2904 = 10'h114 == _T_11 ? _ram_T_77[287:0] : _GEN_1854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2905 = 10'h115 == _T_11 ? _ram_T_77[287:0] : _GEN_1855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2906 = 10'h116 == _T_11 ? _ram_T_77[287:0] : _GEN_1856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2907 = 10'h117 == _T_11 ? _ram_T_77[287:0] : _GEN_1857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2908 = 10'h118 == _T_11 ? _ram_T_77[287:0] : _GEN_1858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2909 = 10'h119 == _T_11 ? _ram_T_77[287:0] : _GEN_1859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2910 = 10'h11a == _T_11 ? _ram_T_77[287:0] : _GEN_1860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2911 = 10'h11b == _T_11 ? _ram_T_77[287:0] : _GEN_1861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2912 = 10'h11c == _T_11 ? _ram_T_77[287:0] : _GEN_1862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2913 = 10'h11d == _T_11 ? _ram_T_77[287:0] : _GEN_1863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2914 = 10'h11e == _T_11 ? _ram_T_77[287:0] : _GEN_1864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2915 = 10'h11f == _T_11 ? _ram_T_77[287:0] : _GEN_1865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2916 = 10'h120 == _T_11 ? _ram_T_77[287:0] : _GEN_1866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2917 = 10'h121 == _T_11 ? _ram_T_77[287:0] : _GEN_1867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2918 = 10'h122 == _T_11 ? _ram_T_77[287:0] : _GEN_1868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2919 = 10'h123 == _T_11 ? _ram_T_77[287:0] : _GEN_1869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2920 = 10'h124 == _T_11 ? _ram_T_77[287:0] : _GEN_1870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2921 = 10'h125 == _T_11 ? _ram_T_77[287:0] : _GEN_1871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2922 = 10'h126 == _T_11 ? _ram_T_77[287:0] : _GEN_1872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2923 = 10'h127 == _T_11 ? _ram_T_77[287:0] : _GEN_1873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2924 = 10'h128 == _T_11 ? _ram_T_77[287:0] : _GEN_1874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2925 = 10'h129 == _T_11 ? _ram_T_77[287:0] : _GEN_1875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2926 = 10'h12a == _T_11 ? _ram_T_77[287:0] : _GEN_1876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2927 = 10'h12b == _T_11 ? _ram_T_77[287:0] : _GEN_1877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2928 = 10'h12c == _T_11 ? _ram_T_77[287:0] : _GEN_1878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2929 = 10'h12d == _T_11 ? _ram_T_77[287:0] : _GEN_1879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2930 = 10'h12e == _T_11 ? _ram_T_77[287:0] : _GEN_1880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2931 = 10'h12f == _T_11 ? _ram_T_77[287:0] : _GEN_1881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2932 = 10'h130 == _T_11 ? _ram_T_77[287:0] : _GEN_1882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2933 = 10'h131 == _T_11 ? _ram_T_77[287:0] : _GEN_1883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2934 = 10'h132 == _T_11 ? _ram_T_77[287:0] : _GEN_1884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2935 = 10'h133 == _T_11 ? _ram_T_77[287:0] : _GEN_1885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2936 = 10'h134 == _T_11 ? _ram_T_77[287:0] : _GEN_1886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2937 = 10'h135 == _T_11 ? _ram_T_77[287:0] : _GEN_1887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2938 = 10'h136 == _T_11 ? _ram_T_77[287:0] : _GEN_1888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2939 = 10'h137 == _T_11 ? _ram_T_77[287:0] : _GEN_1889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2940 = 10'h138 == _T_11 ? _ram_T_77[287:0] : _GEN_1890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2941 = 10'h139 == _T_11 ? _ram_T_77[287:0] : _GEN_1891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2942 = 10'h13a == _T_11 ? _ram_T_77[287:0] : _GEN_1892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2943 = 10'h13b == _T_11 ? _ram_T_77[287:0] : _GEN_1893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2944 = 10'h13c == _T_11 ? _ram_T_77[287:0] : _GEN_1894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2945 = 10'h13d == _T_11 ? _ram_T_77[287:0] : _GEN_1895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2946 = 10'h13e == _T_11 ? _ram_T_77[287:0] : _GEN_1896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2947 = 10'h13f == _T_11 ? _ram_T_77[287:0] : _GEN_1897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2948 = 10'h140 == _T_11 ? _ram_T_77[287:0] : _GEN_1898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2949 = 10'h141 == _T_11 ? _ram_T_77[287:0] : _GEN_1899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2950 = 10'h142 == _T_11 ? _ram_T_77[287:0] : _GEN_1900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2951 = 10'h143 == _T_11 ? _ram_T_77[287:0] : _GEN_1901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2952 = 10'h144 == _T_11 ? _ram_T_77[287:0] : _GEN_1902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2953 = 10'h145 == _T_11 ? _ram_T_77[287:0] : _GEN_1903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2954 = 10'h146 == _T_11 ? _ram_T_77[287:0] : _GEN_1904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2955 = 10'h147 == _T_11 ? _ram_T_77[287:0] : _GEN_1905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2956 = 10'h148 == _T_11 ? _ram_T_77[287:0] : _GEN_1906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2957 = 10'h149 == _T_11 ? _ram_T_77[287:0] : _GEN_1907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2958 = 10'h14a == _T_11 ? _ram_T_77[287:0] : _GEN_1908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2959 = 10'h14b == _T_11 ? _ram_T_77[287:0] : _GEN_1909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2960 = 10'h14c == _T_11 ? _ram_T_77[287:0] : _GEN_1910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2961 = 10'h14d == _T_11 ? _ram_T_77[287:0] : _GEN_1911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2962 = 10'h14e == _T_11 ? _ram_T_77[287:0] : _GEN_1912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2963 = 10'h14f == _T_11 ? _ram_T_77[287:0] : _GEN_1913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2964 = 10'h150 == _T_11 ? _ram_T_77[287:0] : _GEN_1914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2965 = 10'h151 == _T_11 ? _ram_T_77[287:0] : _GEN_1915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2966 = 10'h152 == _T_11 ? _ram_T_77[287:0] : _GEN_1916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2967 = 10'h153 == _T_11 ? _ram_T_77[287:0] : _GEN_1917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2968 = 10'h154 == _T_11 ? _ram_T_77[287:0] : _GEN_1918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2969 = 10'h155 == _T_11 ? _ram_T_77[287:0] : _GEN_1919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2970 = 10'h156 == _T_11 ? _ram_T_77[287:0] : _GEN_1920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2971 = 10'h157 == _T_11 ? _ram_T_77[287:0] : _GEN_1921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2972 = 10'h158 == _T_11 ? _ram_T_77[287:0] : _GEN_1922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2973 = 10'h159 == _T_11 ? _ram_T_77[287:0] : _GEN_1923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2974 = 10'h15a == _T_11 ? _ram_T_77[287:0] : _GEN_1924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2975 = 10'h15b == _T_11 ? _ram_T_77[287:0] : _GEN_1925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2976 = 10'h15c == _T_11 ? _ram_T_77[287:0] : _GEN_1926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2977 = 10'h15d == _T_11 ? _ram_T_77[287:0] : _GEN_1927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2978 = 10'h15e == _T_11 ? _ram_T_77[287:0] : _GEN_1928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2979 = 10'h15f == _T_11 ? _ram_T_77[287:0] : _GEN_1929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2980 = 10'h160 == _T_11 ? _ram_T_77[287:0] : _GEN_1930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2981 = 10'h161 == _T_11 ? _ram_T_77[287:0] : _GEN_1931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2982 = 10'h162 == _T_11 ? _ram_T_77[287:0] : _GEN_1932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2983 = 10'h163 == _T_11 ? _ram_T_77[287:0] : _GEN_1933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2984 = 10'h164 == _T_11 ? _ram_T_77[287:0] : _GEN_1934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2985 = 10'h165 == _T_11 ? _ram_T_77[287:0] : _GEN_1935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2986 = 10'h166 == _T_11 ? _ram_T_77[287:0] : _GEN_1936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2987 = 10'h167 == _T_11 ? _ram_T_77[287:0] : _GEN_1937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2988 = 10'h168 == _T_11 ? _ram_T_77[287:0] : _GEN_1938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2989 = 10'h169 == _T_11 ? _ram_T_77[287:0] : _GEN_1939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2990 = 10'h16a == _T_11 ? _ram_T_77[287:0] : _GEN_1940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2991 = 10'h16b == _T_11 ? _ram_T_77[287:0] : _GEN_1941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2992 = 10'h16c == _T_11 ? _ram_T_77[287:0] : _GEN_1942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2993 = 10'h16d == _T_11 ? _ram_T_77[287:0] : _GEN_1943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2994 = 10'h16e == _T_11 ? _ram_T_77[287:0] : _GEN_1944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2995 = 10'h16f == _T_11 ? _ram_T_77[287:0] : _GEN_1945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2996 = 10'h170 == _T_11 ? _ram_T_77[287:0] : _GEN_1946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2997 = 10'h171 == _T_11 ? _ram_T_77[287:0] : _GEN_1947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2998 = 10'h172 == _T_11 ? _ram_T_77[287:0] : _GEN_1948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_2999 = 10'h173 == _T_11 ? _ram_T_77[287:0] : _GEN_1949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3000 = 10'h174 == _T_11 ? _ram_T_77[287:0] : _GEN_1950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3001 = 10'h175 == _T_11 ? _ram_T_77[287:0] : _GEN_1951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3002 = 10'h176 == _T_11 ? _ram_T_77[287:0] : _GEN_1952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3003 = 10'h177 == _T_11 ? _ram_T_77[287:0] : _GEN_1953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3004 = 10'h178 == _T_11 ? _ram_T_77[287:0] : _GEN_1954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3005 = 10'h179 == _T_11 ? _ram_T_77[287:0] : _GEN_1955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3006 = 10'h17a == _T_11 ? _ram_T_77[287:0] : _GEN_1956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3007 = 10'h17b == _T_11 ? _ram_T_77[287:0] : _GEN_1957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3008 = 10'h17c == _T_11 ? _ram_T_77[287:0] : _GEN_1958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3009 = 10'h17d == _T_11 ? _ram_T_77[287:0] : _GEN_1959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3010 = 10'h17e == _T_11 ? _ram_T_77[287:0] : _GEN_1960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3011 = 10'h17f == _T_11 ? _ram_T_77[287:0] : _GEN_1961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3012 = 10'h180 == _T_11 ? _ram_T_77[287:0] : _GEN_1962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3013 = 10'h181 == _T_11 ? _ram_T_77[287:0] : _GEN_1963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3014 = 10'h182 == _T_11 ? _ram_T_77[287:0] : _GEN_1964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3015 = 10'h183 == _T_11 ? _ram_T_77[287:0] : _GEN_1965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3016 = 10'h184 == _T_11 ? _ram_T_77[287:0] : _GEN_1966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3017 = 10'h185 == _T_11 ? _ram_T_77[287:0] : _GEN_1967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3018 = 10'h186 == _T_11 ? _ram_T_77[287:0] : _GEN_1968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3019 = 10'h187 == _T_11 ? _ram_T_77[287:0] : _GEN_1969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3020 = 10'h188 == _T_11 ? _ram_T_77[287:0] : _GEN_1970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3021 = 10'h189 == _T_11 ? _ram_T_77[287:0] : _GEN_1971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3022 = 10'h18a == _T_11 ? _ram_T_77[287:0] : _GEN_1972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3023 = 10'h18b == _T_11 ? _ram_T_77[287:0] : _GEN_1973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3024 = 10'h18c == _T_11 ? _ram_T_77[287:0] : _GEN_1974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3025 = 10'h18d == _T_11 ? _ram_T_77[287:0] : _GEN_1975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3026 = 10'h18e == _T_11 ? _ram_T_77[287:0] : _GEN_1976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3027 = 10'h18f == _T_11 ? _ram_T_77[287:0] : _GEN_1977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3028 = 10'h190 == _T_11 ? _ram_T_77[287:0] : _GEN_1978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3029 = 10'h191 == _T_11 ? _ram_T_77[287:0] : _GEN_1979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3030 = 10'h192 == _T_11 ? _ram_T_77[287:0] : _GEN_1980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3031 = 10'h193 == _T_11 ? _ram_T_77[287:0] : _GEN_1981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3032 = 10'h194 == _T_11 ? _ram_T_77[287:0] : _GEN_1982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3033 = 10'h195 == _T_11 ? _ram_T_77[287:0] : _GEN_1983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3034 = 10'h196 == _T_11 ? _ram_T_77[287:0] : _GEN_1984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3035 = 10'h197 == _T_11 ? _ram_T_77[287:0] : _GEN_1985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3036 = 10'h198 == _T_11 ? _ram_T_77[287:0] : _GEN_1986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3037 = 10'h199 == _T_11 ? _ram_T_77[287:0] : _GEN_1987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3038 = 10'h19a == _T_11 ? _ram_T_77[287:0] : _GEN_1988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3039 = 10'h19b == _T_11 ? _ram_T_77[287:0] : _GEN_1989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3040 = 10'h19c == _T_11 ? _ram_T_77[287:0] : _GEN_1990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3041 = 10'h19d == _T_11 ? _ram_T_77[287:0] : _GEN_1991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3042 = 10'h19e == _T_11 ? _ram_T_77[287:0] : _GEN_1992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3043 = 10'h19f == _T_11 ? _ram_T_77[287:0] : _GEN_1993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3044 = 10'h1a0 == _T_11 ? _ram_T_77[287:0] : _GEN_1994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3045 = 10'h1a1 == _T_11 ? _ram_T_77[287:0] : _GEN_1995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3046 = 10'h1a2 == _T_11 ? _ram_T_77[287:0] : _GEN_1996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3047 = 10'h1a3 == _T_11 ? _ram_T_77[287:0] : _GEN_1997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3048 = 10'h1a4 == _T_11 ? _ram_T_77[287:0] : _GEN_1998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3049 = 10'h1a5 == _T_11 ? _ram_T_77[287:0] : _GEN_1999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3050 = 10'h1a6 == _T_11 ? _ram_T_77[287:0] : _GEN_2000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3051 = 10'h1a7 == _T_11 ? _ram_T_77[287:0] : _GEN_2001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3052 = 10'h1a8 == _T_11 ? _ram_T_77[287:0] : _GEN_2002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3053 = 10'h1a9 == _T_11 ? _ram_T_77[287:0] : _GEN_2003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3054 = 10'h1aa == _T_11 ? _ram_T_77[287:0] : _GEN_2004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3055 = 10'h1ab == _T_11 ? _ram_T_77[287:0] : _GEN_2005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3056 = 10'h1ac == _T_11 ? _ram_T_77[287:0] : _GEN_2006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3057 = 10'h1ad == _T_11 ? _ram_T_77[287:0] : _GEN_2007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3058 = 10'h1ae == _T_11 ? _ram_T_77[287:0] : _GEN_2008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3059 = 10'h1af == _T_11 ? _ram_T_77[287:0] : _GEN_2009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3060 = 10'h1b0 == _T_11 ? _ram_T_77[287:0] : _GEN_2010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3061 = 10'h1b1 == _T_11 ? _ram_T_77[287:0] : _GEN_2011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3062 = 10'h1b2 == _T_11 ? _ram_T_77[287:0] : _GEN_2012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3063 = 10'h1b3 == _T_11 ? _ram_T_77[287:0] : _GEN_2013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3064 = 10'h1b4 == _T_11 ? _ram_T_77[287:0] : _GEN_2014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3065 = 10'h1b5 == _T_11 ? _ram_T_77[287:0] : _GEN_2015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3066 = 10'h1b6 == _T_11 ? _ram_T_77[287:0] : _GEN_2016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3067 = 10'h1b7 == _T_11 ? _ram_T_77[287:0] : _GEN_2017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3068 = 10'h1b8 == _T_11 ? _ram_T_77[287:0] : _GEN_2018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3069 = 10'h1b9 == _T_11 ? _ram_T_77[287:0] : _GEN_2019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3070 = 10'h1ba == _T_11 ? _ram_T_77[287:0] : _GEN_2020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3071 = 10'h1bb == _T_11 ? _ram_T_77[287:0] : _GEN_2021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3072 = 10'h1bc == _T_11 ? _ram_T_77[287:0] : _GEN_2022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3073 = 10'h1bd == _T_11 ? _ram_T_77[287:0] : _GEN_2023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3074 = 10'h1be == _T_11 ? _ram_T_77[287:0] : _GEN_2024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3075 = 10'h1bf == _T_11 ? _ram_T_77[287:0] : _GEN_2025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3076 = 10'h1c0 == _T_11 ? _ram_T_77[287:0] : _GEN_2026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3077 = 10'h1c1 == _T_11 ? _ram_T_77[287:0] : _GEN_2027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3078 = 10'h1c2 == _T_11 ? _ram_T_77[287:0] : _GEN_2028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3079 = 10'h1c3 == _T_11 ? _ram_T_77[287:0] : _GEN_2029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3080 = 10'h1c4 == _T_11 ? _ram_T_77[287:0] : _GEN_2030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3081 = 10'h1c5 == _T_11 ? _ram_T_77[287:0] : _GEN_2031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3082 = 10'h1c6 == _T_11 ? _ram_T_77[287:0] : _GEN_2032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3083 = 10'h1c7 == _T_11 ? _ram_T_77[287:0] : _GEN_2033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3084 = 10'h1c8 == _T_11 ? _ram_T_77[287:0] : _GEN_2034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3085 = 10'h1c9 == _T_11 ? _ram_T_77[287:0] : _GEN_2035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3086 = 10'h1ca == _T_11 ? _ram_T_77[287:0] : _GEN_2036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3087 = 10'h1cb == _T_11 ? _ram_T_77[287:0] : _GEN_2037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3088 = 10'h1cc == _T_11 ? _ram_T_77[287:0] : _GEN_2038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3089 = 10'h1cd == _T_11 ? _ram_T_77[287:0] : _GEN_2039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3090 = 10'h1ce == _T_11 ? _ram_T_77[287:0] : _GEN_2040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3091 = 10'h1cf == _T_11 ? _ram_T_77[287:0] : _GEN_2041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3092 = 10'h1d0 == _T_11 ? _ram_T_77[287:0] : _GEN_2042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3093 = 10'h1d1 == _T_11 ? _ram_T_77[287:0] : _GEN_2043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3094 = 10'h1d2 == _T_11 ? _ram_T_77[287:0] : _GEN_2044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3095 = 10'h1d3 == _T_11 ? _ram_T_77[287:0] : _GEN_2045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3096 = 10'h1d4 == _T_11 ? _ram_T_77[287:0] : _GEN_2046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3097 = 10'h1d5 == _T_11 ? _ram_T_77[287:0] : _GEN_2047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3098 = 10'h1d6 == _T_11 ? _ram_T_77[287:0] : _GEN_2048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3099 = 10'h1d7 == _T_11 ? _ram_T_77[287:0] : _GEN_2049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3100 = 10'h1d8 == _T_11 ? _ram_T_77[287:0] : _GEN_2050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3101 = 10'h1d9 == _T_11 ? _ram_T_77[287:0] : _GEN_2051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3102 = 10'h1da == _T_11 ? _ram_T_77[287:0] : _GEN_2052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3103 = 10'h1db == _T_11 ? _ram_T_77[287:0] : _GEN_2053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3104 = 10'h1dc == _T_11 ? _ram_T_77[287:0] : _GEN_2054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3105 = 10'h1dd == _T_11 ? _ram_T_77[287:0] : _GEN_2055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3106 = 10'h1de == _T_11 ? _ram_T_77[287:0] : _GEN_2056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3107 = 10'h1df == _T_11 ? _ram_T_77[287:0] : _GEN_2057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3108 = 10'h1e0 == _T_11 ? _ram_T_77[287:0] : _GEN_2058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3109 = 10'h1e1 == _T_11 ? _ram_T_77[287:0] : _GEN_2059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3110 = 10'h1e2 == _T_11 ? _ram_T_77[287:0] : _GEN_2060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3111 = 10'h1e3 == _T_11 ? _ram_T_77[287:0] : _GEN_2061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3112 = 10'h1e4 == _T_11 ? _ram_T_77[287:0] : _GEN_2062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3113 = 10'h1e5 == _T_11 ? _ram_T_77[287:0] : _GEN_2063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3114 = 10'h1e6 == _T_11 ? _ram_T_77[287:0] : _GEN_2064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3115 = 10'h1e7 == _T_11 ? _ram_T_77[287:0] : _GEN_2065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3116 = 10'h1e8 == _T_11 ? _ram_T_77[287:0] : _GEN_2066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3117 = 10'h1e9 == _T_11 ? _ram_T_77[287:0] : _GEN_2067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3118 = 10'h1ea == _T_11 ? _ram_T_77[287:0] : _GEN_2068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3119 = 10'h1eb == _T_11 ? _ram_T_77[287:0] : _GEN_2069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3120 = 10'h1ec == _T_11 ? _ram_T_77[287:0] : _GEN_2070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3121 = 10'h1ed == _T_11 ? _ram_T_77[287:0] : _GEN_2071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3122 = 10'h1ee == _T_11 ? _ram_T_77[287:0] : _GEN_2072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3123 = 10'h1ef == _T_11 ? _ram_T_77[287:0] : _GEN_2073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3124 = 10'h1f0 == _T_11 ? _ram_T_77[287:0] : _GEN_2074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3125 = 10'h1f1 == _T_11 ? _ram_T_77[287:0] : _GEN_2075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3126 = 10'h1f2 == _T_11 ? _ram_T_77[287:0] : _GEN_2076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3127 = 10'h1f3 == _T_11 ? _ram_T_77[287:0] : _GEN_2077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3128 = 10'h1f4 == _T_11 ? _ram_T_77[287:0] : _GEN_2078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3129 = 10'h1f5 == _T_11 ? _ram_T_77[287:0] : _GEN_2079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3130 = 10'h1f6 == _T_11 ? _ram_T_77[287:0] : _GEN_2080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3131 = 10'h1f7 == _T_11 ? _ram_T_77[287:0] : _GEN_2081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3132 = 10'h1f8 == _T_11 ? _ram_T_77[287:0] : _GEN_2082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3133 = 10'h1f9 == _T_11 ? _ram_T_77[287:0] : _GEN_2083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3134 = 10'h1fa == _T_11 ? _ram_T_77[287:0] : _GEN_2084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3135 = 10'h1fb == _T_11 ? _ram_T_77[287:0] : _GEN_2085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3136 = 10'h1fc == _T_11 ? _ram_T_77[287:0] : _GEN_2086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3137 = 10'h1fd == _T_11 ? _ram_T_77[287:0] : _GEN_2087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3138 = 10'h1fe == _T_11 ? _ram_T_77[287:0] : _GEN_2088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3139 = 10'h1ff == _T_11 ? _ram_T_77[287:0] : _GEN_2089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3140 = 10'h200 == _T_11 ? _ram_T_77[287:0] : _GEN_2090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3141 = 10'h201 == _T_11 ? _ram_T_77[287:0] : _GEN_2091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3142 = 10'h202 == _T_11 ? _ram_T_77[287:0] : _GEN_2092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3143 = 10'h203 == _T_11 ? _ram_T_77[287:0] : _GEN_2093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3144 = 10'h204 == _T_11 ? _ram_T_77[287:0] : _GEN_2094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3145 = 10'h205 == _T_11 ? _ram_T_77[287:0] : _GEN_2095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3146 = 10'h206 == _T_11 ? _ram_T_77[287:0] : _GEN_2096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3147 = 10'h207 == _T_11 ? _ram_T_77[287:0] : _GEN_2097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3148 = 10'h208 == _T_11 ? _ram_T_77[287:0] : _GEN_2098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3149 = 10'h209 == _T_11 ? _ram_T_77[287:0] : _GEN_2099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3150 = 10'h20a == _T_11 ? _ram_T_77[287:0] : _GEN_2100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3151 = 10'h20b == _T_11 ? _ram_T_77[287:0] : _GEN_2101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3152 = 10'h20c == _T_11 ? _ram_T_77[287:0] : _GEN_2102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_13 = h + 10'h3; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_3 = vga_mem_ram_MPORT_27_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_3 = vga_mem_ram_MPORT_28_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_3 = vga_mem_ram_MPORT_29_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_3 = vga_mem_ram_MPORT_30_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_3 = vga_mem_ram_MPORT_31_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_3 = vga_mem_ram_MPORT_32_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_3 = vga_mem_ram_MPORT_33_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_3 = vga_mem_ram_MPORT_34_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_3 = vga_mem_ram_MPORT_35_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_98 = {278'h0,ram_hi_hi_hi_lo_3,ram_hi_hi_lo_3,ram_hi_lo_hi_3,ram_hi_lo_lo_3,ram_lo_hi_hi_hi_3,
    ram_lo_hi_hi_lo_3,ram_lo_hi_lo_3,ram_lo_lo_hi_3,ram_lo_lo_lo_3}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19066 = {{8191'd0}, _ram_T_98}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_102 = _GEN_19066 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_3154 = 10'h1 == _T_13 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3155 = 10'h2 == _T_13 ? ram_2 : _GEN_3154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3156 = 10'h3 == _T_13 ? ram_3 : _GEN_3155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3157 = 10'h4 == _T_13 ? ram_4 : _GEN_3156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3158 = 10'h5 == _T_13 ? ram_5 : _GEN_3157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3159 = 10'h6 == _T_13 ? ram_6 : _GEN_3158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3160 = 10'h7 == _T_13 ? ram_7 : _GEN_3159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3161 = 10'h8 == _T_13 ? ram_8 : _GEN_3160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3162 = 10'h9 == _T_13 ? ram_9 : _GEN_3161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3163 = 10'ha == _T_13 ? ram_10 : _GEN_3162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3164 = 10'hb == _T_13 ? ram_11 : _GEN_3163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3165 = 10'hc == _T_13 ? ram_12 : _GEN_3164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3166 = 10'hd == _T_13 ? ram_13 : _GEN_3165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3167 = 10'he == _T_13 ? ram_14 : _GEN_3166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3168 = 10'hf == _T_13 ? ram_15 : _GEN_3167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3169 = 10'h10 == _T_13 ? ram_16 : _GEN_3168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3170 = 10'h11 == _T_13 ? ram_17 : _GEN_3169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3171 = 10'h12 == _T_13 ? ram_18 : _GEN_3170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3172 = 10'h13 == _T_13 ? ram_19 : _GEN_3171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3173 = 10'h14 == _T_13 ? ram_20 : _GEN_3172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3174 = 10'h15 == _T_13 ? ram_21 : _GEN_3173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3175 = 10'h16 == _T_13 ? ram_22 : _GEN_3174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3176 = 10'h17 == _T_13 ? ram_23 : _GEN_3175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3177 = 10'h18 == _T_13 ? ram_24 : _GEN_3176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3178 = 10'h19 == _T_13 ? ram_25 : _GEN_3177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3179 = 10'h1a == _T_13 ? ram_26 : _GEN_3178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3180 = 10'h1b == _T_13 ? ram_27 : _GEN_3179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3181 = 10'h1c == _T_13 ? ram_28 : _GEN_3180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3182 = 10'h1d == _T_13 ? ram_29 : _GEN_3181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3183 = 10'h1e == _T_13 ? ram_30 : _GEN_3182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3184 = 10'h1f == _T_13 ? ram_31 : _GEN_3183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3185 = 10'h20 == _T_13 ? ram_32 : _GEN_3184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3186 = 10'h21 == _T_13 ? ram_33 : _GEN_3185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3187 = 10'h22 == _T_13 ? ram_34 : _GEN_3186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3188 = 10'h23 == _T_13 ? ram_35 : _GEN_3187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3189 = 10'h24 == _T_13 ? ram_36 : _GEN_3188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3190 = 10'h25 == _T_13 ? ram_37 : _GEN_3189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3191 = 10'h26 == _T_13 ? ram_38 : _GEN_3190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3192 = 10'h27 == _T_13 ? ram_39 : _GEN_3191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3193 = 10'h28 == _T_13 ? ram_40 : _GEN_3192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3194 = 10'h29 == _T_13 ? ram_41 : _GEN_3193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3195 = 10'h2a == _T_13 ? ram_42 : _GEN_3194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3196 = 10'h2b == _T_13 ? ram_43 : _GEN_3195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3197 = 10'h2c == _T_13 ? ram_44 : _GEN_3196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3198 = 10'h2d == _T_13 ? ram_45 : _GEN_3197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3199 = 10'h2e == _T_13 ? ram_46 : _GEN_3198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3200 = 10'h2f == _T_13 ? ram_47 : _GEN_3199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3201 = 10'h30 == _T_13 ? ram_48 : _GEN_3200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3202 = 10'h31 == _T_13 ? ram_49 : _GEN_3201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3203 = 10'h32 == _T_13 ? ram_50 : _GEN_3202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3204 = 10'h33 == _T_13 ? ram_51 : _GEN_3203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3205 = 10'h34 == _T_13 ? ram_52 : _GEN_3204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3206 = 10'h35 == _T_13 ? ram_53 : _GEN_3205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3207 = 10'h36 == _T_13 ? ram_54 : _GEN_3206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3208 = 10'h37 == _T_13 ? ram_55 : _GEN_3207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3209 = 10'h38 == _T_13 ? ram_56 : _GEN_3208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3210 = 10'h39 == _T_13 ? ram_57 : _GEN_3209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3211 = 10'h3a == _T_13 ? ram_58 : _GEN_3210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3212 = 10'h3b == _T_13 ? ram_59 : _GEN_3211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3213 = 10'h3c == _T_13 ? ram_60 : _GEN_3212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3214 = 10'h3d == _T_13 ? ram_61 : _GEN_3213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3215 = 10'h3e == _T_13 ? ram_62 : _GEN_3214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3216 = 10'h3f == _T_13 ? ram_63 : _GEN_3215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3217 = 10'h40 == _T_13 ? ram_64 : _GEN_3216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3218 = 10'h41 == _T_13 ? ram_65 : _GEN_3217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3219 = 10'h42 == _T_13 ? ram_66 : _GEN_3218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3220 = 10'h43 == _T_13 ? ram_67 : _GEN_3219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3221 = 10'h44 == _T_13 ? ram_68 : _GEN_3220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3222 = 10'h45 == _T_13 ? ram_69 : _GEN_3221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3223 = 10'h46 == _T_13 ? ram_70 : _GEN_3222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3224 = 10'h47 == _T_13 ? ram_71 : _GEN_3223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3225 = 10'h48 == _T_13 ? ram_72 : _GEN_3224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3226 = 10'h49 == _T_13 ? ram_73 : _GEN_3225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3227 = 10'h4a == _T_13 ? ram_74 : _GEN_3226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3228 = 10'h4b == _T_13 ? ram_75 : _GEN_3227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3229 = 10'h4c == _T_13 ? ram_76 : _GEN_3228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3230 = 10'h4d == _T_13 ? ram_77 : _GEN_3229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3231 = 10'h4e == _T_13 ? ram_78 : _GEN_3230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3232 = 10'h4f == _T_13 ? ram_79 : _GEN_3231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3233 = 10'h50 == _T_13 ? ram_80 : _GEN_3232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3234 = 10'h51 == _T_13 ? ram_81 : _GEN_3233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3235 = 10'h52 == _T_13 ? ram_82 : _GEN_3234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3236 = 10'h53 == _T_13 ? ram_83 : _GEN_3235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3237 = 10'h54 == _T_13 ? ram_84 : _GEN_3236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3238 = 10'h55 == _T_13 ? ram_85 : _GEN_3237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3239 = 10'h56 == _T_13 ? ram_86 : _GEN_3238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3240 = 10'h57 == _T_13 ? ram_87 : _GEN_3239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3241 = 10'h58 == _T_13 ? ram_88 : _GEN_3240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3242 = 10'h59 == _T_13 ? ram_89 : _GEN_3241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3243 = 10'h5a == _T_13 ? ram_90 : _GEN_3242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3244 = 10'h5b == _T_13 ? ram_91 : _GEN_3243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3245 = 10'h5c == _T_13 ? ram_92 : _GEN_3244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3246 = 10'h5d == _T_13 ? ram_93 : _GEN_3245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3247 = 10'h5e == _T_13 ? ram_94 : _GEN_3246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3248 = 10'h5f == _T_13 ? ram_95 : _GEN_3247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3249 = 10'h60 == _T_13 ? ram_96 : _GEN_3248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3250 = 10'h61 == _T_13 ? ram_97 : _GEN_3249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3251 = 10'h62 == _T_13 ? ram_98 : _GEN_3250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3252 = 10'h63 == _T_13 ? ram_99 : _GEN_3251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3253 = 10'h64 == _T_13 ? ram_100 : _GEN_3252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3254 = 10'h65 == _T_13 ? ram_101 : _GEN_3253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3255 = 10'h66 == _T_13 ? ram_102 : _GEN_3254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3256 = 10'h67 == _T_13 ? ram_103 : _GEN_3255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3257 = 10'h68 == _T_13 ? ram_104 : _GEN_3256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3258 = 10'h69 == _T_13 ? ram_105 : _GEN_3257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3259 = 10'h6a == _T_13 ? ram_106 : _GEN_3258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3260 = 10'h6b == _T_13 ? ram_107 : _GEN_3259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3261 = 10'h6c == _T_13 ? ram_108 : _GEN_3260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3262 = 10'h6d == _T_13 ? ram_109 : _GEN_3261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3263 = 10'h6e == _T_13 ? ram_110 : _GEN_3262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3264 = 10'h6f == _T_13 ? ram_111 : _GEN_3263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3265 = 10'h70 == _T_13 ? ram_112 : _GEN_3264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3266 = 10'h71 == _T_13 ? ram_113 : _GEN_3265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3267 = 10'h72 == _T_13 ? ram_114 : _GEN_3266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3268 = 10'h73 == _T_13 ? ram_115 : _GEN_3267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3269 = 10'h74 == _T_13 ? ram_116 : _GEN_3268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3270 = 10'h75 == _T_13 ? ram_117 : _GEN_3269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3271 = 10'h76 == _T_13 ? ram_118 : _GEN_3270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3272 = 10'h77 == _T_13 ? ram_119 : _GEN_3271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3273 = 10'h78 == _T_13 ? ram_120 : _GEN_3272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3274 = 10'h79 == _T_13 ? ram_121 : _GEN_3273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3275 = 10'h7a == _T_13 ? ram_122 : _GEN_3274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3276 = 10'h7b == _T_13 ? ram_123 : _GEN_3275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3277 = 10'h7c == _T_13 ? ram_124 : _GEN_3276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3278 = 10'h7d == _T_13 ? ram_125 : _GEN_3277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3279 = 10'h7e == _T_13 ? ram_126 : _GEN_3278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3280 = 10'h7f == _T_13 ? ram_127 : _GEN_3279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3281 = 10'h80 == _T_13 ? ram_128 : _GEN_3280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3282 = 10'h81 == _T_13 ? ram_129 : _GEN_3281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3283 = 10'h82 == _T_13 ? ram_130 : _GEN_3282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3284 = 10'h83 == _T_13 ? ram_131 : _GEN_3283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3285 = 10'h84 == _T_13 ? ram_132 : _GEN_3284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3286 = 10'h85 == _T_13 ? ram_133 : _GEN_3285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3287 = 10'h86 == _T_13 ? ram_134 : _GEN_3286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3288 = 10'h87 == _T_13 ? ram_135 : _GEN_3287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3289 = 10'h88 == _T_13 ? ram_136 : _GEN_3288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3290 = 10'h89 == _T_13 ? ram_137 : _GEN_3289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3291 = 10'h8a == _T_13 ? ram_138 : _GEN_3290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3292 = 10'h8b == _T_13 ? ram_139 : _GEN_3291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3293 = 10'h8c == _T_13 ? ram_140 : _GEN_3292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3294 = 10'h8d == _T_13 ? ram_141 : _GEN_3293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3295 = 10'h8e == _T_13 ? ram_142 : _GEN_3294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3296 = 10'h8f == _T_13 ? ram_143 : _GEN_3295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3297 = 10'h90 == _T_13 ? ram_144 : _GEN_3296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3298 = 10'h91 == _T_13 ? ram_145 : _GEN_3297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3299 = 10'h92 == _T_13 ? ram_146 : _GEN_3298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3300 = 10'h93 == _T_13 ? ram_147 : _GEN_3299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3301 = 10'h94 == _T_13 ? ram_148 : _GEN_3300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3302 = 10'h95 == _T_13 ? ram_149 : _GEN_3301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3303 = 10'h96 == _T_13 ? ram_150 : _GEN_3302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3304 = 10'h97 == _T_13 ? ram_151 : _GEN_3303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3305 = 10'h98 == _T_13 ? ram_152 : _GEN_3304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3306 = 10'h99 == _T_13 ? ram_153 : _GEN_3305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3307 = 10'h9a == _T_13 ? ram_154 : _GEN_3306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3308 = 10'h9b == _T_13 ? ram_155 : _GEN_3307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3309 = 10'h9c == _T_13 ? ram_156 : _GEN_3308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3310 = 10'h9d == _T_13 ? ram_157 : _GEN_3309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3311 = 10'h9e == _T_13 ? ram_158 : _GEN_3310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3312 = 10'h9f == _T_13 ? ram_159 : _GEN_3311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3313 = 10'ha0 == _T_13 ? ram_160 : _GEN_3312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3314 = 10'ha1 == _T_13 ? ram_161 : _GEN_3313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3315 = 10'ha2 == _T_13 ? ram_162 : _GEN_3314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3316 = 10'ha3 == _T_13 ? ram_163 : _GEN_3315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3317 = 10'ha4 == _T_13 ? ram_164 : _GEN_3316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3318 = 10'ha5 == _T_13 ? ram_165 : _GEN_3317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3319 = 10'ha6 == _T_13 ? ram_166 : _GEN_3318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3320 = 10'ha7 == _T_13 ? ram_167 : _GEN_3319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3321 = 10'ha8 == _T_13 ? ram_168 : _GEN_3320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3322 = 10'ha9 == _T_13 ? ram_169 : _GEN_3321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3323 = 10'haa == _T_13 ? ram_170 : _GEN_3322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3324 = 10'hab == _T_13 ? ram_171 : _GEN_3323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3325 = 10'hac == _T_13 ? ram_172 : _GEN_3324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3326 = 10'had == _T_13 ? ram_173 : _GEN_3325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3327 = 10'hae == _T_13 ? ram_174 : _GEN_3326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3328 = 10'haf == _T_13 ? ram_175 : _GEN_3327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3329 = 10'hb0 == _T_13 ? ram_176 : _GEN_3328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3330 = 10'hb1 == _T_13 ? ram_177 : _GEN_3329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3331 = 10'hb2 == _T_13 ? ram_178 : _GEN_3330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3332 = 10'hb3 == _T_13 ? ram_179 : _GEN_3331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3333 = 10'hb4 == _T_13 ? ram_180 : _GEN_3332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3334 = 10'hb5 == _T_13 ? ram_181 : _GEN_3333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3335 = 10'hb6 == _T_13 ? ram_182 : _GEN_3334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3336 = 10'hb7 == _T_13 ? ram_183 : _GEN_3335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3337 = 10'hb8 == _T_13 ? ram_184 : _GEN_3336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3338 = 10'hb9 == _T_13 ? ram_185 : _GEN_3337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3339 = 10'hba == _T_13 ? ram_186 : _GEN_3338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3340 = 10'hbb == _T_13 ? ram_187 : _GEN_3339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3341 = 10'hbc == _T_13 ? ram_188 : _GEN_3340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3342 = 10'hbd == _T_13 ? ram_189 : _GEN_3341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3343 = 10'hbe == _T_13 ? ram_190 : _GEN_3342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3344 = 10'hbf == _T_13 ? ram_191 : _GEN_3343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3345 = 10'hc0 == _T_13 ? ram_192 : _GEN_3344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3346 = 10'hc1 == _T_13 ? ram_193 : _GEN_3345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3347 = 10'hc2 == _T_13 ? ram_194 : _GEN_3346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3348 = 10'hc3 == _T_13 ? ram_195 : _GEN_3347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3349 = 10'hc4 == _T_13 ? ram_196 : _GEN_3348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3350 = 10'hc5 == _T_13 ? ram_197 : _GEN_3349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3351 = 10'hc6 == _T_13 ? ram_198 : _GEN_3350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3352 = 10'hc7 == _T_13 ? ram_199 : _GEN_3351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3353 = 10'hc8 == _T_13 ? ram_200 : _GEN_3352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3354 = 10'hc9 == _T_13 ? ram_201 : _GEN_3353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3355 = 10'hca == _T_13 ? ram_202 : _GEN_3354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3356 = 10'hcb == _T_13 ? ram_203 : _GEN_3355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3357 = 10'hcc == _T_13 ? ram_204 : _GEN_3356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3358 = 10'hcd == _T_13 ? ram_205 : _GEN_3357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3359 = 10'hce == _T_13 ? ram_206 : _GEN_3358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3360 = 10'hcf == _T_13 ? ram_207 : _GEN_3359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3361 = 10'hd0 == _T_13 ? ram_208 : _GEN_3360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3362 = 10'hd1 == _T_13 ? ram_209 : _GEN_3361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3363 = 10'hd2 == _T_13 ? ram_210 : _GEN_3362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3364 = 10'hd3 == _T_13 ? ram_211 : _GEN_3363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3365 = 10'hd4 == _T_13 ? ram_212 : _GEN_3364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3366 = 10'hd5 == _T_13 ? ram_213 : _GEN_3365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3367 = 10'hd6 == _T_13 ? ram_214 : _GEN_3366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3368 = 10'hd7 == _T_13 ? ram_215 : _GEN_3367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3369 = 10'hd8 == _T_13 ? ram_216 : _GEN_3368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3370 = 10'hd9 == _T_13 ? ram_217 : _GEN_3369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3371 = 10'hda == _T_13 ? ram_218 : _GEN_3370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3372 = 10'hdb == _T_13 ? ram_219 : _GEN_3371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3373 = 10'hdc == _T_13 ? ram_220 : _GEN_3372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3374 = 10'hdd == _T_13 ? ram_221 : _GEN_3373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3375 = 10'hde == _T_13 ? ram_222 : _GEN_3374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3376 = 10'hdf == _T_13 ? ram_223 : _GEN_3375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3377 = 10'he0 == _T_13 ? ram_224 : _GEN_3376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3378 = 10'he1 == _T_13 ? ram_225 : _GEN_3377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3379 = 10'he2 == _T_13 ? ram_226 : _GEN_3378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3380 = 10'he3 == _T_13 ? ram_227 : _GEN_3379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3381 = 10'he4 == _T_13 ? ram_228 : _GEN_3380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3382 = 10'he5 == _T_13 ? ram_229 : _GEN_3381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3383 = 10'he6 == _T_13 ? ram_230 : _GEN_3382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3384 = 10'he7 == _T_13 ? ram_231 : _GEN_3383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3385 = 10'he8 == _T_13 ? ram_232 : _GEN_3384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3386 = 10'he9 == _T_13 ? ram_233 : _GEN_3385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3387 = 10'hea == _T_13 ? ram_234 : _GEN_3386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3388 = 10'heb == _T_13 ? ram_235 : _GEN_3387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3389 = 10'hec == _T_13 ? ram_236 : _GEN_3388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3390 = 10'hed == _T_13 ? ram_237 : _GEN_3389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3391 = 10'hee == _T_13 ? ram_238 : _GEN_3390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3392 = 10'hef == _T_13 ? ram_239 : _GEN_3391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3393 = 10'hf0 == _T_13 ? ram_240 : _GEN_3392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3394 = 10'hf1 == _T_13 ? ram_241 : _GEN_3393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3395 = 10'hf2 == _T_13 ? ram_242 : _GEN_3394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3396 = 10'hf3 == _T_13 ? ram_243 : _GEN_3395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3397 = 10'hf4 == _T_13 ? ram_244 : _GEN_3396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3398 = 10'hf5 == _T_13 ? ram_245 : _GEN_3397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3399 = 10'hf6 == _T_13 ? ram_246 : _GEN_3398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3400 = 10'hf7 == _T_13 ? ram_247 : _GEN_3399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3401 = 10'hf8 == _T_13 ? ram_248 : _GEN_3400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3402 = 10'hf9 == _T_13 ? ram_249 : _GEN_3401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3403 = 10'hfa == _T_13 ? ram_250 : _GEN_3402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3404 = 10'hfb == _T_13 ? ram_251 : _GEN_3403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3405 = 10'hfc == _T_13 ? ram_252 : _GEN_3404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3406 = 10'hfd == _T_13 ? ram_253 : _GEN_3405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3407 = 10'hfe == _T_13 ? ram_254 : _GEN_3406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3408 = 10'hff == _T_13 ? ram_255 : _GEN_3407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3409 = 10'h100 == _T_13 ? ram_256 : _GEN_3408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3410 = 10'h101 == _T_13 ? ram_257 : _GEN_3409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3411 = 10'h102 == _T_13 ? ram_258 : _GEN_3410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3412 = 10'h103 == _T_13 ? ram_259 : _GEN_3411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3413 = 10'h104 == _T_13 ? ram_260 : _GEN_3412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3414 = 10'h105 == _T_13 ? ram_261 : _GEN_3413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3415 = 10'h106 == _T_13 ? ram_262 : _GEN_3414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3416 = 10'h107 == _T_13 ? ram_263 : _GEN_3415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3417 = 10'h108 == _T_13 ? ram_264 : _GEN_3416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3418 = 10'h109 == _T_13 ? ram_265 : _GEN_3417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3419 = 10'h10a == _T_13 ? ram_266 : _GEN_3418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3420 = 10'h10b == _T_13 ? ram_267 : _GEN_3419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3421 = 10'h10c == _T_13 ? ram_268 : _GEN_3420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3422 = 10'h10d == _T_13 ? ram_269 : _GEN_3421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3423 = 10'h10e == _T_13 ? ram_270 : _GEN_3422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3424 = 10'h10f == _T_13 ? ram_271 : _GEN_3423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3425 = 10'h110 == _T_13 ? ram_272 : _GEN_3424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3426 = 10'h111 == _T_13 ? ram_273 : _GEN_3425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3427 = 10'h112 == _T_13 ? ram_274 : _GEN_3426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3428 = 10'h113 == _T_13 ? ram_275 : _GEN_3427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3429 = 10'h114 == _T_13 ? ram_276 : _GEN_3428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3430 = 10'h115 == _T_13 ? ram_277 : _GEN_3429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3431 = 10'h116 == _T_13 ? ram_278 : _GEN_3430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3432 = 10'h117 == _T_13 ? ram_279 : _GEN_3431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3433 = 10'h118 == _T_13 ? ram_280 : _GEN_3432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3434 = 10'h119 == _T_13 ? ram_281 : _GEN_3433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3435 = 10'h11a == _T_13 ? ram_282 : _GEN_3434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3436 = 10'h11b == _T_13 ? ram_283 : _GEN_3435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3437 = 10'h11c == _T_13 ? ram_284 : _GEN_3436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3438 = 10'h11d == _T_13 ? ram_285 : _GEN_3437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3439 = 10'h11e == _T_13 ? ram_286 : _GEN_3438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3440 = 10'h11f == _T_13 ? ram_287 : _GEN_3439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3441 = 10'h120 == _T_13 ? ram_288 : _GEN_3440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3442 = 10'h121 == _T_13 ? ram_289 : _GEN_3441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3443 = 10'h122 == _T_13 ? ram_290 : _GEN_3442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3444 = 10'h123 == _T_13 ? ram_291 : _GEN_3443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3445 = 10'h124 == _T_13 ? ram_292 : _GEN_3444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3446 = 10'h125 == _T_13 ? ram_293 : _GEN_3445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3447 = 10'h126 == _T_13 ? ram_294 : _GEN_3446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3448 = 10'h127 == _T_13 ? ram_295 : _GEN_3447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3449 = 10'h128 == _T_13 ? ram_296 : _GEN_3448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3450 = 10'h129 == _T_13 ? ram_297 : _GEN_3449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3451 = 10'h12a == _T_13 ? ram_298 : _GEN_3450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3452 = 10'h12b == _T_13 ? ram_299 : _GEN_3451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3453 = 10'h12c == _T_13 ? ram_300 : _GEN_3452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3454 = 10'h12d == _T_13 ? ram_301 : _GEN_3453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3455 = 10'h12e == _T_13 ? ram_302 : _GEN_3454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3456 = 10'h12f == _T_13 ? ram_303 : _GEN_3455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3457 = 10'h130 == _T_13 ? ram_304 : _GEN_3456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3458 = 10'h131 == _T_13 ? ram_305 : _GEN_3457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3459 = 10'h132 == _T_13 ? ram_306 : _GEN_3458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3460 = 10'h133 == _T_13 ? ram_307 : _GEN_3459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3461 = 10'h134 == _T_13 ? ram_308 : _GEN_3460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3462 = 10'h135 == _T_13 ? ram_309 : _GEN_3461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3463 = 10'h136 == _T_13 ? ram_310 : _GEN_3462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3464 = 10'h137 == _T_13 ? ram_311 : _GEN_3463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3465 = 10'h138 == _T_13 ? ram_312 : _GEN_3464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3466 = 10'h139 == _T_13 ? ram_313 : _GEN_3465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3467 = 10'h13a == _T_13 ? ram_314 : _GEN_3466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3468 = 10'h13b == _T_13 ? ram_315 : _GEN_3467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3469 = 10'h13c == _T_13 ? ram_316 : _GEN_3468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3470 = 10'h13d == _T_13 ? ram_317 : _GEN_3469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3471 = 10'h13e == _T_13 ? ram_318 : _GEN_3470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3472 = 10'h13f == _T_13 ? ram_319 : _GEN_3471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3473 = 10'h140 == _T_13 ? ram_320 : _GEN_3472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3474 = 10'h141 == _T_13 ? ram_321 : _GEN_3473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3475 = 10'h142 == _T_13 ? ram_322 : _GEN_3474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3476 = 10'h143 == _T_13 ? ram_323 : _GEN_3475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3477 = 10'h144 == _T_13 ? ram_324 : _GEN_3476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3478 = 10'h145 == _T_13 ? ram_325 : _GEN_3477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3479 = 10'h146 == _T_13 ? ram_326 : _GEN_3478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3480 = 10'h147 == _T_13 ? ram_327 : _GEN_3479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3481 = 10'h148 == _T_13 ? ram_328 : _GEN_3480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3482 = 10'h149 == _T_13 ? ram_329 : _GEN_3481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3483 = 10'h14a == _T_13 ? ram_330 : _GEN_3482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3484 = 10'h14b == _T_13 ? ram_331 : _GEN_3483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3485 = 10'h14c == _T_13 ? ram_332 : _GEN_3484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3486 = 10'h14d == _T_13 ? ram_333 : _GEN_3485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3487 = 10'h14e == _T_13 ? ram_334 : _GEN_3486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3488 = 10'h14f == _T_13 ? ram_335 : _GEN_3487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3489 = 10'h150 == _T_13 ? ram_336 : _GEN_3488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3490 = 10'h151 == _T_13 ? ram_337 : _GEN_3489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3491 = 10'h152 == _T_13 ? ram_338 : _GEN_3490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3492 = 10'h153 == _T_13 ? ram_339 : _GEN_3491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3493 = 10'h154 == _T_13 ? ram_340 : _GEN_3492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3494 = 10'h155 == _T_13 ? ram_341 : _GEN_3493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3495 = 10'h156 == _T_13 ? ram_342 : _GEN_3494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3496 = 10'h157 == _T_13 ? ram_343 : _GEN_3495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3497 = 10'h158 == _T_13 ? ram_344 : _GEN_3496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3498 = 10'h159 == _T_13 ? ram_345 : _GEN_3497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3499 = 10'h15a == _T_13 ? ram_346 : _GEN_3498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3500 = 10'h15b == _T_13 ? ram_347 : _GEN_3499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3501 = 10'h15c == _T_13 ? ram_348 : _GEN_3500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3502 = 10'h15d == _T_13 ? ram_349 : _GEN_3501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3503 = 10'h15e == _T_13 ? ram_350 : _GEN_3502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3504 = 10'h15f == _T_13 ? ram_351 : _GEN_3503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3505 = 10'h160 == _T_13 ? ram_352 : _GEN_3504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3506 = 10'h161 == _T_13 ? ram_353 : _GEN_3505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3507 = 10'h162 == _T_13 ? ram_354 : _GEN_3506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3508 = 10'h163 == _T_13 ? ram_355 : _GEN_3507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3509 = 10'h164 == _T_13 ? ram_356 : _GEN_3508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3510 = 10'h165 == _T_13 ? ram_357 : _GEN_3509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3511 = 10'h166 == _T_13 ? ram_358 : _GEN_3510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3512 = 10'h167 == _T_13 ? ram_359 : _GEN_3511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3513 = 10'h168 == _T_13 ? ram_360 : _GEN_3512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3514 = 10'h169 == _T_13 ? ram_361 : _GEN_3513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3515 = 10'h16a == _T_13 ? ram_362 : _GEN_3514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3516 = 10'h16b == _T_13 ? ram_363 : _GEN_3515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3517 = 10'h16c == _T_13 ? ram_364 : _GEN_3516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3518 = 10'h16d == _T_13 ? ram_365 : _GEN_3517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3519 = 10'h16e == _T_13 ? ram_366 : _GEN_3518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3520 = 10'h16f == _T_13 ? ram_367 : _GEN_3519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3521 = 10'h170 == _T_13 ? ram_368 : _GEN_3520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3522 = 10'h171 == _T_13 ? ram_369 : _GEN_3521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3523 = 10'h172 == _T_13 ? ram_370 : _GEN_3522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3524 = 10'h173 == _T_13 ? ram_371 : _GEN_3523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3525 = 10'h174 == _T_13 ? ram_372 : _GEN_3524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3526 = 10'h175 == _T_13 ? ram_373 : _GEN_3525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3527 = 10'h176 == _T_13 ? ram_374 : _GEN_3526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3528 = 10'h177 == _T_13 ? ram_375 : _GEN_3527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3529 = 10'h178 == _T_13 ? ram_376 : _GEN_3528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3530 = 10'h179 == _T_13 ? ram_377 : _GEN_3529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3531 = 10'h17a == _T_13 ? ram_378 : _GEN_3530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3532 = 10'h17b == _T_13 ? ram_379 : _GEN_3531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3533 = 10'h17c == _T_13 ? ram_380 : _GEN_3532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3534 = 10'h17d == _T_13 ? ram_381 : _GEN_3533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3535 = 10'h17e == _T_13 ? ram_382 : _GEN_3534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3536 = 10'h17f == _T_13 ? ram_383 : _GEN_3535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3537 = 10'h180 == _T_13 ? ram_384 : _GEN_3536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3538 = 10'h181 == _T_13 ? ram_385 : _GEN_3537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3539 = 10'h182 == _T_13 ? ram_386 : _GEN_3538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3540 = 10'h183 == _T_13 ? ram_387 : _GEN_3539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3541 = 10'h184 == _T_13 ? ram_388 : _GEN_3540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3542 = 10'h185 == _T_13 ? ram_389 : _GEN_3541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3543 = 10'h186 == _T_13 ? ram_390 : _GEN_3542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3544 = 10'h187 == _T_13 ? ram_391 : _GEN_3543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3545 = 10'h188 == _T_13 ? ram_392 : _GEN_3544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3546 = 10'h189 == _T_13 ? ram_393 : _GEN_3545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3547 = 10'h18a == _T_13 ? ram_394 : _GEN_3546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3548 = 10'h18b == _T_13 ? ram_395 : _GEN_3547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3549 = 10'h18c == _T_13 ? ram_396 : _GEN_3548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3550 = 10'h18d == _T_13 ? ram_397 : _GEN_3549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3551 = 10'h18e == _T_13 ? ram_398 : _GEN_3550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3552 = 10'h18f == _T_13 ? ram_399 : _GEN_3551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3553 = 10'h190 == _T_13 ? ram_400 : _GEN_3552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3554 = 10'h191 == _T_13 ? ram_401 : _GEN_3553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3555 = 10'h192 == _T_13 ? ram_402 : _GEN_3554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3556 = 10'h193 == _T_13 ? ram_403 : _GEN_3555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3557 = 10'h194 == _T_13 ? ram_404 : _GEN_3556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3558 = 10'h195 == _T_13 ? ram_405 : _GEN_3557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3559 = 10'h196 == _T_13 ? ram_406 : _GEN_3558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3560 = 10'h197 == _T_13 ? ram_407 : _GEN_3559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3561 = 10'h198 == _T_13 ? ram_408 : _GEN_3560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3562 = 10'h199 == _T_13 ? ram_409 : _GEN_3561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3563 = 10'h19a == _T_13 ? ram_410 : _GEN_3562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3564 = 10'h19b == _T_13 ? ram_411 : _GEN_3563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3565 = 10'h19c == _T_13 ? ram_412 : _GEN_3564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3566 = 10'h19d == _T_13 ? ram_413 : _GEN_3565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3567 = 10'h19e == _T_13 ? ram_414 : _GEN_3566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3568 = 10'h19f == _T_13 ? ram_415 : _GEN_3567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3569 = 10'h1a0 == _T_13 ? ram_416 : _GEN_3568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3570 = 10'h1a1 == _T_13 ? ram_417 : _GEN_3569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3571 = 10'h1a2 == _T_13 ? ram_418 : _GEN_3570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3572 = 10'h1a3 == _T_13 ? ram_419 : _GEN_3571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3573 = 10'h1a4 == _T_13 ? ram_420 : _GEN_3572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3574 = 10'h1a5 == _T_13 ? ram_421 : _GEN_3573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3575 = 10'h1a6 == _T_13 ? ram_422 : _GEN_3574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3576 = 10'h1a7 == _T_13 ? ram_423 : _GEN_3575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3577 = 10'h1a8 == _T_13 ? ram_424 : _GEN_3576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3578 = 10'h1a9 == _T_13 ? ram_425 : _GEN_3577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3579 = 10'h1aa == _T_13 ? ram_426 : _GEN_3578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3580 = 10'h1ab == _T_13 ? ram_427 : _GEN_3579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3581 = 10'h1ac == _T_13 ? ram_428 : _GEN_3580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3582 = 10'h1ad == _T_13 ? ram_429 : _GEN_3581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3583 = 10'h1ae == _T_13 ? ram_430 : _GEN_3582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3584 = 10'h1af == _T_13 ? ram_431 : _GEN_3583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3585 = 10'h1b0 == _T_13 ? ram_432 : _GEN_3584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3586 = 10'h1b1 == _T_13 ? ram_433 : _GEN_3585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3587 = 10'h1b2 == _T_13 ? ram_434 : _GEN_3586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3588 = 10'h1b3 == _T_13 ? ram_435 : _GEN_3587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3589 = 10'h1b4 == _T_13 ? ram_436 : _GEN_3588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3590 = 10'h1b5 == _T_13 ? ram_437 : _GEN_3589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3591 = 10'h1b6 == _T_13 ? ram_438 : _GEN_3590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3592 = 10'h1b7 == _T_13 ? ram_439 : _GEN_3591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3593 = 10'h1b8 == _T_13 ? ram_440 : _GEN_3592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3594 = 10'h1b9 == _T_13 ? ram_441 : _GEN_3593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3595 = 10'h1ba == _T_13 ? ram_442 : _GEN_3594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3596 = 10'h1bb == _T_13 ? ram_443 : _GEN_3595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3597 = 10'h1bc == _T_13 ? ram_444 : _GEN_3596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3598 = 10'h1bd == _T_13 ? ram_445 : _GEN_3597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3599 = 10'h1be == _T_13 ? ram_446 : _GEN_3598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3600 = 10'h1bf == _T_13 ? ram_447 : _GEN_3599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3601 = 10'h1c0 == _T_13 ? ram_448 : _GEN_3600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3602 = 10'h1c1 == _T_13 ? ram_449 : _GEN_3601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3603 = 10'h1c2 == _T_13 ? ram_450 : _GEN_3602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3604 = 10'h1c3 == _T_13 ? ram_451 : _GEN_3603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3605 = 10'h1c4 == _T_13 ? ram_452 : _GEN_3604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3606 = 10'h1c5 == _T_13 ? ram_453 : _GEN_3605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3607 = 10'h1c6 == _T_13 ? ram_454 : _GEN_3606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3608 = 10'h1c7 == _T_13 ? ram_455 : _GEN_3607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3609 = 10'h1c8 == _T_13 ? ram_456 : _GEN_3608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3610 = 10'h1c9 == _T_13 ? ram_457 : _GEN_3609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3611 = 10'h1ca == _T_13 ? ram_458 : _GEN_3610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3612 = 10'h1cb == _T_13 ? ram_459 : _GEN_3611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3613 = 10'h1cc == _T_13 ? ram_460 : _GEN_3612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3614 = 10'h1cd == _T_13 ? ram_461 : _GEN_3613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3615 = 10'h1ce == _T_13 ? ram_462 : _GEN_3614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3616 = 10'h1cf == _T_13 ? ram_463 : _GEN_3615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3617 = 10'h1d0 == _T_13 ? ram_464 : _GEN_3616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3618 = 10'h1d1 == _T_13 ? ram_465 : _GEN_3617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3619 = 10'h1d2 == _T_13 ? ram_466 : _GEN_3618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3620 = 10'h1d3 == _T_13 ? ram_467 : _GEN_3619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3621 = 10'h1d4 == _T_13 ? ram_468 : _GEN_3620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3622 = 10'h1d5 == _T_13 ? ram_469 : _GEN_3621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3623 = 10'h1d6 == _T_13 ? ram_470 : _GEN_3622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3624 = 10'h1d7 == _T_13 ? ram_471 : _GEN_3623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3625 = 10'h1d8 == _T_13 ? ram_472 : _GEN_3624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3626 = 10'h1d9 == _T_13 ? ram_473 : _GEN_3625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3627 = 10'h1da == _T_13 ? ram_474 : _GEN_3626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3628 = 10'h1db == _T_13 ? ram_475 : _GEN_3627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3629 = 10'h1dc == _T_13 ? ram_476 : _GEN_3628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3630 = 10'h1dd == _T_13 ? ram_477 : _GEN_3629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3631 = 10'h1de == _T_13 ? ram_478 : _GEN_3630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3632 = 10'h1df == _T_13 ? ram_479 : _GEN_3631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3633 = 10'h1e0 == _T_13 ? ram_480 : _GEN_3632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3634 = 10'h1e1 == _T_13 ? ram_481 : _GEN_3633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3635 = 10'h1e2 == _T_13 ? ram_482 : _GEN_3634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3636 = 10'h1e3 == _T_13 ? ram_483 : _GEN_3635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3637 = 10'h1e4 == _T_13 ? ram_484 : _GEN_3636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3638 = 10'h1e5 == _T_13 ? ram_485 : _GEN_3637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3639 = 10'h1e6 == _T_13 ? ram_486 : _GEN_3638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3640 = 10'h1e7 == _T_13 ? ram_487 : _GEN_3639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3641 = 10'h1e8 == _T_13 ? ram_488 : _GEN_3640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3642 = 10'h1e9 == _T_13 ? ram_489 : _GEN_3641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3643 = 10'h1ea == _T_13 ? ram_490 : _GEN_3642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3644 = 10'h1eb == _T_13 ? ram_491 : _GEN_3643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3645 = 10'h1ec == _T_13 ? ram_492 : _GEN_3644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3646 = 10'h1ed == _T_13 ? ram_493 : _GEN_3645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3647 = 10'h1ee == _T_13 ? ram_494 : _GEN_3646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3648 = 10'h1ef == _T_13 ? ram_495 : _GEN_3647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3649 = 10'h1f0 == _T_13 ? ram_496 : _GEN_3648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3650 = 10'h1f1 == _T_13 ? ram_497 : _GEN_3649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3651 = 10'h1f2 == _T_13 ? ram_498 : _GEN_3650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3652 = 10'h1f3 == _T_13 ? ram_499 : _GEN_3651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3653 = 10'h1f4 == _T_13 ? ram_500 : _GEN_3652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3654 = 10'h1f5 == _T_13 ? ram_501 : _GEN_3653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3655 = 10'h1f6 == _T_13 ? ram_502 : _GEN_3654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3656 = 10'h1f7 == _T_13 ? ram_503 : _GEN_3655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3657 = 10'h1f8 == _T_13 ? ram_504 : _GEN_3656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3658 = 10'h1f9 == _T_13 ? ram_505 : _GEN_3657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3659 = 10'h1fa == _T_13 ? ram_506 : _GEN_3658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3660 = 10'h1fb == _T_13 ? ram_507 : _GEN_3659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3661 = 10'h1fc == _T_13 ? ram_508 : _GEN_3660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3662 = 10'h1fd == _T_13 ? ram_509 : _GEN_3661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3663 = 10'h1fe == _T_13 ? ram_510 : _GEN_3662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3664 = 10'h1ff == _T_13 ? ram_511 : _GEN_3663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3665 = 10'h200 == _T_13 ? ram_512 : _GEN_3664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3666 = 10'h201 == _T_13 ? ram_513 : _GEN_3665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3667 = 10'h202 == _T_13 ? ram_514 : _GEN_3666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3668 = 10'h203 == _T_13 ? ram_515 : _GEN_3667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3669 = 10'h204 == _T_13 ? ram_516 : _GEN_3668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3670 = 10'h205 == _T_13 ? ram_517 : _GEN_3669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3671 = 10'h206 == _T_13 ? ram_518 : _GEN_3670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3672 = 10'h207 == _T_13 ? ram_519 : _GEN_3671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3673 = 10'h208 == _T_13 ? ram_520 : _GEN_3672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3674 = 10'h209 == _T_13 ? ram_521 : _GEN_3673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3675 = 10'h20a == _T_13 ? ram_522 : _GEN_3674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3676 = 10'h20b == _T_13 ? ram_523 : _GEN_3675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_3677 = 10'h20c == _T_13 ? ram_524 : _GEN_3676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19067 = {{8190'd0}, _GEN_3677}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_103 = _GEN_19067 ^ _ram_T_102; // @[vga.scala 64:41]
  wire [287:0] _GEN_3678 = 10'h0 == _T_13 ? _ram_T_103[287:0] : _GEN_2628; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3679 = 10'h1 == _T_13 ? _ram_T_103[287:0] : _GEN_2629; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3680 = 10'h2 == _T_13 ? _ram_T_103[287:0] : _GEN_2630; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3681 = 10'h3 == _T_13 ? _ram_T_103[287:0] : _GEN_2631; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3682 = 10'h4 == _T_13 ? _ram_T_103[287:0] : _GEN_2632; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3683 = 10'h5 == _T_13 ? _ram_T_103[287:0] : _GEN_2633; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3684 = 10'h6 == _T_13 ? _ram_T_103[287:0] : _GEN_2634; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3685 = 10'h7 == _T_13 ? _ram_T_103[287:0] : _GEN_2635; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3686 = 10'h8 == _T_13 ? _ram_T_103[287:0] : _GEN_2636; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3687 = 10'h9 == _T_13 ? _ram_T_103[287:0] : _GEN_2637; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3688 = 10'ha == _T_13 ? _ram_T_103[287:0] : _GEN_2638; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3689 = 10'hb == _T_13 ? _ram_T_103[287:0] : _GEN_2639; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3690 = 10'hc == _T_13 ? _ram_T_103[287:0] : _GEN_2640; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3691 = 10'hd == _T_13 ? _ram_T_103[287:0] : _GEN_2641; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3692 = 10'he == _T_13 ? _ram_T_103[287:0] : _GEN_2642; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3693 = 10'hf == _T_13 ? _ram_T_103[287:0] : _GEN_2643; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3694 = 10'h10 == _T_13 ? _ram_T_103[287:0] : _GEN_2644; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3695 = 10'h11 == _T_13 ? _ram_T_103[287:0] : _GEN_2645; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3696 = 10'h12 == _T_13 ? _ram_T_103[287:0] : _GEN_2646; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3697 = 10'h13 == _T_13 ? _ram_T_103[287:0] : _GEN_2647; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3698 = 10'h14 == _T_13 ? _ram_T_103[287:0] : _GEN_2648; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3699 = 10'h15 == _T_13 ? _ram_T_103[287:0] : _GEN_2649; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3700 = 10'h16 == _T_13 ? _ram_T_103[287:0] : _GEN_2650; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3701 = 10'h17 == _T_13 ? _ram_T_103[287:0] : _GEN_2651; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3702 = 10'h18 == _T_13 ? _ram_T_103[287:0] : _GEN_2652; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3703 = 10'h19 == _T_13 ? _ram_T_103[287:0] : _GEN_2653; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3704 = 10'h1a == _T_13 ? _ram_T_103[287:0] : _GEN_2654; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3705 = 10'h1b == _T_13 ? _ram_T_103[287:0] : _GEN_2655; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3706 = 10'h1c == _T_13 ? _ram_T_103[287:0] : _GEN_2656; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3707 = 10'h1d == _T_13 ? _ram_T_103[287:0] : _GEN_2657; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3708 = 10'h1e == _T_13 ? _ram_T_103[287:0] : _GEN_2658; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3709 = 10'h1f == _T_13 ? _ram_T_103[287:0] : _GEN_2659; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3710 = 10'h20 == _T_13 ? _ram_T_103[287:0] : _GEN_2660; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3711 = 10'h21 == _T_13 ? _ram_T_103[287:0] : _GEN_2661; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3712 = 10'h22 == _T_13 ? _ram_T_103[287:0] : _GEN_2662; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3713 = 10'h23 == _T_13 ? _ram_T_103[287:0] : _GEN_2663; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3714 = 10'h24 == _T_13 ? _ram_T_103[287:0] : _GEN_2664; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3715 = 10'h25 == _T_13 ? _ram_T_103[287:0] : _GEN_2665; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3716 = 10'h26 == _T_13 ? _ram_T_103[287:0] : _GEN_2666; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3717 = 10'h27 == _T_13 ? _ram_T_103[287:0] : _GEN_2667; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3718 = 10'h28 == _T_13 ? _ram_T_103[287:0] : _GEN_2668; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3719 = 10'h29 == _T_13 ? _ram_T_103[287:0] : _GEN_2669; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3720 = 10'h2a == _T_13 ? _ram_T_103[287:0] : _GEN_2670; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3721 = 10'h2b == _T_13 ? _ram_T_103[287:0] : _GEN_2671; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3722 = 10'h2c == _T_13 ? _ram_T_103[287:0] : _GEN_2672; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3723 = 10'h2d == _T_13 ? _ram_T_103[287:0] : _GEN_2673; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3724 = 10'h2e == _T_13 ? _ram_T_103[287:0] : _GEN_2674; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3725 = 10'h2f == _T_13 ? _ram_T_103[287:0] : _GEN_2675; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3726 = 10'h30 == _T_13 ? _ram_T_103[287:0] : _GEN_2676; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3727 = 10'h31 == _T_13 ? _ram_T_103[287:0] : _GEN_2677; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3728 = 10'h32 == _T_13 ? _ram_T_103[287:0] : _GEN_2678; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3729 = 10'h33 == _T_13 ? _ram_T_103[287:0] : _GEN_2679; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3730 = 10'h34 == _T_13 ? _ram_T_103[287:0] : _GEN_2680; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3731 = 10'h35 == _T_13 ? _ram_T_103[287:0] : _GEN_2681; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3732 = 10'h36 == _T_13 ? _ram_T_103[287:0] : _GEN_2682; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3733 = 10'h37 == _T_13 ? _ram_T_103[287:0] : _GEN_2683; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3734 = 10'h38 == _T_13 ? _ram_T_103[287:0] : _GEN_2684; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3735 = 10'h39 == _T_13 ? _ram_T_103[287:0] : _GEN_2685; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3736 = 10'h3a == _T_13 ? _ram_T_103[287:0] : _GEN_2686; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3737 = 10'h3b == _T_13 ? _ram_T_103[287:0] : _GEN_2687; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3738 = 10'h3c == _T_13 ? _ram_T_103[287:0] : _GEN_2688; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3739 = 10'h3d == _T_13 ? _ram_T_103[287:0] : _GEN_2689; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3740 = 10'h3e == _T_13 ? _ram_T_103[287:0] : _GEN_2690; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3741 = 10'h3f == _T_13 ? _ram_T_103[287:0] : _GEN_2691; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3742 = 10'h40 == _T_13 ? _ram_T_103[287:0] : _GEN_2692; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3743 = 10'h41 == _T_13 ? _ram_T_103[287:0] : _GEN_2693; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3744 = 10'h42 == _T_13 ? _ram_T_103[287:0] : _GEN_2694; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3745 = 10'h43 == _T_13 ? _ram_T_103[287:0] : _GEN_2695; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3746 = 10'h44 == _T_13 ? _ram_T_103[287:0] : _GEN_2696; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3747 = 10'h45 == _T_13 ? _ram_T_103[287:0] : _GEN_2697; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3748 = 10'h46 == _T_13 ? _ram_T_103[287:0] : _GEN_2698; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3749 = 10'h47 == _T_13 ? _ram_T_103[287:0] : _GEN_2699; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3750 = 10'h48 == _T_13 ? _ram_T_103[287:0] : _GEN_2700; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3751 = 10'h49 == _T_13 ? _ram_T_103[287:0] : _GEN_2701; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3752 = 10'h4a == _T_13 ? _ram_T_103[287:0] : _GEN_2702; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3753 = 10'h4b == _T_13 ? _ram_T_103[287:0] : _GEN_2703; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3754 = 10'h4c == _T_13 ? _ram_T_103[287:0] : _GEN_2704; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3755 = 10'h4d == _T_13 ? _ram_T_103[287:0] : _GEN_2705; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3756 = 10'h4e == _T_13 ? _ram_T_103[287:0] : _GEN_2706; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3757 = 10'h4f == _T_13 ? _ram_T_103[287:0] : _GEN_2707; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3758 = 10'h50 == _T_13 ? _ram_T_103[287:0] : _GEN_2708; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3759 = 10'h51 == _T_13 ? _ram_T_103[287:0] : _GEN_2709; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3760 = 10'h52 == _T_13 ? _ram_T_103[287:0] : _GEN_2710; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3761 = 10'h53 == _T_13 ? _ram_T_103[287:0] : _GEN_2711; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3762 = 10'h54 == _T_13 ? _ram_T_103[287:0] : _GEN_2712; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3763 = 10'h55 == _T_13 ? _ram_T_103[287:0] : _GEN_2713; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3764 = 10'h56 == _T_13 ? _ram_T_103[287:0] : _GEN_2714; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3765 = 10'h57 == _T_13 ? _ram_T_103[287:0] : _GEN_2715; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3766 = 10'h58 == _T_13 ? _ram_T_103[287:0] : _GEN_2716; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3767 = 10'h59 == _T_13 ? _ram_T_103[287:0] : _GEN_2717; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3768 = 10'h5a == _T_13 ? _ram_T_103[287:0] : _GEN_2718; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3769 = 10'h5b == _T_13 ? _ram_T_103[287:0] : _GEN_2719; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3770 = 10'h5c == _T_13 ? _ram_T_103[287:0] : _GEN_2720; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3771 = 10'h5d == _T_13 ? _ram_T_103[287:0] : _GEN_2721; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3772 = 10'h5e == _T_13 ? _ram_T_103[287:0] : _GEN_2722; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3773 = 10'h5f == _T_13 ? _ram_T_103[287:0] : _GEN_2723; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3774 = 10'h60 == _T_13 ? _ram_T_103[287:0] : _GEN_2724; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3775 = 10'h61 == _T_13 ? _ram_T_103[287:0] : _GEN_2725; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3776 = 10'h62 == _T_13 ? _ram_T_103[287:0] : _GEN_2726; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3777 = 10'h63 == _T_13 ? _ram_T_103[287:0] : _GEN_2727; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3778 = 10'h64 == _T_13 ? _ram_T_103[287:0] : _GEN_2728; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3779 = 10'h65 == _T_13 ? _ram_T_103[287:0] : _GEN_2729; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3780 = 10'h66 == _T_13 ? _ram_T_103[287:0] : _GEN_2730; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3781 = 10'h67 == _T_13 ? _ram_T_103[287:0] : _GEN_2731; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3782 = 10'h68 == _T_13 ? _ram_T_103[287:0] : _GEN_2732; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3783 = 10'h69 == _T_13 ? _ram_T_103[287:0] : _GEN_2733; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3784 = 10'h6a == _T_13 ? _ram_T_103[287:0] : _GEN_2734; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3785 = 10'h6b == _T_13 ? _ram_T_103[287:0] : _GEN_2735; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3786 = 10'h6c == _T_13 ? _ram_T_103[287:0] : _GEN_2736; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3787 = 10'h6d == _T_13 ? _ram_T_103[287:0] : _GEN_2737; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3788 = 10'h6e == _T_13 ? _ram_T_103[287:0] : _GEN_2738; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3789 = 10'h6f == _T_13 ? _ram_T_103[287:0] : _GEN_2739; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3790 = 10'h70 == _T_13 ? _ram_T_103[287:0] : _GEN_2740; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3791 = 10'h71 == _T_13 ? _ram_T_103[287:0] : _GEN_2741; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3792 = 10'h72 == _T_13 ? _ram_T_103[287:0] : _GEN_2742; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3793 = 10'h73 == _T_13 ? _ram_T_103[287:0] : _GEN_2743; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3794 = 10'h74 == _T_13 ? _ram_T_103[287:0] : _GEN_2744; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3795 = 10'h75 == _T_13 ? _ram_T_103[287:0] : _GEN_2745; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3796 = 10'h76 == _T_13 ? _ram_T_103[287:0] : _GEN_2746; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3797 = 10'h77 == _T_13 ? _ram_T_103[287:0] : _GEN_2747; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3798 = 10'h78 == _T_13 ? _ram_T_103[287:0] : _GEN_2748; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3799 = 10'h79 == _T_13 ? _ram_T_103[287:0] : _GEN_2749; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3800 = 10'h7a == _T_13 ? _ram_T_103[287:0] : _GEN_2750; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3801 = 10'h7b == _T_13 ? _ram_T_103[287:0] : _GEN_2751; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3802 = 10'h7c == _T_13 ? _ram_T_103[287:0] : _GEN_2752; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3803 = 10'h7d == _T_13 ? _ram_T_103[287:0] : _GEN_2753; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3804 = 10'h7e == _T_13 ? _ram_T_103[287:0] : _GEN_2754; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3805 = 10'h7f == _T_13 ? _ram_T_103[287:0] : _GEN_2755; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3806 = 10'h80 == _T_13 ? _ram_T_103[287:0] : _GEN_2756; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3807 = 10'h81 == _T_13 ? _ram_T_103[287:0] : _GEN_2757; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3808 = 10'h82 == _T_13 ? _ram_T_103[287:0] : _GEN_2758; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3809 = 10'h83 == _T_13 ? _ram_T_103[287:0] : _GEN_2759; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3810 = 10'h84 == _T_13 ? _ram_T_103[287:0] : _GEN_2760; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3811 = 10'h85 == _T_13 ? _ram_T_103[287:0] : _GEN_2761; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3812 = 10'h86 == _T_13 ? _ram_T_103[287:0] : _GEN_2762; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3813 = 10'h87 == _T_13 ? _ram_T_103[287:0] : _GEN_2763; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3814 = 10'h88 == _T_13 ? _ram_T_103[287:0] : _GEN_2764; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3815 = 10'h89 == _T_13 ? _ram_T_103[287:0] : _GEN_2765; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3816 = 10'h8a == _T_13 ? _ram_T_103[287:0] : _GEN_2766; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3817 = 10'h8b == _T_13 ? _ram_T_103[287:0] : _GEN_2767; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3818 = 10'h8c == _T_13 ? _ram_T_103[287:0] : _GEN_2768; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3819 = 10'h8d == _T_13 ? _ram_T_103[287:0] : _GEN_2769; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3820 = 10'h8e == _T_13 ? _ram_T_103[287:0] : _GEN_2770; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3821 = 10'h8f == _T_13 ? _ram_T_103[287:0] : _GEN_2771; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3822 = 10'h90 == _T_13 ? _ram_T_103[287:0] : _GEN_2772; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3823 = 10'h91 == _T_13 ? _ram_T_103[287:0] : _GEN_2773; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3824 = 10'h92 == _T_13 ? _ram_T_103[287:0] : _GEN_2774; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3825 = 10'h93 == _T_13 ? _ram_T_103[287:0] : _GEN_2775; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3826 = 10'h94 == _T_13 ? _ram_T_103[287:0] : _GEN_2776; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3827 = 10'h95 == _T_13 ? _ram_T_103[287:0] : _GEN_2777; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3828 = 10'h96 == _T_13 ? _ram_T_103[287:0] : _GEN_2778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3829 = 10'h97 == _T_13 ? _ram_T_103[287:0] : _GEN_2779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3830 = 10'h98 == _T_13 ? _ram_T_103[287:0] : _GEN_2780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3831 = 10'h99 == _T_13 ? _ram_T_103[287:0] : _GEN_2781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3832 = 10'h9a == _T_13 ? _ram_T_103[287:0] : _GEN_2782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3833 = 10'h9b == _T_13 ? _ram_T_103[287:0] : _GEN_2783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3834 = 10'h9c == _T_13 ? _ram_T_103[287:0] : _GEN_2784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3835 = 10'h9d == _T_13 ? _ram_T_103[287:0] : _GEN_2785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3836 = 10'h9e == _T_13 ? _ram_T_103[287:0] : _GEN_2786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3837 = 10'h9f == _T_13 ? _ram_T_103[287:0] : _GEN_2787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3838 = 10'ha0 == _T_13 ? _ram_T_103[287:0] : _GEN_2788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3839 = 10'ha1 == _T_13 ? _ram_T_103[287:0] : _GEN_2789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3840 = 10'ha2 == _T_13 ? _ram_T_103[287:0] : _GEN_2790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3841 = 10'ha3 == _T_13 ? _ram_T_103[287:0] : _GEN_2791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3842 = 10'ha4 == _T_13 ? _ram_T_103[287:0] : _GEN_2792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3843 = 10'ha5 == _T_13 ? _ram_T_103[287:0] : _GEN_2793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3844 = 10'ha6 == _T_13 ? _ram_T_103[287:0] : _GEN_2794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3845 = 10'ha7 == _T_13 ? _ram_T_103[287:0] : _GEN_2795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3846 = 10'ha8 == _T_13 ? _ram_T_103[287:0] : _GEN_2796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3847 = 10'ha9 == _T_13 ? _ram_T_103[287:0] : _GEN_2797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3848 = 10'haa == _T_13 ? _ram_T_103[287:0] : _GEN_2798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3849 = 10'hab == _T_13 ? _ram_T_103[287:0] : _GEN_2799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3850 = 10'hac == _T_13 ? _ram_T_103[287:0] : _GEN_2800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3851 = 10'had == _T_13 ? _ram_T_103[287:0] : _GEN_2801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3852 = 10'hae == _T_13 ? _ram_T_103[287:0] : _GEN_2802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3853 = 10'haf == _T_13 ? _ram_T_103[287:0] : _GEN_2803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3854 = 10'hb0 == _T_13 ? _ram_T_103[287:0] : _GEN_2804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3855 = 10'hb1 == _T_13 ? _ram_T_103[287:0] : _GEN_2805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3856 = 10'hb2 == _T_13 ? _ram_T_103[287:0] : _GEN_2806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3857 = 10'hb3 == _T_13 ? _ram_T_103[287:0] : _GEN_2807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3858 = 10'hb4 == _T_13 ? _ram_T_103[287:0] : _GEN_2808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3859 = 10'hb5 == _T_13 ? _ram_T_103[287:0] : _GEN_2809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3860 = 10'hb6 == _T_13 ? _ram_T_103[287:0] : _GEN_2810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3861 = 10'hb7 == _T_13 ? _ram_T_103[287:0] : _GEN_2811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3862 = 10'hb8 == _T_13 ? _ram_T_103[287:0] : _GEN_2812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3863 = 10'hb9 == _T_13 ? _ram_T_103[287:0] : _GEN_2813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3864 = 10'hba == _T_13 ? _ram_T_103[287:0] : _GEN_2814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3865 = 10'hbb == _T_13 ? _ram_T_103[287:0] : _GEN_2815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3866 = 10'hbc == _T_13 ? _ram_T_103[287:0] : _GEN_2816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3867 = 10'hbd == _T_13 ? _ram_T_103[287:0] : _GEN_2817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3868 = 10'hbe == _T_13 ? _ram_T_103[287:0] : _GEN_2818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3869 = 10'hbf == _T_13 ? _ram_T_103[287:0] : _GEN_2819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3870 = 10'hc0 == _T_13 ? _ram_T_103[287:0] : _GEN_2820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3871 = 10'hc1 == _T_13 ? _ram_T_103[287:0] : _GEN_2821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3872 = 10'hc2 == _T_13 ? _ram_T_103[287:0] : _GEN_2822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3873 = 10'hc3 == _T_13 ? _ram_T_103[287:0] : _GEN_2823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3874 = 10'hc4 == _T_13 ? _ram_T_103[287:0] : _GEN_2824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3875 = 10'hc5 == _T_13 ? _ram_T_103[287:0] : _GEN_2825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3876 = 10'hc6 == _T_13 ? _ram_T_103[287:0] : _GEN_2826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3877 = 10'hc7 == _T_13 ? _ram_T_103[287:0] : _GEN_2827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3878 = 10'hc8 == _T_13 ? _ram_T_103[287:0] : _GEN_2828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3879 = 10'hc9 == _T_13 ? _ram_T_103[287:0] : _GEN_2829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3880 = 10'hca == _T_13 ? _ram_T_103[287:0] : _GEN_2830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3881 = 10'hcb == _T_13 ? _ram_T_103[287:0] : _GEN_2831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3882 = 10'hcc == _T_13 ? _ram_T_103[287:0] : _GEN_2832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3883 = 10'hcd == _T_13 ? _ram_T_103[287:0] : _GEN_2833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3884 = 10'hce == _T_13 ? _ram_T_103[287:0] : _GEN_2834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3885 = 10'hcf == _T_13 ? _ram_T_103[287:0] : _GEN_2835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3886 = 10'hd0 == _T_13 ? _ram_T_103[287:0] : _GEN_2836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3887 = 10'hd1 == _T_13 ? _ram_T_103[287:0] : _GEN_2837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3888 = 10'hd2 == _T_13 ? _ram_T_103[287:0] : _GEN_2838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3889 = 10'hd3 == _T_13 ? _ram_T_103[287:0] : _GEN_2839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3890 = 10'hd4 == _T_13 ? _ram_T_103[287:0] : _GEN_2840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3891 = 10'hd5 == _T_13 ? _ram_T_103[287:0] : _GEN_2841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3892 = 10'hd6 == _T_13 ? _ram_T_103[287:0] : _GEN_2842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3893 = 10'hd7 == _T_13 ? _ram_T_103[287:0] : _GEN_2843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3894 = 10'hd8 == _T_13 ? _ram_T_103[287:0] : _GEN_2844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3895 = 10'hd9 == _T_13 ? _ram_T_103[287:0] : _GEN_2845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3896 = 10'hda == _T_13 ? _ram_T_103[287:0] : _GEN_2846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3897 = 10'hdb == _T_13 ? _ram_T_103[287:0] : _GEN_2847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3898 = 10'hdc == _T_13 ? _ram_T_103[287:0] : _GEN_2848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3899 = 10'hdd == _T_13 ? _ram_T_103[287:0] : _GEN_2849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3900 = 10'hde == _T_13 ? _ram_T_103[287:0] : _GEN_2850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3901 = 10'hdf == _T_13 ? _ram_T_103[287:0] : _GEN_2851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3902 = 10'he0 == _T_13 ? _ram_T_103[287:0] : _GEN_2852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3903 = 10'he1 == _T_13 ? _ram_T_103[287:0] : _GEN_2853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3904 = 10'he2 == _T_13 ? _ram_T_103[287:0] : _GEN_2854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3905 = 10'he3 == _T_13 ? _ram_T_103[287:0] : _GEN_2855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3906 = 10'he4 == _T_13 ? _ram_T_103[287:0] : _GEN_2856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3907 = 10'he5 == _T_13 ? _ram_T_103[287:0] : _GEN_2857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3908 = 10'he6 == _T_13 ? _ram_T_103[287:0] : _GEN_2858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3909 = 10'he7 == _T_13 ? _ram_T_103[287:0] : _GEN_2859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3910 = 10'he8 == _T_13 ? _ram_T_103[287:0] : _GEN_2860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3911 = 10'he9 == _T_13 ? _ram_T_103[287:0] : _GEN_2861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3912 = 10'hea == _T_13 ? _ram_T_103[287:0] : _GEN_2862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3913 = 10'heb == _T_13 ? _ram_T_103[287:0] : _GEN_2863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3914 = 10'hec == _T_13 ? _ram_T_103[287:0] : _GEN_2864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3915 = 10'hed == _T_13 ? _ram_T_103[287:0] : _GEN_2865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3916 = 10'hee == _T_13 ? _ram_T_103[287:0] : _GEN_2866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3917 = 10'hef == _T_13 ? _ram_T_103[287:0] : _GEN_2867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3918 = 10'hf0 == _T_13 ? _ram_T_103[287:0] : _GEN_2868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3919 = 10'hf1 == _T_13 ? _ram_T_103[287:0] : _GEN_2869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3920 = 10'hf2 == _T_13 ? _ram_T_103[287:0] : _GEN_2870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3921 = 10'hf3 == _T_13 ? _ram_T_103[287:0] : _GEN_2871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3922 = 10'hf4 == _T_13 ? _ram_T_103[287:0] : _GEN_2872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3923 = 10'hf5 == _T_13 ? _ram_T_103[287:0] : _GEN_2873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3924 = 10'hf6 == _T_13 ? _ram_T_103[287:0] : _GEN_2874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3925 = 10'hf7 == _T_13 ? _ram_T_103[287:0] : _GEN_2875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3926 = 10'hf8 == _T_13 ? _ram_T_103[287:0] : _GEN_2876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3927 = 10'hf9 == _T_13 ? _ram_T_103[287:0] : _GEN_2877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3928 = 10'hfa == _T_13 ? _ram_T_103[287:0] : _GEN_2878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3929 = 10'hfb == _T_13 ? _ram_T_103[287:0] : _GEN_2879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3930 = 10'hfc == _T_13 ? _ram_T_103[287:0] : _GEN_2880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3931 = 10'hfd == _T_13 ? _ram_T_103[287:0] : _GEN_2881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3932 = 10'hfe == _T_13 ? _ram_T_103[287:0] : _GEN_2882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3933 = 10'hff == _T_13 ? _ram_T_103[287:0] : _GEN_2883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3934 = 10'h100 == _T_13 ? _ram_T_103[287:0] : _GEN_2884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3935 = 10'h101 == _T_13 ? _ram_T_103[287:0] : _GEN_2885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3936 = 10'h102 == _T_13 ? _ram_T_103[287:0] : _GEN_2886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3937 = 10'h103 == _T_13 ? _ram_T_103[287:0] : _GEN_2887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3938 = 10'h104 == _T_13 ? _ram_T_103[287:0] : _GEN_2888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3939 = 10'h105 == _T_13 ? _ram_T_103[287:0] : _GEN_2889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3940 = 10'h106 == _T_13 ? _ram_T_103[287:0] : _GEN_2890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3941 = 10'h107 == _T_13 ? _ram_T_103[287:0] : _GEN_2891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3942 = 10'h108 == _T_13 ? _ram_T_103[287:0] : _GEN_2892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3943 = 10'h109 == _T_13 ? _ram_T_103[287:0] : _GEN_2893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3944 = 10'h10a == _T_13 ? _ram_T_103[287:0] : _GEN_2894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3945 = 10'h10b == _T_13 ? _ram_T_103[287:0] : _GEN_2895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3946 = 10'h10c == _T_13 ? _ram_T_103[287:0] : _GEN_2896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3947 = 10'h10d == _T_13 ? _ram_T_103[287:0] : _GEN_2897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3948 = 10'h10e == _T_13 ? _ram_T_103[287:0] : _GEN_2898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3949 = 10'h10f == _T_13 ? _ram_T_103[287:0] : _GEN_2899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3950 = 10'h110 == _T_13 ? _ram_T_103[287:0] : _GEN_2900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3951 = 10'h111 == _T_13 ? _ram_T_103[287:0] : _GEN_2901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3952 = 10'h112 == _T_13 ? _ram_T_103[287:0] : _GEN_2902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3953 = 10'h113 == _T_13 ? _ram_T_103[287:0] : _GEN_2903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3954 = 10'h114 == _T_13 ? _ram_T_103[287:0] : _GEN_2904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3955 = 10'h115 == _T_13 ? _ram_T_103[287:0] : _GEN_2905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3956 = 10'h116 == _T_13 ? _ram_T_103[287:0] : _GEN_2906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3957 = 10'h117 == _T_13 ? _ram_T_103[287:0] : _GEN_2907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3958 = 10'h118 == _T_13 ? _ram_T_103[287:0] : _GEN_2908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3959 = 10'h119 == _T_13 ? _ram_T_103[287:0] : _GEN_2909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3960 = 10'h11a == _T_13 ? _ram_T_103[287:0] : _GEN_2910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3961 = 10'h11b == _T_13 ? _ram_T_103[287:0] : _GEN_2911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3962 = 10'h11c == _T_13 ? _ram_T_103[287:0] : _GEN_2912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3963 = 10'h11d == _T_13 ? _ram_T_103[287:0] : _GEN_2913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3964 = 10'h11e == _T_13 ? _ram_T_103[287:0] : _GEN_2914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3965 = 10'h11f == _T_13 ? _ram_T_103[287:0] : _GEN_2915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3966 = 10'h120 == _T_13 ? _ram_T_103[287:0] : _GEN_2916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3967 = 10'h121 == _T_13 ? _ram_T_103[287:0] : _GEN_2917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3968 = 10'h122 == _T_13 ? _ram_T_103[287:0] : _GEN_2918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3969 = 10'h123 == _T_13 ? _ram_T_103[287:0] : _GEN_2919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3970 = 10'h124 == _T_13 ? _ram_T_103[287:0] : _GEN_2920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3971 = 10'h125 == _T_13 ? _ram_T_103[287:0] : _GEN_2921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3972 = 10'h126 == _T_13 ? _ram_T_103[287:0] : _GEN_2922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3973 = 10'h127 == _T_13 ? _ram_T_103[287:0] : _GEN_2923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3974 = 10'h128 == _T_13 ? _ram_T_103[287:0] : _GEN_2924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3975 = 10'h129 == _T_13 ? _ram_T_103[287:0] : _GEN_2925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3976 = 10'h12a == _T_13 ? _ram_T_103[287:0] : _GEN_2926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3977 = 10'h12b == _T_13 ? _ram_T_103[287:0] : _GEN_2927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3978 = 10'h12c == _T_13 ? _ram_T_103[287:0] : _GEN_2928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3979 = 10'h12d == _T_13 ? _ram_T_103[287:0] : _GEN_2929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3980 = 10'h12e == _T_13 ? _ram_T_103[287:0] : _GEN_2930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3981 = 10'h12f == _T_13 ? _ram_T_103[287:0] : _GEN_2931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3982 = 10'h130 == _T_13 ? _ram_T_103[287:0] : _GEN_2932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3983 = 10'h131 == _T_13 ? _ram_T_103[287:0] : _GEN_2933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3984 = 10'h132 == _T_13 ? _ram_T_103[287:0] : _GEN_2934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3985 = 10'h133 == _T_13 ? _ram_T_103[287:0] : _GEN_2935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3986 = 10'h134 == _T_13 ? _ram_T_103[287:0] : _GEN_2936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3987 = 10'h135 == _T_13 ? _ram_T_103[287:0] : _GEN_2937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3988 = 10'h136 == _T_13 ? _ram_T_103[287:0] : _GEN_2938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3989 = 10'h137 == _T_13 ? _ram_T_103[287:0] : _GEN_2939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3990 = 10'h138 == _T_13 ? _ram_T_103[287:0] : _GEN_2940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3991 = 10'h139 == _T_13 ? _ram_T_103[287:0] : _GEN_2941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3992 = 10'h13a == _T_13 ? _ram_T_103[287:0] : _GEN_2942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3993 = 10'h13b == _T_13 ? _ram_T_103[287:0] : _GEN_2943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3994 = 10'h13c == _T_13 ? _ram_T_103[287:0] : _GEN_2944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3995 = 10'h13d == _T_13 ? _ram_T_103[287:0] : _GEN_2945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3996 = 10'h13e == _T_13 ? _ram_T_103[287:0] : _GEN_2946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3997 = 10'h13f == _T_13 ? _ram_T_103[287:0] : _GEN_2947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3998 = 10'h140 == _T_13 ? _ram_T_103[287:0] : _GEN_2948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_3999 = 10'h141 == _T_13 ? _ram_T_103[287:0] : _GEN_2949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4000 = 10'h142 == _T_13 ? _ram_T_103[287:0] : _GEN_2950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4001 = 10'h143 == _T_13 ? _ram_T_103[287:0] : _GEN_2951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4002 = 10'h144 == _T_13 ? _ram_T_103[287:0] : _GEN_2952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4003 = 10'h145 == _T_13 ? _ram_T_103[287:0] : _GEN_2953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4004 = 10'h146 == _T_13 ? _ram_T_103[287:0] : _GEN_2954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4005 = 10'h147 == _T_13 ? _ram_T_103[287:0] : _GEN_2955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4006 = 10'h148 == _T_13 ? _ram_T_103[287:0] : _GEN_2956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4007 = 10'h149 == _T_13 ? _ram_T_103[287:0] : _GEN_2957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4008 = 10'h14a == _T_13 ? _ram_T_103[287:0] : _GEN_2958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4009 = 10'h14b == _T_13 ? _ram_T_103[287:0] : _GEN_2959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4010 = 10'h14c == _T_13 ? _ram_T_103[287:0] : _GEN_2960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4011 = 10'h14d == _T_13 ? _ram_T_103[287:0] : _GEN_2961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4012 = 10'h14e == _T_13 ? _ram_T_103[287:0] : _GEN_2962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4013 = 10'h14f == _T_13 ? _ram_T_103[287:0] : _GEN_2963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4014 = 10'h150 == _T_13 ? _ram_T_103[287:0] : _GEN_2964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4015 = 10'h151 == _T_13 ? _ram_T_103[287:0] : _GEN_2965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4016 = 10'h152 == _T_13 ? _ram_T_103[287:0] : _GEN_2966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4017 = 10'h153 == _T_13 ? _ram_T_103[287:0] : _GEN_2967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4018 = 10'h154 == _T_13 ? _ram_T_103[287:0] : _GEN_2968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4019 = 10'h155 == _T_13 ? _ram_T_103[287:0] : _GEN_2969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4020 = 10'h156 == _T_13 ? _ram_T_103[287:0] : _GEN_2970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4021 = 10'h157 == _T_13 ? _ram_T_103[287:0] : _GEN_2971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4022 = 10'h158 == _T_13 ? _ram_T_103[287:0] : _GEN_2972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4023 = 10'h159 == _T_13 ? _ram_T_103[287:0] : _GEN_2973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4024 = 10'h15a == _T_13 ? _ram_T_103[287:0] : _GEN_2974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4025 = 10'h15b == _T_13 ? _ram_T_103[287:0] : _GEN_2975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4026 = 10'h15c == _T_13 ? _ram_T_103[287:0] : _GEN_2976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4027 = 10'h15d == _T_13 ? _ram_T_103[287:0] : _GEN_2977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4028 = 10'h15e == _T_13 ? _ram_T_103[287:0] : _GEN_2978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4029 = 10'h15f == _T_13 ? _ram_T_103[287:0] : _GEN_2979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4030 = 10'h160 == _T_13 ? _ram_T_103[287:0] : _GEN_2980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4031 = 10'h161 == _T_13 ? _ram_T_103[287:0] : _GEN_2981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4032 = 10'h162 == _T_13 ? _ram_T_103[287:0] : _GEN_2982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4033 = 10'h163 == _T_13 ? _ram_T_103[287:0] : _GEN_2983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4034 = 10'h164 == _T_13 ? _ram_T_103[287:0] : _GEN_2984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4035 = 10'h165 == _T_13 ? _ram_T_103[287:0] : _GEN_2985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4036 = 10'h166 == _T_13 ? _ram_T_103[287:0] : _GEN_2986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4037 = 10'h167 == _T_13 ? _ram_T_103[287:0] : _GEN_2987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4038 = 10'h168 == _T_13 ? _ram_T_103[287:0] : _GEN_2988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4039 = 10'h169 == _T_13 ? _ram_T_103[287:0] : _GEN_2989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4040 = 10'h16a == _T_13 ? _ram_T_103[287:0] : _GEN_2990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4041 = 10'h16b == _T_13 ? _ram_T_103[287:0] : _GEN_2991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4042 = 10'h16c == _T_13 ? _ram_T_103[287:0] : _GEN_2992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4043 = 10'h16d == _T_13 ? _ram_T_103[287:0] : _GEN_2993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4044 = 10'h16e == _T_13 ? _ram_T_103[287:0] : _GEN_2994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4045 = 10'h16f == _T_13 ? _ram_T_103[287:0] : _GEN_2995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4046 = 10'h170 == _T_13 ? _ram_T_103[287:0] : _GEN_2996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4047 = 10'h171 == _T_13 ? _ram_T_103[287:0] : _GEN_2997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4048 = 10'h172 == _T_13 ? _ram_T_103[287:0] : _GEN_2998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4049 = 10'h173 == _T_13 ? _ram_T_103[287:0] : _GEN_2999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4050 = 10'h174 == _T_13 ? _ram_T_103[287:0] : _GEN_3000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4051 = 10'h175 == _T_13 ? _ram_T_103[287:0] : _GEN_3001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4052 = 10'h176 == _T_13 ? _ram_T_103[287:0] : _GEN_3002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4053 = 10'h177 == _T_13 ? _ram_T_103[287:0] : _GEN_3003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4054 = 10'h178 == _T_13 ? _ram_T_103[287:0] : _GEN_3004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4055 = 10'h179 == _T_13 ? _ram_T_103[287:0] : _GEN_3005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4056 = 10'h17a == _T_13 ? _ram_T_103[287:0] : _GEN_3006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4057 = 10'h17b == _T_13 ? _ram_T_103[287:0] : _GEN_3007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4058 = 10'h17c == _T_13 ? _ram_T_103[287:0] : _GEN_3008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4059 = 10'h17d == _T_13 ? _ram_T_103[287:0] : _GEN_3009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4060 = 10'h17e == _T_13 ? _ram_T_103[287:0] : _GEN_3010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4061 = 10'h17f == _T_13 ? _ram_T_103[287:0] : _GEN_3011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4062 = 10'h180 == _T_13 ? _ram_T_103[287:0] : _GEN_3012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4063 = 10'h181 == _T_13 ? _ram_T_103[287:0] : _GEN_3013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4064 = 10'h182 == _T_13 ? _ram_T_103[287:0] : _GEN_3014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4065 = 10'h183 == _T_13 ? _ram_T_103[287:0] : _GEN_3015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4066 = 10'h184 == _T_13 ? _ram_T_103[287:0] : _GEN_3016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4067 = 10'h185 == _T_13 ? _ram_T_103[287:0] : _GEN_3017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4068 = 10'h186 == _T_13 ? _ram_T_103[287:0] : _GEN_3018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4069 = 10'h187 == _T_13 ? _ram_T_103[287:0] : _GEN_3019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4070 = 10'h188 == _T_13 ? _ram_T_103[287:0] : _GEN_3020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4071 = 10'h189 == _T_13 ? _ram_T_103[287:0] : _GEN_3021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4072 = 10'h18a == _T_13 ? _ram_T_103[287:0] : _GEN_3022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4073 = 10'h18b == _T_13 ? _ram_T_103[287:0] : _GEN_3023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4074 = 10'h18c == _T_13 ? _ram_T_103[287:0] : _GEN_3024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4075 = 10'h18d == _T_13 ? _ram_T_103[287:0] : _GEN_3025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4076 = 10'h18e == _T_13 ? _ram_T_103[287:0] : _GEN_3026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4077 = 10'h18f == _T_13 ? _ram_T_103[287:0] : _GEN_3027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4078 = 10'h190 == _T_13 ? _ram_T_103[287:0] : _GEN_3028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4079 = 10'h191 == _T_13 ? _ram_T_103[287:0] : _GEN_3029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4080 = 10'h192 == _T_13 ? _ram_T_103[287:0] : _GEN_3030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4081 = 10'h193 == _T_13 ? _ram_T_103[287:0] : _GEN_3031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4082 = 10'h194 == _T_13 ? _ram_T_103[287:0] : _GEN_3032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4083 = 10'h195 == _T_13 ? _ram_T_103[287:0] : _GEN_3033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4084 = 10'h196 == _T_13 ? _ram_T_103[287:0] : _GEN_3034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4085 = 10'h197 == _T_13 ? _ram_T_103[287:0] : _GEN_3035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4086 = 10'h198 == _T_13 ? _ram_T_103[287:0] : _GEN_3036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4087 = 10'h199 == _T_13 ? _ram_T_103[287:0] : _GEN_3037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4088 = 10'h19a == _T_13 ? _ram_T_103[287:0] : _GEN_3038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4089 = 10'h19b == _T_13 ? _ram_T_103[287:0] : _GEN_3039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4090 = 10'h19c == _T_13 ? _ram_T_103[287:0] : _GEN_3040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4091 = 10'h19d == _T_13 ? _ram_T_103[287:0] : _GEN_3041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4092 = 10'h19e == _T_13 ? _ram_T_103[287:0] : _GEN_3042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4093 = 10'h19f == _T_13 ? _ram_T_103[287:0] : _GEN_3043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4094 = 10'h1a0 == _T_13 ? _ram_T_103[287:0] : _GEN_3044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4095 = 10'h1a1 == _T_13 ? _ram_T_103[287:0] : _GEN_3045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4096 = 10'h1a2 == _T_13 ? _ram_T_103[287:0] : _GEN_3046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4097 = 10'h1a3 == _T_13 ? _ram_T_103[287:0] : _GEN_3047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4098 = 10'h1a4 == _T_13 ? _ram_T_103[287:0] : _GEN_3048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4099 = 10'h1a5 == _T_13 ? _ram_T_103[287:0] : _GEN_3049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4100 = 10'h1a6 == _T_13 ? _ram_T_103[287:0] : _GEN_3050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4101 = 10'h1a7 == _T_13 ? _ram_T_103[287:0] : _GEN_3051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4102 = 10'h1a8 == _T_13 ? _ram_T_103[287:0] : _GEN_3052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4103 = 10'h1a9 == _T_13 ? _ram_T_103[287:0] : _GEN_3053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4104 = 10'h1aa == _T_13 ? _ram_T_103[287:0] : _GEN_3054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4105 = 10'h1ab == _T_13 ? _ram_T_103[287:0] : _GEN_3055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4106 = 10'h1ac == _T_13 ? _ram_T_103[287:0] : _GEN_3056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4107 = 10'h1ad == _T_13 ? _ram_T_103[287:0] : _GEN_3057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4108 = 10'h1ae == _T_13 ? _ram_T_103[287:0] : _GEN_3058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4109 = 10'h1af == _T_13 ? _ram_T_103[287:0] : _GEN_3059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4110 = 10'h1b0 == _T_13 ? _ram_T_103[287:0] : _GEN_3060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4111 = 10'h1b1 == _T_13 ? _ram_T_103[287:0] : _GEN_3061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4112 = 10'h1b2 == _T_13 ? _ram_T_103[287:0] : _GEN_3062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4113 = 10'h1b3 == _T_13 ? _ram_T_103[287:0] : _GEN_3063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4114 = 10'h1b4 == _T_13 ? _ram_T_103[287:0] : _GEN_3064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4115 = 10'h1b5 == _T_13 ? _ram_T_103[287:0] : _GEN_3065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4116 = 10'h1b6 == _T_13 ? _ram_T_103[287:0] : _GEN_3066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4117 = 10'h1b7 == _T_13 ? _ram_T_103[287:0] : _GEN_3067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4118 = 10'h1b8 == _T_13 ? _ram_T_103[287:0] : _GEN_3068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4119 = 10'h1b9 == _T_13 ? _ram_T_103[287:0] : _GEN_3069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4120 = 10'h1ba == _T_13 ? _ram_T_103[287:0] : _GEN_3070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4121 = 10'h1bb == _T_13 ? _ram_T_103[287:0] : _GEN_3071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4122 = 10'h1bc == _T_13 ? _ram_T_103[287:0] : _GEN_3072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4123 = 10'h1bd == _T_13 ? _ram_T_103[287:0] : _GEN_3073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4124 = 10'h1be == _T_13 ? _ram_T_103[287:0] : _GEN_3074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4125 = 10'h1bf == _T_13 ? _ram_T_103[287:0] : _GEN_3075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4126 = 10'h1c0 == _T_13 ? _ram_T_103[287:0] : _GEN_3076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4127 = 10'h1c1 == _T_13 ? _ram_T_103[287:0] : _GEN_3077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4128 = 10'h1c2 == _T_13 ? _ram_T_103[287:0] : _GEN_3078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4129 = 10'h1c3 == _T_13 ? _ram_T_103[287:0] : _GEN_3079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4130 = 10'h1c4 == _T_13 ? _ram_T_103[287:0] : _GEN_3080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4131 = 10'h1c5 == _T_13 ? _ram_T_103[287:0] : _GEN_3081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4132 = 10'h1c6 == _T_13 ? _ram_T_103[287:0] : _GEN_3082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4133 = 10'h1c7 == _T_13 ? _ram_T_103[287:0] : _GEN_3083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4134 = 10'h1c8 == _T_13 ? _ram_T_103[287:0] : _GEN_3084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4135 = 10'h1c9 == _T_13 ? _ram_T_103[287:0] : _GEN_3085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4136 = 10'h1ca == _T_13 ? _ram_T_103[287:0] : _GEN_3086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4137 = 10'h1cb == _T_13 ? _ram_T_103[287:0] : _GEN_3087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4138 = 10'h1cc == _T_13 ? _ram_T_103[287:0] : _GEN_3088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4139 = 10'h1cd == _T_13 ? _ram_T_103[287:0] : _GEN_3089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4140 = 10'h1ce == _T_13 ? _ram_T_103[287:0] : _GEN_3090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4141 = 10'h1cf == _T_13 ? _ram_T_103[287:0] : _GEN_3091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4142 = 10'h1d0 == _T_13 ? _ram_T_103[287:0] : _GEN_3092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4143 = 10'h1d1 == _T_13 ? _ram_T_103[287:0] : _GEN_3093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4144 = 10'h1d2 == _T_13 ? _ram_T_103[287:0] : _GEN_3094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4145 = 10'h1d3 == _T_13 ? _ram_T_103[287:0] : _GEN_3095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4146 = 10'h1d4 == _T_13 ? _ram_T_103[287:0] : _GEN_3096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4147 = 10'h1d5 == _T_13 ? _ram_T_103[287:0] : _GEN_3097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4148 = 10'h1d6 == _T_13 ? _ram_T_103[287:0] : _GEN_3098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4149 = 10'h1d7 == _T_13 ? _ram_T_103[287:0] : _GEN_3099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4150 = 10'h1d8 == _T_13 ? _ram_T_103[287:0] : _GEN_3100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4151 = 10'h1d9 == _T_13 ? _ram_T_103[287:0] : _GEN_3101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4152 = 10'h1da == _T_13 ? _ram_T_103[287:0] : _GEN_3102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4153 = 10'h1db == _T_13 ? _ram_T_103[287:0] : _GEN_3103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4154 = 10'h1dc == _T_13 ? _ram_T_103[287:0] : _GEN_3104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4155 = 10'h1dd == _T_13 ? _ram_T_103[287:0] : _GEN_3105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4156 = 10'h1de == _T_13 ? _ram_T_103[287:0] : _GEN_3106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4157 = 10'h1df == _T_13 ? _ram_T_103[287:0] : _GEN_3107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4158 = 10'h1e0 == _T_13 ? _ram_T_103[287:0] : _GEN_3108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4159 = 10'h1e1 == _T_13 ? _ram_T_103[287:0] : _GEN_3109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4160 = 10'h1e2 == _T_13 ? _ram_T_103[287:0] : _GEN_3110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4161 = 10'h1e3 == _T_13 ? _ram_T_103[287:0] : _GEN_3111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4162 = 10'h1e4 == _T_13 ? _ram_T_103[287:0] : _GEN_3112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4163 = 10'h1e5 == _T_13 ? _ram_T_103[287:0] : _GEN_3113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4164 = 10'h1e6 == _T_13 ? _ram_T_103[287:0] : _GEN_3114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4165 = 10'h1e7 == _T_13 ? _ram_T_103[287:0] : _GEN_3115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4166 = 10'h1e8 == _T_13 ? _ram_T_103[287:0] : _GEN_3116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4167 = 10'h1e9 == _T_13 ? _ram_T_103[287:0] : _GEN_3117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4168 = 10'h1ea == _T_13 ? _ram_T_103[287:0] : _GEN_3118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4169 = 10'h1eb == _T_13 ? _ram_T_103[287:0] : _GEN_3119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4170 = 10'h1ec == _T_13 ? _ram_T_103[287:0] : _GEN_3120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4171 = 10'h1ed == _T_13 ? _ram_T_103[287:0] : _GEN_3121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4172 = 10'h1ee == _T_13 ? _ram_T_103[287:0] : _GEN_3122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4173 = 10'h1ef == _T_13 ? _ram_T_103[287:0] : _GEN_3123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4174 = 10'h1f0 == _T_13 ? _ram_T_103[287:0] : _GEN_3124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4175 = 10'h1f1 == _T_13 ? _ram_T_103[287:0] : _GEN_3125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4176 = 10'h1f2 == _T_13 ? _ram_T_103[287:0] : _GEN_3126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4177 = 10'h1f3 == _T_13 ? _ram_T_103[287:0] : _GEN_3127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4178 = 10'h1f4 == _T_13 ? _ram_T_103[287:0] : _GEN_3128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4179 = 10'h1f5 == _T_13 ? _ram_T_103[287:0] : _GEN_3129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4180 = 10'h1f6 == _T_13 ? _ram_T_103[287:0] : _GEN_3130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4181 = 10'h1f7 == _T_13 ? _ram_T_103[287:0] : _GEN_3131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4182 = 10'h1f8 == _T_13 ? _ram_T_103[287:0] : _GEN_3132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4183 = 10'h1f9 == _T_13 ? _ram_T_103[287:0] : _GEN_3133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4184 = 10'h1fa == _T_13 ? _ram_T_103[287:0] : _GEN_3134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4185 = 10'h1fb == _T_13 ? _ram_T_103[287:0] : _GEN_3135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4186 = 10'h1fc == _T_13 ? _ram_T_103[287:0] : _GEN_3136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4187 = 10'h1fd == _T_13 ? _ram_T_103[287:0] : _GEN_3137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4188 = 10'h1fe == _T_13 ? _ram_T_103[287:0] : _GEN_3138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4189 = 10'h1ff == _T_13 ? _ram_T_103[287:0] : _GEN_3139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4190 = 10'h200 == _T_13 ? _ram_T_103[287:0] : _GEN_3140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4191 = 10'h201 == _T_13 ? _ram_T_103[287:0] : _GEN_3141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4192 = 10'h202 == _T_13 ? _ram_T_103[287:0] : _GEN_3142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4193 = 10'h203 == _T_13 ? _ram_T_103[287:0] : _GEN_3143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4194 = 10'h204 == _T_13 ? _ram_T_103[287:0] : _GEN_3144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4195 = 10'h205 == _T_13 ? _ram_T_103[287:0] : _GEN_3145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4196 = 10'h206 == _T_13 ? _ram_T_103[287:0] : _GEN_3146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4197 = 10'h207 == _T_13 ? _ram_T_103[287:0] : _GEN_3147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4198 = 10'h208 == _T_13 ? _ram_T_103[287:0] : _GEN_3148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4199 = 10'h209 == _T_13 ? _ram_T_103[287:0] : _GEN_3149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4200 = 10'h20a == _T_13 ? _ram_T_103[287:0] : _GEN_3150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4201 = 10'h20b == _T_13 ? _ram_T_103[287:0] : _GEN_3151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4202 = 10'h20c == _T_13 ? _ram_T_103[287:0] : _GEN_3152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_15 = h + 10'h4; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_4 = vga_mem_ram_MPORT_36_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_4 = vga_mem_ram_MPORT_37_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_4 = vga_mem_ram_MPORT_38_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_4 = vga_mem_ram_MPORT_39_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_4 = vga_mem_ram_MPORT_40_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_4 = vga_mem_ram_MPORT_41_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_4 = vga_mem_ram_MPORT_42_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_4 = vga_mem_ram_MPORT_43_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_4 = vga_mem_ram_MPORT_44_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_124 = {278'h0,ram_hi_hi_hi_lo_4,ram_hi_hi_lo_4,ram_hi_lo_hi_4,ram_hi_lo_lo_4,ram_lo_hi_hi_hi_4,
    ram_lo_hi_hi_lo_4,ram_lo_hi_lo_4,ram_lo_lo_hi_4,ram_lo_lo_lo_4}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19068 = {{8191'd0}, _ram_T_124}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_128 = _GEN_19068 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_4204 = 10'h1 == _T_15 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4205 = 10'h2 == _T_15 ? ram_2 : _GEN_4204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4206 = 10'h3 == _T_15 ? ram_3 : _GEN_4205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4207 = 10'h4 == _T_15 ? ram_4 : _GEN_4206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4208 = 10'h5 == _T_15 ? ram_5 : _GEN_4207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4209 = 10'h6 == _T_15 ? ram_6 : _GEN_4208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4210 = 10'h7 == _T_15 ? ram_7 : _GEN_4209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4211 = 10'h8 == _T_15 ? ram_8 : _GEN_4210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4212 = 10'h9 == _T_15 ? ram_9 : _GEN_4211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4213 = 10'ha == _T_15 ? ram_10 : _GEN_4212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4214 = 10'hb == _T_15 ? ram_11 : _GEN_4213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4215 = 10'hc == _T_15 ? ram_12 : _GEN_4214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4216 = 10'hd == _T_15 ? ram_13 : _GEN_4215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4217 = 10'he == _T_15 ? ram_14 : _GEN_4216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4218 = 10'hf == _T_15 ? ram_15 : _GEN_4217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4219 = 10'h10 == _T_15 ? ram_16 : _GEN_4218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4220 = 10'h11 == _T_15 ? ram_17 : _GEN_4219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4221 = 10'h12 == _T_15 ? ram_18 : _GEN_4220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4222 = 10'h13 == _T_15 ? ram_19 : _GEN_4221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4223 = 10'h14 == _T_15 ? ram_20 : _GEN_4222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4224 = 10'h15 == _T_15 ? ram_21 : _GEN_4223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4225 = 10'h16 == _T_15 ? ram_22 : _GEN_4224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4226 = 10'h17 == _T_15 ? ram_23 : _GEN_4225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4227 = 10'h18 == _T_15 ? ram_24 : _GEN_4226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4228 = 10'h19 == _T_15 ? ram_25 : _GEN_4227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4229 = 10'h1a == _T_15 ? ram_26 : _GEN_4228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4230 = 10'h1b == _T_15 ? ram_27 : _GEN_4229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4231 = 10'h1c == _T_15 ? ram_28 : _GEN_4230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4232 = 10'h1d == _T_15 ? ram_29 : _GEN_4231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4233 = 10'h1e == _T_15 ? ram_30 : _GEN_4232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4234 = 10'h1f == _T_15 ? ram_31 : _GEN_4233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4235 = 10'h20 == _T_15 ? ram_32 : _GEN_4234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4236 = 10'h21 == _T_15 ? ram_33 : _GEN_4235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4237 = 10'h22 == _T_15 ? ram_34 : _GEN_4236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4238 = 10'h23 == _T_15 ? ram_35 : _GEN_4237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4239 = 10'h24 == _T_15 ? ram_36 : _GEN_4238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4240 = 10'h25 == _T_15 ? ram_37 : _GEN_4239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4241 = 10'h26 == _T_15 ? ram_38 : _GEN_4240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4242 = 10'h27 == _T_15 ? ram_39 : _GEN_4241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4243 = 10'h28 == _T_15 ? ram_40 : _GEN_4242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4244 = 10'h29 == _T_15 ? ram_41 : _GEN_4243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4245 = 10'h2a == _T_15 ? ram_42 : _GEN_4244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4246 = 10'h2b == _T_15 ? ram_43 : _GEN_4245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4247 = 10'h2c == _T_15 ? ram_44 : _GEN_4246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4248 = 10'h2d == _T_15 ? ram_45 : _GEN_4247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4249 = 10'h2e == _T_15 ? ram_46 : _GEN_4248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4250 = 10'h2f == _T_15 ? ram_47 : _GEN_4249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4251 = 10'h30 == _T_15 ? ram_48 : _GEN_4250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4252 = 10'h31 == _T_15 ? ram_49 : _GEN_4251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4253 = 10'h32 == _T_15 ? ram_50 : _GEN_4252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4254 = 10'h33 == _T_15 ? ram_51 : _GEN_4253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4255 = 10'h34 == _T_15 ? ram_52 : _GEN_4254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4256 = 10'h35 == _T_15 ? ram_53 : _GEN_4255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4257 = 10'h36 == _T_15 ? ram_54 : _GEN_4256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4258 = 10'h37 == _T_15 ? ram_55 : _GEN_4257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4259 = 10'h38 == _T_15 ? ram_56 : _GEN_4258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4260 = 10'h39 == _T_15 ? ram_57 : _GEN_4259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4261 = 10'h3a == _T_15 ? ram_58 : _GEN_4260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4262 = 10'h3b == _T_15 ? ram_59 : _GEN_4261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4263 = 10'h3c == _T_15 ? ram_60 : _GEN_4262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4264 = 10'h3d == _T_15 ? ram_61 : _GEN_4263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4265 = 10'h3e == _T_15 ? ram_62 : _GEN_4264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4266 = 10'h3f == _T_15 ? ram_63 : _GEN_4265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4267 = 10'h40 == _T_15 ? ram_64 : _GEN_4266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4268 = 10'h41 == _T_15 ? ram_65 : _GEN_4267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4269 = 10'h42 == _T_15 ? ram_66 : _GEN_4268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4270 = 10'h43 == _T_15 ? ram_67 : _GEN_4269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4271 = 10'h44 == _T_15 ? ram_68 : _GEN_4270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4272 = 10'h45 == _T_15 ? ram_69 : _GEN_4271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4273 = 10'h46 == _T_15 ? ram_70 : _GEN_4272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4274 = 10'h47 == _T_15 ? ram_71 : _GEN_4273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4275 = 10'h48 == _T_15 ? ram_72 : _GEN_4274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4276 = 10'h49 == _T_15 ? ram_73 : _GEN_4275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4277 = 10'h4a == _T_15 ? ram_74 : _GEN_4276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4278 = 10'h4b == _T_15 ? ram_75 : _GEN_4277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4279 = 10'h4c == _T_15 ? ram_76 : _GEN_4278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4280 = 10'h4d == _T_15 ? ram_77 : _GEN_4279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4281 = 10'h4e == _T_15 ? ram_78 : _GEN_4280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4282 = 10'h4f == _T_15 ? ram_79 : _GEN_4281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4283 = 10'h50 == _T_15 ? ram_80 : _GEN_4282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4284 = 10'h51 == _T_15 ? ram_81 : _GEN_4283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4285 = 10'h52 == _T_15 ? ram_82 : _GEN_4284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4286 = 10'h53 == _T_15 ? ram_83 : _GEN_4285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4287 = 10'h54 == _T_15 ? ram_84 : _GEN_4286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4288 = 10'h55 == _T_15 ? ram_85 : _GEN_4287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4289 = 10'h56 == _T_15 ? ram_86 : _GEN_4288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4290 = 10'h57 == _T_15 ? ram_87 : _GEN_4289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4291 = 10'h58 == _T_15 ? ram_88 : _GEN_4290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4292 = 10'h59 == _T_15 ? ram_89 : _GEN_4291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4293 = 10'h5a == _T_15 ? ram_90 : _GEN_4292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4294 = 10'h5b == _T_15 ? ram_91 : _GEN_4293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4295 = 10'h5c == _T_15 ? ram_92 : _GEN_4294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4296 = 10'h5d == _T_15 ? ram_93 : _GEN_4295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4297 = 10'h5e == _T_15 ? ram_94 : _GEN_4296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4298 = 10'h5f == _T_15 ? ram_95 : _GEN_4297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4299 = 10'h60 == _T_15 ? ram_96 : _GEN_4298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4300 = 10'h61 == _T_15 ? ram_97 : _GEN_4299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4301 = 10'h62 == _T_15 ? ram_98 : _GEN_4300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4302 = 10'h63 == _T_15 ? ram_99 : _GEN_4301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4303 = 10'h64 == _T_15 ? ram_100 : _GEN_4302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4304 = 10'h65 == _T_15 ? ram_101 : _GEN_4303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4305 = 10'h66 == _T_15 ? ram_102 : _GEN_4304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4306 = 10'h67 == _T_15 ? ram_103 : _GEN_4305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4307 = 10'h68 == _T_15 ? ram_104 : _GEN_4306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4308 = 10'h69 == _T_15 ? ram_105 : _GEN_4307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4309 = 10'h6a == _T_15 ? ram_106 : _GEN_4308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4310 = 10'h6b == _T_15 ? ram_107 : _GEN_4309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4311 = 10'h6c == _T_15 ? ram_108 : _GEN_4310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4312 = 10'h6d == _T_15 ? ram_109 : _GEN_4311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4313 = 10'h6e == _T_15 ? ram_110 : _GEN_4312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4314 = 10'h6f == _T_15 ? ram_111 : _GEN_4313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4315 = 10'h70 == _T_15 ? ram_112 : _GEN_4314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4316 = 10'h71 == _T_15 ? ram_113 : _GEN_4315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4317 = 10'h72 == _T_15 ? ram_114 : _GEN_4316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4318 = 10'h73 == _T_15 ? ram_115 : _GEN_4317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4319 = 10'h74 == _T_15 ? ram_116 : _GEN_4318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4320 = 10'h75 == _T_15 ? ram_117 : _GEN_4319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4321 = 10'h76 == _T_15 ? ram_118 : _GEN_4320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4322 = 10'h77 == _T_15 ? ram_119 : _GEN_4321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4323 = 10'h78 == _T_15 ? ram_120 : _GEN_4322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4324 = 10'h79 == _T_15 ? ram_121 : _GEN_4323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4325 = 10'h7a == _T_15 ? ram_122 : _GEN_4324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4326 = 10'h7b == _T_15 ? ram_123 : _GEN_4325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4327 = 10'h7c == _T_15 ? ram_124 : _GEN_4326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4328 = 10'h7d == _T_15 ? ram_125 : _GEN_4327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4329 = 10'h7e == _T_15 ? ram_126 : _GEN_4328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4330 = 10'h7f == _T_15 ? ram_127 : _GEN_4329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4331 = 10'h80 == _T_15 ? ram_128 : _GEN_4330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4332 = 10'h81 == _T_15 ? ram_129 : _GEN_4331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4333 = 10'h82 == _T_15 ? ram_130 : _GEN_4332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4334 = 10'h83 == _T_15 ? ram_131 : _GEN_4333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4335 = 10'h84 == _T_15 ? ram_132 : _GEN_4334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4336 = 10'h85 == _T_15 ? ram_133 : _GEN_4335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4337 = 10'h86 == _T_15 ? ram_134 : _GEN_4336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4338 = 10'h87 == _T_15 ? ram_135 : _GEN_4337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4339 = 10'h88 == _T_15 ? ram_136 : _GEN_4338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4340 = 10'h89 == _T_15 ? ram_137 : _GEN_4339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4341 = 10'h8a == _T_15 ? ram_138 : _GEN_4340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4342 = 10'h8b == _T_15 ? ram_139 : _GEN_4341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4343 = 10'h8c == _T_15 ? ram_140 : _GEN_4342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4344 = 10'h8d == _T_15 ? ram_141 : _GEN_4343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4345 = 10'h8e == _T_15 ? ram_142 : _GEN_4344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4346 = 10'h8f == _T_15 ? ram_143 : _GEN_4345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4347 = 10'h90 == _T_15 ? ram_144 : _GEN_4346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4348 = 10'h91 == _T_15 ? ram_145 : _GEN_4347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4349 = 10'h92 == _T_15 ? ram_146 : _GEN_4348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4350 = 10'h93 == _T_15 ? ram_147 : _GEN_4349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4351 = 10'h94 == _T_15 ? ram_148 : _GEN_4350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4352 = 10'h95 == _T_15 ? ram_149 : _GEN_4351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4353 = 10'h96 == _T_15 ? ram_150 : _GEN_4352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4354 = 10'h97 == _T_15 ? ram_151 : _GEN_4353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4355 = 10'h98 == _T_15 ? ram_152 : _GEN_4354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4356 = 10'h99 == _T_15 ? ram_153 : _GEN_4355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4357 = 10'h9a == _T_15 ? ram_154 : _GEN_4356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4358 = 10'h9b == _T_15 ? ram_155 : _GEN_4357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4359 = 10'h9c == _T_15 ? ram_156 : _GEN_4358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4360 = 10'h9d == _T_15 ? ram_157 : _GEN_4359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4361 = 10'h9e == _T_15 ? ram_158 : _GEN_4360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4362 = 10'h9f == _T_15 ? ram_159 : _GEN_4361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4363 = 10'ha0 == _T_15 ? ram_160 : _GEN_4362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4364 = 10'ha1 == _T_15 ? ram_161 : _GEN_4363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4365 = 10'ha2 == _T_15 ? ram_162 : _GEN_4364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4366 = 10'ha3 == _T_15 ? ram_163 : _GEN_4365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4367 = 10'ha4 == _T_15 ? ram_164 : _GEN_4366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4368 = 10'ha5 == _T_15 ? ram_165 : _GEN_4367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4369 = 10'ha6 == _T_15 ? ram_166 : _GEN_4368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4370 = 10'ha7 == _T_15 ? ram_167 : _GEN_4369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4371 = 10'ha8 == _T_15 ? ram_168 : _GEN_4370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4372 = 10'ha9 == _T_15 ? ram_169 : _GEN_4371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4373 = 10'haa == _T_15 ? ram_170 : _GEN_4372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4374 = 10'hab == _T_15 ? ram_171 : _GEN_4373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4375 = 10'hac == _T_15 ? ram_172 : _GEN_4374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4376 = 10'had == _T_15 ? ram_173 : _GEN_4375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4377 = 10'hae == _T_15 ? ram_174 : _GEN_4376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4378 = 10'haf == _T_15 ? ram_175 : _GEN_4377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4379 = 10'hb0 == _T_15 ? ram_176 : _GEN_4378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4380 = 10'hb1 == _T_15 ? ram_177 : _GEN_4379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4381 = 10'hb2 == _T_15 ? ram_178 : _GEN_4380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4382 = 10'hb3 == _T_15 ? ram_179 : _GEN_4381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4383 = 10'hb4 == _T_15 ? ram_180 : _GEN_4382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4384 = 10'hb5 == _T_15 ? ram_181 : _GEN_4383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4385 = 10'hb6 == _T_15 ? ram_182 : _GEN_4384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4386 = 10'hb7 == _T_15 ? ram_183 : _GEN_4385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4387 = 10'hb8 == _T_15 ? ram_184 : _GEN_4386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4388 = 10'hb9 == _T_15 ? ram_185 : _GEN_4387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4389 = 10'hba == _T_15 ? ram_186 : _GEN_4388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4390 = 10'hbb == _T_15 ? ram_187 : _GEN_4389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4391 = 10'hbc == _T_15 ? ram_188 : _GEN_4390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4392 = 10'hbd == _T_15 ? ram_189 : _GEN_4391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4393 = 10'hbe == _T_15 ? ram_190 : _GEN_4392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4394 = 10'hbf == _T_15 ? ram_191 : _GEN_4393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4395 = 10'hc0 == _T_15 ? ram_192 : _GEN_4394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4396 = 10'hc1 == _T_15 ? ram_193 : _GEN_4395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4397 = 10'hc2 == _T_15 ? ram_194 : _GEN_4396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4398 = 10'hc3 == _T_15 ? ram_195 : _GEN_4397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4399 = 10'hc4 == _T_15 ? ram_196 : _GEN_4398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4400 = 10'hc5 == _T_15 ? ram_197 : _GEN_4399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4401 = 10'hc6 == _T_15 ? ram_198 : _GEN_4400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4402 = 10'hc7 == _T_15 ? ram_199 : _GEN_4401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4403 = 10'hc8 == _T_15 ? ram_200 : _GEN_4402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4404 = 10'hc9 == _T_15 ? ram_201 : _GEN_4403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4405 = 10'hca == _T_15 ? ram_202 : _GEN_4404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4406 = 10'hcb == _T_15 ? ram_203 : _GEN_4405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4407 = 10'hcc == _T_15 ? ram_204 : _GEN_4406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4408 = 10'hcd == _T_15 ? ram_205 : _GEN_4407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4409 = 10'hce == _T_15 ? ram_206 : _GEN_4408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4410 = 10'hcf == _T_15 ? ram_207 : _GEN_4409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4411 = 10'hd0 == _T_15 ? ram_208 : _GEN_4410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4412 = 10'hd1 == _T_15 ? ram_209 : _GEN_4411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4413 = 10'hd2 == _T_15 ? ram_210 : _GEN_4412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4414 = 10'hd3 == _T_15 ? ram_211 : _GEN_4413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4415 = 10'hd4 == _T_15 ? ram_212 : _GEN_4414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4416 = 10'hd5 == _T_15 ? ram_213 : _GEN_4415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4417 = 10'hd6 == _T_15 ? ram_214 : _GEN_4416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4418 = 10'hd7 == _T_15 ? ram_215 : _GEN_4417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4419 = 10'hd8 == _T_15 ? ram_216 : _GEN_4418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4420 = 10'hd9 == _T_15 ? ram_217 : _GEN_4419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4421 = 10'hda == _T_15 ? ram_218 : _GEN_4420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4422 = 10'hdb == _T_15 ? ram_219 : _GEN_4421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4423 = 10'hdc == _T_15 ? ram_220 : _GEN_4422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4424 = 10'hdd == _T_15 ? ram_221 : _GEN_4423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4425 = 10'hde == _T_15 ? ram_222 : _GEN_4424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4426 = 10'hdf == _T_15 ? ram_223 : _GEN_4425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4427 = 10'he0 == _T_15 ? ram_224 : _GEN_4426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4428 = 10'he1 == _T_15 ? ram_225 : _GEN_4427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4429 = 10'he2 == _T_15 ? ram_226 : _GEN_4428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4430 = 10'he3 == _T_15 ? ram_227 : _GEN_4429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4431 = 10'he4 == _T_15 ? ram_228 : _GEN_4430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4432 = 10'he5 == _T_15 ? ram_229 : _GEN_4431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4433 = 10'he6 == _T_15 ? ram_230 : _GEN_4432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4434 = 10'he7 == _T_15 ? ram_231 : _GEN_4433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4435 = 10'he8 == _T_15 ? ram_232 : _GEN_4434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4436 = 10'he9 == _T_15 ? ram_233 : _GEN_4435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4437 = 10'hea == _T_15 ? ram_234 : _GEN_4436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4438 = 10'heb == _T_15 ? ram_235 : _GEN_4437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4439 = 10'hec == _T_15 ? ram_236 : _GEN_4438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4440 = 10'hed == _T_15 ? ram_237 : _GEN_4439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4441 = 10'hee == _T_15 ? ram_238 : _GEN_4440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4442 = 10'hef == _T_15 ? ram_239 : _GEN_4441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4443 = 10'hf0 == _T_15 ? ram_240 : _GEN_4442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4444 = 10'hf1 == _T_15 ? ram_241 : _GEN_4443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4445 = 10'hf2 == _T_15 ? ram_242 : _GEN_4444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4446 = 10'hf3 == _T_15 ? ram_243 : _GEN_4445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4447 = 10'hf4 == _T_15 ? ram_244 : _GEN_4446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4448 = 10'hf5 == _T_15 ? ram_245 : _GEN_4447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4449 = 10'hf6 == _T_15 ? ram_246 : _GEN_4448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4450 = 10'hf7 == _T_15 ? ram_247 : _GEN_4449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4451 = 10'hf8 == _T_15 ? ram_248 : _GEN_4450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4452 = 10'hf9 == _T_15 ? ram_249 : _GEN_4451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4453 = 10'hfa == _T_15 ? ram_250 : _GEN_4452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4454 = 10'hfb == _T_15 ? ram_251 : _GEN_4453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4455 = 10'hfc == _T_15 ? ram_252 : _GEN_4454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4456 = 10'hfd == _T_15 ? ram_253 : _GEN_4455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4457 = 10'hfe == _T_15 ? ram_254 : _GEN_4456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4458 = 10'hff == _T_15 ? ram_255 : _GEN_4457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4459 = 10'h100 == _T_15 ? ram_256 : _GEN_4458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4460 = 10'h101 == _T_15 ? ram_257 : _GEN_4459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4461 = 10'h102 == _T_15 ? ram_258 : _GEN_4460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4462 = 10'h103 == _T_15 ? ram_259 : _GEN_4461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4463 = 10'h104 == _T_15 ? ram_260 : _GEN_4462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4464 = 10'h105 == _T_15 ? ram_261 : _GEN_4463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4465 = 10'h106 == _T_15 ? ram_262 : _GEN_4464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4466 = 10'h107 == _T_15 ? ram_263 : _GEN_4465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4467 = 10'h108 == _T_15 ? ram_264 : _GEN_4466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4468 = 10'h109 == _T_15 ? ram_265 : _GEN_4467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4469 = 10'h10a == _T_15 ? ram_266 : _GEN_4468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4470 = 10'h10b == _T_15 ? ram_267 : _GEN_4469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4471 = 10'h10c == _T_15 ? ram_268 : _GEN_4470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4472 = 10'h10d == _T_15 ? ram_269 : _GEN_4471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4473 = 10'h10e == _T_15 ? ram_270 : _GEN_4472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4474 = 10'h10f == _T_15 ? ram_271 : _GEN_4473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4475 = 10'h110 == _T_15 ? ram_272 : _GEN_4474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4476 = 10'h111 == _T_15 ? ram_273 : _GEN_4475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4477 = 10'h112 == _T_15 ? ram_274 : _GEN_4476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4478 = 10'h113 == _T_15 ? ram_275 : _GEN_4477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4479 = 10'h114 == _T_15 ? ram_276 : _GEN_4478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4480 = 10'h115 == _T_15 ? ram_277 : _GEN_4479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4481 = 10'h116 == _T_15 ? ram_278 : _GEN_4480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4482 = 10'h117 == _T_15 ? ram_279 : _GEN_4481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4483 = 10'h118 == _T_15 ? ram_280 : _GEN_4482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4484 = 10'h119 == _T_15 ? ram_281 : _GEN_4483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4485 = 10'h11a == _T_15 ? ram_282 : _GEN_4484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4486 = 10'h11b == _T_15 ? ram_283 : _GEN_4485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4487 = 10'h11c == _T_15 ? ram_284 : _GEN_4486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4488 = 10'h11d == _T_15 ? ram_285 : _GEN_4487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4489 = 10'h11e == _T_15 ? ram_286 : _GEN_4488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4490 = 10'h11f == _T_15 ? ram_287 : _GEN_4489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4491 = 10'h120 == _T_15 ? ram_288 : _GEN_4490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4492 = 10'h121 == _T_15 ? ram_289 : _GEN_4491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4493 = 10'h122 == _T_15 ? ram_290 : _GEN_4492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4494 = 10'h123 == _T_15 ? ram_291 : _GEN_4493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4495 = 10'h124 == _T_15 ? ram_292 : _GEN_4494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4496 = 10'h125 == _T_15 ? ram_293 : _GEN_4495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4497 = 10'h126 == _T_15 ? ram_294 : _GEN_4496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4498 = 10'h127 == _T_15 ? ram_295 : _GEN_4497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4499 = 10'h128 == _T_15 ? ram_296 : _GEN_4498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4500 = 10'h129 == _T_15 ? ram_297 : _GEN_4499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4501 = 10'h12a == _T_15 ? ram_298 : _GEN_4500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4502 = 10'h12b == _T_15 ? ram_299 : _GEN_4501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4503 = 10'h12c == _T_15 ? ram_300 : _GEN_4502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4504 = 10'h12d == _T_15 ? ram_301 : _GEN_4503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4505 = 10'h12e == _T_15 ? ram_302 : _GEN_4504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4506 = 10'h12f == _T_15 ? ram_303 : _GEN_4505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4507 = 10'h130 == _T_15 ? ram_304 : _GEN_4506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4508 = 10'h131 == _T_15 ? ram_305 : _GEN_4507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4509 = 10'h132 == _T_15 ? ram_306 : _GEN_4508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4510 = 10'h133 == _T_15 ? ram_307 : _GEN_4509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4511 = 10'h134 == _T_15 ? ram_308 : _GEN_4510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4512 = 10'h135 == _T_15 ? ram_309 : _GEN_4511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4513 = 10'h136 == _T_15 ? ram_310 : _GEN_4512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4514 = 10'h137 == _T_15 ? ram_311 : _GEN_4513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4515 = 10'h138 == _T_15 ? ram_312 : _GEN_4514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4516 = 10'h139 == _T_15 ? ram_313 : _GEN_4515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4517 = 10'h13a == _T_15 ? ram_314 : _GEN_4516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4518 = 10'h13b == _T_15 ? ram_315 : _GEN_4517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4519 = 10'h13c == _T_15 ? ram_316 : _GEN_4518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4520 = 10'h13d == _T_15 ? ram_317 : _GEN_4519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4521 = 10'h13e == _T_15 ? ram_318 : _GEN_4520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4522 = 10'h13f == _T_15 ? ram_319 : _GEN_4521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4523 = 10'h140 == _T_15 ? ram_320 : _GEN_4522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4524 = 10'h141 == _T_15 ? ram_321 : _GEN_4523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4525 = 10'h142 == _T_15 ? ram_322 : _GEN_4524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4526 = 10'h143 == _T_15 ? ram_323 : _GEN_4525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4527 = 10'h144 == _T_15 ? ram_324 : _GEN_4526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4528 = 10'h145 == _T_15 ? ram_325 : _GEN_4527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4529 = 10'h146 == _T_15 ? ram_326 : _GEN_4528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4530 = 10'h147 == _T_15 ? ram_327 : _GEN_4529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4531 = 10'h148 == _T_15 ? ram_328 : _GEN_4530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4532 = 10'h149 == _T_15 ? ram_329 : _GEN_4531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4533 = 10'h14a == _T_15 ? ram_330 : _GEN_4532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4534 = 10'h14b == _T_15 ? ram_331 : _GEN_4533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4535 = 10'h14c == _T_15 ? ram_332 : _GEN_4534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4536 = 10'h14d == _T_15 ? ram_333 : _GEN_4535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4537 = 10'h14e == _T_15 ? ram_334 : _GEN_4536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4538 = 10'h14f == _T_15 ? ram_335 : _GEN_4537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4539 = 10'h150 == _T_15 ? ram_336 : _GEN_4538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4540 = 10'h151 == _T_15 ? ram_337 : _GEN_4539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4541 = 10'h152 == _T_15 ? ram_338 : _GEN_4540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4542 = 10'h153 == _T_15 ? ram_339 : _GEN_4541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4543 = 10'h154 == _T_15 ? ram_340 : _GEN_4542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4544 = 10'h155 == _T_15 ? ram_341 : _GEN_4543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4545 = 10'h156 == _T_15 ? ram_342 : _GEN_4544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4546 = 10'h157 == _T_15 ? ram_343 : _GEN_4545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4547 = 10'h158 == _T_15 ? ram_344 : _GEN_4546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4548 = 10'h159 == _T_15 ? ram_345 : _GEN_4547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4549 = 10'h15a == _T_15 ? ram_346 : _GEN_4548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4550 = 10'h15b == _T_15 ? ram_347 : _GEN_4549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4551 = 10'h15c == _T_15 ? ram_348 : _GEN_4550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4552 = 10'h15d == _T_15 ? ram_349 : _GEN_4551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4553 = 10'h15e == _T_15 ? ram_350 : _GEN_4552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4554 = 10'h15f == _T_15 ? ram_351 : _GEN_4553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4555 = 10'h160 == _T_15 ? ram_352 : _GEN_4554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4556 = 10'h161 == _T_15 ? ram_353 : _GEN_4555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4557 = 10'h162 == _T_15 ? ram_354 : _GEN_4556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4558 = 10'h163 == _T_15 ? ram_355 : _GEN_4557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4559 = 10'h164 == _T_15 ? ram_356 : _GEN_4558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4560 = 10'h165 == _T_15 ? ram_357 : _GEN_4559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4561 = 10'h166 == _T_15 ? ram_358 : _GEN_4560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4562 = 10'h167 == _T_15 ? ram_359 : _GEN_4561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4563 = 10'h168 == _T_15 ? ram_360 : _GEN_4562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4564 = 10'h169 == _T_15 ? ram_361 : _GEN_4563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4565 = 10'h16a == _T_15 ? ram_362 : _GEN_4564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4566 = 10'h16b == _T_15 ? ram_363 : _GEN_4565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4567 = 10'h16c == _T_15 ? ram_364 : _GEN_4566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4568 = 10'h16d == _T_15 ? ram_365 : _GEN_4567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4569 = 10'h16e == _T_15 ? ram_366 : _GEN_4568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4570 = 10'h16f == _T_15 ? ram_367 : _GEN_4569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4571 = 10'h170 == _T_15 ? ram_368 : _GEN_4570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4572 = 10'h171 == _T_15 ? ram_369 : _GEN_4571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4573 = 10'h172 == _T_15 ? ram_370 : _GEN_4572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4574 = 10'h173 == _T_15 ? ram_371 : _GEN_4573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4575 = 10'h174 == _T_15 ? ram_372 : _GEN_4574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4576 = 10'h175 == _T_15 ? ram_373 : _GEN_4575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4577 = 10'h176 == _T_15 ? ram_374 : _GEN_4576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4578 = 10'h177 == _T_15 ? ram_375 : _GEN_4577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4579 = 10'h178 == _T_15 ? ram_376 : _GEN_4578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4580 = 10'h179 == _T_15 ? ram_377 : _GEN_4579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4581 = 10'h17a == _T_15 ? ram_378 : _GEN_4580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4582 = 10'h17b == _T_15 ? ram_379 : _GEN_4581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4583 = 10'h17c == _T_15 ? ram_380 : _GEN_4582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4584 = 10'h17d == _T_15 ? ram_381 : _GEN_4583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4585 = 10'h17e == _T_15 ? ram_382 : _GEN_4584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4586 = 10'h17f == _T_15 ? ram_383 : _GEN_4585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4587 = 10'h180 == _T_15 ? ram_384 : _GEN_4586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4588 = 10'h181 == _T_15 ? ram_385 : _GEN_4587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4589 = 10'h182 == _T_15 ? ram_386 : _GEN_4588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4590 = 10'h183 == _T_15 ? ram_387 : _GEN_4589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4591 = 10'h184 == _T_15 ? ram_388 : _GEN_4590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4592 = 10'h185 == _T_15 ? ram_389 : _GEN_4591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4593 = 10'h186 == _T_15 ? ram_390 : _GEN_4592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4594 = 10'h187 == _T_15 ? ram_391 : _GEN_4593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4595 = 10'h188 == _T_15 ? ram_392 : _GEN_4594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4596 = 10'h189 == _T_15 ? ram_393 : _GEN_4595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4597 = 10'h18a == _T_15 ? ram_394 : _GEN_4596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4598 = 10'h18b == _T_15 ? ram_395 : _GEN_4597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4599 = 10'h18c == _T_15 ? ram_396 : _GEN_4598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4600 = 10'h18d == _T_15 ? ram_397 : _GEN_4599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4601 = 10'h18e == _T_15 ? ram_398 : _GEN_4600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4602 = 10'h18f == _T_15 ? ram_399 : _GEN_4601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4603 = 10'h190 == _T_15 ? ram_400 : _GEN_4602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4604 = 10'h191 == _T_15 ? ram_401 : _GEN_4603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4605 = 10'h192 == _T_15 ? ram_402 : _GEN_4604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4606 = 10'h193 == _T_15 ? ram_403 : _GEN_4605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4607 = 10'h194 == _T_15 ? ram_404 : _GEN_4606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4608 = 10'h195 == _T_15 ? ram_405 : _GEN_4607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4609 = 10'h196 == _T_15 ? ram_406 : _GEN_4608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4610 = 10'h197 == _T_15 ? ram_407 : _GEN_4609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4611 = 10'h198 == _T_15 ? ram_408 : _GEN_4610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4612 = 10'h199 == _T_15 ? ram_409 : _GEN_4611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4613 = 10'h19a == _T_15 ? ram_410 : _GEN_4612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4614 = 10'h19b == _T_15 ? ram_411 : _GEN_4613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4615 = 10'h19c == _T_15 ? ram_412 : _GEN_4614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4616 = 10'h19d == _T_15 ? ram_413 : _GEN_4615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4617 = 10'h19e == _T_15 ? ram_414 : _GEN_4616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4618 = 10'h19f == _T_15 ? ram_415 : _GEN_4617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4619 = 10'h1a0 == _T_15 ? ram_416 : _GEN_4618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4620 = 10'h1a1 == _T_15 ? ram_417 : _GEN_4619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4621 = 10'h1a2 == _T_15 ? ram_418 : _GEN_4620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4622 = 10'h1a3 == _T_15 ? ram_419 : _GEN_4621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4623 = 10'h1a4 == _T_15 ? ram_420 : _GEN_4622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4624 = 10'h1a5 == _T_15 ? ram_421 : _GEN_4623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4625 = 10'h1a6 == _T_15 ? ram_422 : _GEN_4624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4626 = 10'h1a7 == _T_15 ? ram_423 : _GEN_4625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4627 = 10'h1a8 == _T_15 ? ram_424 : _GEN_4626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4628 = 10'h1a9 == _T_15 ? ram_425 : _GEN_4627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4629 = 10'h1aa == _T_15 ? ram_426 : _GEN_4628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4630 = 10'h1ab == _T_15 ? ram_427 : _GEN_4629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4631 = 10'h1ac == _T_15 ? ram_428 : _GEN_4630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4632 = 10'h1ad == _T_15 ? ram_429 : _GEN_4631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4633 = 10'h1ae == _T_15 ? ram_430 : _GEN_4632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4634 = 10'h1af == _T_15 ? ram_431 : _GEN_4633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4635 = 10'h1b0 == _T_15 ? ram_432 : _GEN_4634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4636 = 10'h1b1 == _T_15 ? ram_433 : _GEN_4635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4637 = 10'h1b2 == _T_15 ? ram_434 : _GEN_4636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4638 = 10'h1b3 == _T_15 ? ram_435 : _GEN_4637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4639 = 10'h1b4 == _T_15 ? ram_436 : _GEN_4638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4640 = 10'h1b5 == _T_15 ? ram_437 : _GEN_4639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4641 = 10'h1b6 == _T_15 ? ram_438 : _GEN_4640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4642 = 10'h1b7 == _T_15 ? ram_439 : _GEN_4641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4643 = 10'h1b8 == _T_15 ? ram_440 : _GEN_4642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4644 = 10'h1b9 == _T_15 ? ram_441 : _GEN_4643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4645 = 10'h1ba == _T_15 ? ram_442 : _GEN_4644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4646 = 10'h1bb == _T_15 ? ram_443 : _GEN_4645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4647 = 10'h1bc == _T_15 ? ram_444 : _GEN_4646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4648 = 10'h1bd == _T_15 ? ram_445 : _GEN_4647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4649 = 10'h1be == _T_15 ? ram_446 : _GEN_4648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4650 = 10'h1bf == _T_15 ? ram_447 : _GEN_4649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4651 = 10'h1c0 == _T_15 ? ram_448 : _GEN_4650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4652 = 10'h1c1 == _T_15 ? ram_449 : _GEN_4651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4653 = 10'h1c2 == _T_15 ? ram_450 : _GEN_4652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4654 = 10'h1c3 == _T_15 ? ram_451 : _GEN_4653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4655 = 10'h1c4 == _T_15 ? ram_452 : _GEN_4654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4656 = 10'h1c5 == _T_15 ? ram_453 : _GEN_4655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4657 = 10'h1c6 == _T_15 ? ram_454 : _GEN_4656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4658 = 10'h1c7 == _T_15 ? ram_455 : _GEN_4657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4659 = 10'h1c8 == _T_15 ? ram_456 : _GEN_4658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4660 = 10'h1c9 == _T_15 ? ram_457 : _GEN_4659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4661 = 10'h1ca == _T_15 ? ram_458 : _GEN_4660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4662 = 10'h1cb == _T_15 ? ram_459 : _GEN_4661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4663 = 10'h1cc == _T_15 ? ram_460 : _GEN_4662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4664 = 10'h1cd == _T_15 ? ram_461 : _GEN_4663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4665 = 10'h1ce == _T_15 ? ram_462 : _GEN_4664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4666 = 10'h1cf == _T_15 ? ram_463 : _GEN_4665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4667 = 10'h1d0 == _T_15 ? ram_464 : _GEN_4666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4668 = 10'h1d1 == _T_15 ? ram_465 : _GEN_4667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4669 = 10'h1d2 == _T_15 ? ram_466 : _GEN_4668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4670 = 10'h1d3 == _T_15 ? ram_467 : _GEN_4669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4671 = 10'h1d4 == _T_15 ? ram_468 : _GEN_4670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4672 = 10'h1d5 == _T_15 ? ram_469 : _GEN_4671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4673 = 10'h1d6 == _T_15 ? ram_470 : _GEN_4672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4674 = 10'h1d7 == _T_15 ? ram_471 : _GEN_4673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4675 = 10'h1d8 == _T_15 ? ram_472 : _GEN_4674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4676 = 10'h1d9 == _T_15 ? ram_473 : _GEN_4675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4677 = 10'h1da == _T_15 ? ram_474 : _GEN_4676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4678 = 10'h1db == _T_15 ? ram_475 : _GEN_4677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4679 = 10'h1dc == _T_15 ? ram_476 : _GEN_4678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4680 = 10'h1dd == _T_15 ? ram_477 : _GEN_4679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4681 = 10'h1de == _T_15 ? ram_478 : _GEN_4680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4682 = 10'h1df == _T_15 ? ram_479 : _GEN_4681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4683 = 10'h1e0 == _T_15 ? ram_480 : _GEN_4682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4684 = 10'h1e1 == _T_15 ? ram_481 : _GEN_4683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4685 = 10'h1e2 == _T_15 ? ram_482 : _GEN_4684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4686 = 10'h1e3 == _T_15 ? ram_483 : _GEN_4685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4687 = 10'h1e4 == _T_15 ? ram_484 : _GEN_4686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4688 = 10'h1e5 == _T_15 ? ram_485 : _GEN_4687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4689 = 10'h1e6 == _T_15 ? ram_486 : _GEN_4688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4690 = 10'h1e7 == _T_15 ? ram_487 : _GEN_4689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4691 = 10'h1e8 == _T_15 ? ram_488 : _GEN_4690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4692 = 10'h1e9 == _T_15 ? ram_489 : _GEN_4691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4693 = 10'h1ea == _T_15 ? ram_490 : _GEN_4692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4694 = 10'h1eb == _T_15 ? ram_491 : _GEN_4693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4695 = 10'h1ec == _T_15 ? ram_492 : _GEN_4694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4696 = 10'h1ed == _T_15 ? ram_493 : _GEN_4695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4697 = 10'h1ee == _T_15 ? ram_494 : _GEN_4696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4698 = 10'h1ef == _T_15 ? ram_495 : _GEN_4697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4699 = 10'h1f0 == _T_15 ? ram_496 : _GEN_4698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4700 = 10'h1f1 == _T_15 ? ram_497 : _GEN_4699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4701 = 10'h1f2 == _T_15 ? ram_498 : _GEN_4700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4702 = 10'h1f3 == _T_15 ? ram_499 : _GEN_4701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4703 = 10'h1f4 == _T_15 ? ram_500 : _GEN_4702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4704 = 10'h1f5 == _T_15 ? ram_501 : _GEN_4703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4705 = 10'h1f6 == _T_15 ? ram_502 : _GEN_4704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4706 = 10'h1f7 == _T_15 ? ram_503 : _GEN_4705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4707 = 10'h1f8 == _T_15 ? ram_504 : _GEN_4706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4708 = 10'h1f9 == _T_15 ? ram_505 : _GEN_4707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4709 = 10'h1fa == _T_15 ? ram_506 : _GEN_4708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4710 = 10'h1fb == _T_15 ? ram_507 : _GEN_4709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4711 = 10'h1fc == _T_15 ? ram_508 : _GEN_4710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4712 = 10'h1fd == _T_15 ? ram_509 : _GEN_4711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4713 = 10'h1fe == _T_15 ? ram_510 : _GEN_4712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4714 = 10'h1ff == _T_15 ? ram_511 : _GEN_4713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4715 = 10'h200 == _T_15 ? ram_512 : _GEN_4714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4716 = 10'h201 == _T_15 ? ram_513 : _GEN_4715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4717 = 10'h202 == _T_15 ? ram_514 : _GEN_4716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4718 = 10'h203 == _T_15 ? ram_515 : _GEN_4717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4719 = 10'h204 == _T_15 ? ram_516 : _GEN_4718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4720 = 10'h205 == _T_15 ? ram_517 : _GEN_4719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4721 = 10'h206 == _T_15 ? ram_518 : _GEN_4720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4722 = 10'h207 == _T_15 ? ram_519 : _GEN_4721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4723 = 10'h208 == _T_15 ? ram_520 : _GEN_4722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4724 = 10'h209 == _T_15 ? ram_521 : _GEN_4723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4725 = 10'h20a == _T_15 ? ram_522 : _GEN_4724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4726 = 10'h20b == _T_15 ? ram_523 : _GEN_4725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_4727 = 10'h20c == _T_15 ? ram_524 : _GEN_4726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19069 = {{8190'd0}, _GEN_4727}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_129 = _GEN_19069 ^ _ram_T_128; // @[vga.scala 64:41]
  wire [287:0] _GEN_4728 = 10'h0 == _T_15 ? _ram_T_129[287:0] : _GEN_3678; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4729 = 10'h1 == _T_15 ? _ram_T_129[287:0] : _GEN_3679; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4730 = 10'h2 == _T_15 ? _ram_T_129[287:0] : _GEN_3680; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4731 = 10'h3 == _T_15 ? _ram_T_129[287:0] : _GEN_3681; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4732 = 10'h4 == _T_15 ? _ram_T_129[287:0] : _GEN_3682; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4733 = 10'h5 == _T_15 ? _ram_T_129[287:0] : _GEN_3683; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4734 = 10'h6 == _T_15 ? _ram_T_129[287:0] : _GEN_3684; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4735 = 10'h7 == _T_15 ? _ram_T_129[287:0] : _GEN_3685; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4736 = 10'h8 == _T_15 ? _ram_T_129[287:0] : _GEN_3686; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4737 = 10'h9 == _T_15 ? _ram_T_129[287:0] : _GEN_3687; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4738 = 10'ha == _T_15 ? _ram_T_129[287:0] : _GEN_3688; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4739 = 10'hb == _T_15 ? _ram_T_129[287:0] : _GEN_3689; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4740 = 10'hc == _T_15 ? _ram_T_129[287:0] : _GEN_3690; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4741 = 10'hd == _T_15 ? _ram_T_129[287:0] : _GEN_3691; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4742 = 10'he == _T_15 ? _ram_T_129[287:0] : _GEN_3692; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4743 = 10'hf == _T_15 ? _ram_T_129[287:0] : _GEN_3693; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4744 = 10'h10 == _T_15 ? _ram_T_129[287:0] : _GEN_3694; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4745 = 10'h11 == _T_15 ? _ram_T_129[287:0] : _GEN_3695; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4746 = 10'h12 == _T_15 ? _ram_T_129[287:0] : _GEN_3696; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4747 = 10'h13 == _T_15 ? _ram_T_129[287:0] : _GEN_3697; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4748 = 10'h14 == _T_15 ? _ram_T_129[287:0] : _GEN_3698; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4749 = 10'h15 == _T_15 ? _ram_T_129[287:0] : _GEN_3699; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4750 = 10'h16 == _T_15 ? _ram_T_129[287:0] : _GEN_3700; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4751 = 10'h17 == _T_15 ? _ram_T_129[287:0] : _GEN_3701; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4752 = 10'h18 == _T_15 ? _ram_T_129[287:0] : _GEN_3702; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4753 = 10'h19 == _T_15 ? _ram_T_129[287:0] : _GEN_3703; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4754 = 10'h1a == _T_15 ? _ram_T_129[287:0] : _GEN_3704; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4755 = 10'h1b == _T_15 ? _ram_T_129[287:0] : _GEN_3705; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4756 = 10'h1c == _T_15 ? _ram_T_129[287:0] : _GEN_3706; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4757 = 10'h1d == _T_15 ? _ram_T_129[287:0] : _GEN_3707; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4758 = 10'h1e == _T_15 ? _ram_T_129[287:0] : _GEN_3708; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4759 = 10'h1f == _T_15 ? _ram_T_129[287:0] : _GEN_3709; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4760 = 10'h20 == _T_15 ? _ram_T_129[287:0] : _GEN_3710; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4761 = 10'h21 == _T_15 ? _ram_T_129[287:0] : _GEN_3711; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4762 = 10'h22 == _T_15 ? _ram_T_129[287:0] : _GEN_3712; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4763 = 10'h23 == _T_15 ? _ram_T_129[287:0] : _GEN_3713; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4764 = 10'h24 == _T_15 ? _ram_T_129[287:0] : _GEN_3714; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4765 = 10'h25 == _T_15 ? _ram_T_129[287:0] : _GEN_3715; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4766 = 10'h26 == _T_15 ? _ram_T_129[287:0] : _GEN_3716; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4767 = 10'h27 == _T_15 ? _ram_T_129[287:0] : _GEN_3717; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4768 = 10'h28 == _T_15 ? _ram_T_129[287:0] : _GEN_3718; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4769 = 10'h29 == _T_15 ? _ram_T_129[287:0] : _GEN_3719; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4770 = 10'h2a == _T_15 ? _ram_T_129[287:0] : _GEN_3720; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4771 = 10'h2b == _T_15 ? _ram_T_129[287:0] : _GEN_3721; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4772 = 10'h2c == _T_15 ? _ram_T_129[287:0] : _GEN_3722; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4773 = 10'h2d == _T_15 ? _ram_T_129[287:0] : _GEN_3723; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4774 = 10'h2e == _T_15 ? _ram_T_129[287:0] : _GEN_3724; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4775 = 10'h2f == _T_15 ? _ram_T_129[287:0] : _GEN_3725; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4776 = 10'h30 == _T_15 ? _ram_T_129[287:0] : _GEN_3726; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4777 = 10'h31 == _T_15 ? _ram_T_129[287:0] : _GEN_3727; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4778 = 10'h32 == _T_15 ? _ram_T_129[287:0] : _GEN_3728; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4779 = 10'h33 == _T_15 ? _ram_T_129[287:0] : _GEN_3729; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4780 = 10'h34 == _T_15 ? _ram_T_129[287:0] : _GEN_3730; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4781 = 10'h35 == _T_15 ? _ram_T_129[287:0] : _GEN_3731; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4782 = 10'h36 == _T_15 ? _ram_T_129[287:0] : _GEN_3732; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4783 = 10'h37 == _T_15 ? _ram_T_129[287:0] : _GEN_3733; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4784 = 10'h38 == _T_15 ? _ram_T_129[287:0] : _GEN_3734; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4785 = 10'h39 == _T_15 ? _ram_T_129[287:0] : _GEN_3735; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4786 = 10'h3a == _T_15 ? _ram_T_129[287:0] : _GEN_3736; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4787 = 10'h3b == _T_15 ? _ram_T_129[287:0] : _GEN_3737; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4788 = 10'h3c == _T_15 ? _ram_T_129[287:0] : _GEN_3738; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4789 = 10'h3d == _T_15 ? _ram_T_129[287:0] : _GEN_3739; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4790 = 10'h3e == _T_15 ? _ram_T_129[287:0] : _GEN_3740; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4791 = 10'h3f == _T_15 ? _ram_T_129[287:0] : _GEN_3741; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4792 = 10'h40 == _T_15 ? _ram_T_129[287:0] : _GEN_3742; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4793 = 10'h41 == _T_15 ? _ram_T_129[287:0] : _GEN_3743; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4794 = 10'h42 == _T_15 ? _ram_T_129[287:0] : _GEN_3744; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4795 = 10'h43 == _T_15 ? _ram_T_129[287:0] : _GEN_3745; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4796 = 10'h44 == _T_15 ? _ram_T_129[287:0] : _GEN_3746; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4797 = 10'h45 == _T_15 ? _ram_T_129[287:0] : _GEN_3747; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4798 = 10'h46 == _T_15 ? _ram_T_129[287:0] : _GEN_3748; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4799 = 10'h47 == _T_15 ? _ram_T_129[287:0] : _GEN_3749; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4800 = 10'h48 == _T_15 ? _ram_T_129[287:0] : _GEN_3750; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4801 = 10'h49 == _T_15 ? _ram_T_129[287:0] : _GEN_3751; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4802 = 10'h4a == _T_15 ? _ram_T_129[287:0] : _GEN_3752; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4803 = 10'h4b == _T_15 ? _ram_T_129[287:0] : _GEN_3753; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4804 = 10'h4c == _T_15 ? _ram_T_129[287:0] : _GEN_3754; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4805 = 10'h4d == _T_15 ? _ram_T_129[287:0] : _GEN_3755; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4806 = 10'h4e == _T_15 ? _ram_T_129[287:0] : _GEN_3756; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4807 = 10'h4f == _T_15 ? _ram_T_129[287:0] : _GEN_3757; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4808 = 10'h50 == _T_15 ? _ram_T_129[287:0] : _GEN_3758; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4809 = 10'h51 == _T_15 ? _ram_T_129[287:0] : _GEN_3759; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4810 = 10'h52 == _T_15 ? _ram_T_129[287:0] : _GEN_3760; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4811 = 10'h53 == _T_15 ? _ram_T_129[287:0] : _GEN_3761; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4812 = 10'h54 == _T_15 ? _ram_T_129[287:0] : _GEN_3762; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4813 = 10'h55 == _T_15 ? _ram_T_129[287:0] : _GEN_3763; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4814 = 10'h56 == _T_15 ? _ram_T_129[287:0] : _GEN_3764; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4815 = 10'h57 == _T_15 ? _ram_T_129[287:0] : _GEN_3765; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4816 = 10'h58 == _T_15 ? _ram_T_129[287:0] : _GEN_3766; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4817 = 10'h59 == _T_15 ? _ram_T_129[287:0] : _GEN_3767; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4818 = 10'h5a == _T_15 ? _ram_T_129[287:0] : _GEN_3768; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4819 = 10'h5b == _T_15 ? _ram_T_129[287:0] : _GEN_3769; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4820 = 10'h5c == _T_15 ? _ram_T_129[287:0] : _GEN_3770; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4821 = 10'h5d == _T_15 ? _ram_T_129[287:0] : _GEN_3771; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4822 = 10'h5e == _T_15 ? _ram_T_129[287:0] : _GEN_3772; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4823 = 10'h5f == _T_15 ? _ram_T_129[287:0] : _GEN_3773; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4824 = 10'h60 == _T_15 ? _ram_T_129[287:0] : _GEN_3774; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4825 = 10'h61 == _T_15 ? _ram_T_129[287:0] : _GEN_3775; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4826 = 10'h62 == _T_15 ? _ram_T_129[287:0] : _GEN_3776; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4827 = 10'h63 == _T_15 ? _ram_T_129[287:0] : _GEN_3777; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4828 = 10'h64 == _T_15 ? _ram_T_129[287:0] : _GEN_3778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4829 = 10'h65 == _T_15 ? _ram_T_129[287:0] : _GEN_3779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4830 = 10'h66 == _T_15 ? _ram_T_129[287:0] : _GEN_3780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4831 = 10'h67 == _T_15 ? _ram_T_129[287:0] : _GEN_3781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4832 = 10'h68 == _T_15 ? _ram_T_129[287:0] : _GEN_3782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4833 = 10'h69 == _T_15 ? _ram_T_129[287:0] : _GEN_3783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4834 = 10'h6a == _T_15 ? _ram_T_129[287:0] : _GEN_3784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4835 = 10'h6b == _T_15 ? _ram_T_129[287:0] : _GEN_3785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4836 = 10'h6c == _T_15 ? _ram_T_129[287:0] : _GEN_3786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4837 = 10'h6d == _T_15 ? _ram_T_129[287:0] : _GEN_3787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4838 = 10'h6e == _T_15 ? _ram_T_129[287:0] : _GEN_3788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4839 = 10'h6f == _T_15 ? _ram_T_129[287:0] : _GEN_3789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4840 = 10'h70 == _T_15 ? _ram_T_129[287:0] : _GEN_3790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4841 = 10'h71 == _T_15 ? _ram_T_129[287:0] : _GEN_3791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4842 = 10'h72 == _T_15 ? _ram_T_129[287:0] : _GEN_3792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4843 = 10'h73 == _T_15 ? _ram_T_129[287:0] : _GEN_3793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4844 = 10'h74 == _T_15 ? _ram_T_129[287:0] : _GEN_3794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4845 = 10'h75 == _T_15 ? _ram_T_129[287:0] : _GEN_3795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4846 = 10'h76 == _T_15 ? _ram_T_129[287:0] : _GEN_3796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4847 = 10'h77 == _T_15 ? _ram_T_129[287:0] : _GEN_3797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4848 = 10'h78 == _T_15 ? _ram_T_129[287:0] : _GEN_3798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4849 = 10'h79 == _T_15 ? _ram_T_129[287:0] : _GEN_3799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4850 = 10'h7a == _T_15 ? _ram_T_129[287:0] : _GEN_3800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4851 = 10'h7b == _T_15 ? _ram_T_129[287:0] : _GEN_3801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4852 = 10'h7c == _T_15 ? _ram_T_129[287:0] : _GEN_3802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4853 = 10'h7d == _T_15 ? _ram_T_129[287:0] : _GEN_3803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4854 = 10'h7e == _T_15 ? _ram_T_129[287:0] : _GEN_3804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4855 = 10'h7f == _T_15 ? _ram_T_129[287:0] : _GEN_3805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4856 = 10'h80 == _T_15 ? _ram_T_129[287:0] : _GEN_3806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4857 = 10'h81 == _T_15 ? _ram_T_129[287:0] : _GEN_3807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4858 = 10'h82 == _T_15 ? _ram_T_129[287:0] : _GEN_3808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4859 = 10'h83 == _T_15 ? _ram_T_129[287:0] : _GEN_3809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4860 = 10'h84 == _T_15 ? _ram_T_129[287:0] : _GEN_3810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4861 = 10'h85 == _T_15 ? _ram_T_129[287:0] : _GEN_3811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4862 = 10'h86 == _T_15 ? _ram_T_129[287:0] : _GEN_3812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4863 = 10'h87 == _T_15 ? _ram_T_129[287:0] : _GEN_3813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4864 = 10'h88 == _T_15 ? _ram_T_129[287:0] : _GEN_3814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4865 = 10'h89 == _T_15 ? _ram_T_129[287:0] : _GEN_3815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4866 = 10'h8a == _T_15 ? _ram_T_129[287:0] : _GEN_3816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4867 = 10'h8b == _T_15 ? _ram_T_129[287:0] : _GEN_3817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4868 = 10'h8c == _T_15 ? _ram_T_129[287:0] : _GEN_3818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4869 = 10'h8d == _T_15 ? _ram_T_129[287:0] : _GEN_3819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4870 = 10'h8e == _T_15 ? _ram_T_129[287:0] : _GEN_3820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4871 = 10'h8f == _T_15 ? _ram_T_129[287:0] : _GEN_3821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4872 = 10'h90 == _T_15 ? _ram_T_129[287:0] : _GEN_3822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4873 = 10'h91 == _T_15 ? _ram_T_129[287:0] : _GEN_3823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4874 = 10'h92 == _T_15 ? _ram_T_129[287:0] : _GEN_3824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4875 = 10'h93 == _T_15 ? _ram_T_129[287:0] : _GEN_3825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4876 = 10'h94 == _T_15 ? _ram_T_129[287:0] : _GEN_3826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4877 = 10'h95 == _T_15 ? _ram_T_129[287:0] : _GEN_3827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4878 = 10'h96 == _T_15 ? _ram_T_129[287:0] : _GEN_3828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4879 = 10'h97 == _T_15 ? _ram_T_129[287:0] : _GEN_3829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4880 = 10'h98 == _T_15 ? _ram_T_129[287:0] : _GEN_3830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4881 = 10'h99 == _T_15 ? _ram_T_129[287:0] : _GEN_3831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4882 = 10'h9a == _T_15 ? _ram_T_129[287:0] : _GEN_3832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4883 = 10'h9b == _T_15 ? _ram_T_129[287:0] : _GEN_3833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4884 = 10'h9c == _T_15 ? _ram_T_129[287:0] : _GEN_3834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4885 = 10'h9d == _T_15 ? _ram_T_129[287:0] : _GEN_3835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4886 = 10'h9e == _T_15 ? _ram_T_129[287:0] : _GEN_3836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4887 = 10'h9f == _T_15 ? _ram_T_129[287:0] : _GEN_3837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4888 = 10'ha0 == _T_15 ? _ram_T_129[287:0] : _GEN_3838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4889 = 10'ha1 == _T_15 ? _ram_T_129[287:0] : _GEN_3839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4890 = 10'ha2 == _T_15 ? _ram_T_129[287:0] : _GEN_3840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4891 = 10'ha3 == _T_15 ? _ram_T_129[287:0] : _GEN_3841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4892 = 10'ha4 == _T_15 ? _ram_T_129[287:0] : _GEN_3842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4893 = 10'ha5 == _T_15 ? _ram_T_129[287:0] : _GEN_3843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4894 = 10'ha6 == _T_15 ? _ram_T_129[287:0] : _GEN_3844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4895 = 10'ha7 == _T_15 ? _ram_T_129[287:0] : _GEN_3845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4896 = 10'ha8 == _T_15 ? _ram_T_129[287:0] : _GEN_3846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4897 = 10'ha9 == _T_15 ? _ram_T_129[287:0] : _GEN_3847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4898 = 10'haa == _T_15 ? _ram_T_129[287:0] : _GEN_3848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4899 = 10'hab == _T_15 ? _ram_T_129[287:0] : _GEN_3849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4900 = 10'hac == _T_15 ? _ram_T_129[287:0] : _GEN_3850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4901 = 10'had == _T_15 ? _ram_T_129[287:0] : _GEN_3851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4902 = 10'hae == _T_15 ? _ram_T_129[287:0] : _GEN_3852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4903 = 10'haf == _T_15 ? _ram_T_129[287:0] : _GEN_3853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4904 = 10'hb0 == _T_15 ? _ram_T_129[287:0] : _GEN_3854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4905 = 10'hb1 == _T_15 ? _ram_T_129[287:0] : _GEN_3855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4906 = 10'hb2 == _T_15 ? _ram_T_129[287:0] : _GEN_3856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4907 = 10'hb3 == _T_15 ? _ram_T_129[287:0] : _GEN_3857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4908 = 10'hb4 == _T_15 ? _ram_T_129[287:0] : _GEN_3858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4909 = 10'hb5 == _T_15 ? _ram_T_129[287:0] : _GEN_3859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4910 = 10'hb6 == _T_15 ? _ram_T_129[287:0] : _GEN_3860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4911 = 10'hb7 == _T_15 ? _ram_T_129[287:0] : _GEN_3861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4912 = 10'hb8 == _T_15 ? _ram_T_129[287:0] : _GEN_3862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4913 = 10'hb9 == _T_15 ? _ram_T_129[287:0] : _GEN_3863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4914 = 10'hba == _T_15 ? _ram_T_129[287:0] : _GEN_3864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4915 = 10'hbb == _T_15 ? _ram_T_129[287:0] : _GEN_3865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4916 = 10'hbc == _T_15 ? _ram_T_129[287:0] : _GEN_3866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4917 = 10'hbd == _T_15 ? _ram_T_129[287:0] : _GEN_3867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4918 = 10'hbe == _T_15 ? _ram_T_129[287:0] : _GEN_3868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4919 = 10'hbf == _T_15 ? _ram_T_129[287:0] : _GEN_3869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4920 = 10'hc0 == _T_15 ? _ram_T_129[287:0] : _GEN_3870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4921 = 10'hc1 == _T_15 ? _ram_T_129[287:0] : _GEN_3871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4922 = 10'hc2 == _T_15 ? _ram_T_129[287:0] : _GEN_3872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4923 = 10'hc3 == _T_15 ? _ram_T_129[287:0] : _GEN_3873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4924 = 10'hc4 == _T_15 ? _ram_T_129[287:0] : _GEN_3874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4925 = 10'hc5 == _T_15 ? _ram_T_129[287:0] : _GEN_3875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4926 = 10'hc6 == _T_15 ? _ram_T_129[287:0] : _GEN_3876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4927 = 10'hc7 == _T_15 ? _ram_T_129[287:0] : _GEN_3877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4928 = 10'hc8 == _T_15 ? _ram_T_129[287:0] : _GEN_3878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4929 = 10'hc9 == _T_15 ? _ram_T_129[287:0] : _GEN_3879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4930 = 10'hca == _T_15 ? _ram_T_129[287:0] : _GEN_3880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4931 = 10'hcb == _T_15 ? _ram_T_129[287:0] : _GEN_3881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4932 = 10'hcc == _T_15 ? _ram_T_129[287:0] : _GEN_3882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4933 = 10'hcd == _T_15 ? _ram_T_129[287:0] : _GEN_3883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4934 = 10'hce == _T_15 ? _ram_T_129[287:0] : _GEN_3884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4935 = 10'hcf == _T_15 ? _ram_T_129[287:0] : _GEN_3885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4936 = 10'hd0 == _T_15 ? _ram_T_129[287:0] : _GEN_3886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4937 = 10'hd1 == _T_15 ? _ram_T_129[287:0] : _GEN_3887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4938 = 10'hd2 == _T_15 ? _ram_T_129[287:0] : _GEN_3888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4939 = 10'hd3 == _T_15 ? _ram_T_129[287:0] : _GEN_3889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4940 = 10'hd4 == _T_15 ? _ram_T_129[287:0] : _GEN_3890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4941 = 10'hd5 == _T_15 ? _ram_T_129[287:0] : _GEN_3891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4942 = 10'hd6 == _T_15 ? _ram_T_129[287:0] : _GEN_3892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4943 = 10'hd7 == _T_15 ? _ram_T_129[287:0] : _GEN_3893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4944 = 10'hd8 == _T_15 ? _ram_T_129[287:0] : _GEN_3894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4945 = 10'hd9 == _T_15 ? _ram_T_129[287:0] : _GEN_3895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4946 = 10'hda == _T_15 ? _ram_T_129[287:0] : _GEN_3896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4947 = 10'hdb == _T_15 ? _ram_T_129[287:0] : _GEN_3897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4948 = 10'hdc == _T_15 ? _ram_T_129[287:0] : _GEN_3898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4949 = 10'hdd == _T_15 ? _ram_T_129[287:0] : _GEN_3899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4950 = 10'hde == _T_15 ? _ram_T_129[287:0] : _GEN_3900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4951 = 10'hdf == _T_15 ? _ram_T_129[287:0] : _GEN_3901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4952 = 10'he0 == _T_15 ? _ram_T_129[287:0] : _GEN_3902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4953 = 10'he1 == _T_15 ? _ram_T_129[287:0] : _GEN_3903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4954 = 10'he2 == _T_15 ? _ram_T_129[287:0] : _GEN_3904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4955 = 10'he3 == _T_15 ? _ram_T_129[287:0] : _GEN_3905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4956 = 10'he4 == _T_15 ? _ram_T_129[287:0] : _GEN_3906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4957 = 10'he5 == _T_15 ? _ram_T_129[287:0] : _GEN_3907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4958 = 10'he6 == _T_15 ? _ram_T_129[287:0] : _GEN_3908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4959 = 10'he7 == _T_15 ? _ram_T_129[287:0] : _GEN_3909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4960 = 10'he8 == _T_15 ? _ram_T_129[287:0] : _GEN_3910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4961 = 10'he9 == _T_15 ? _ram_T_129[287:0] : _GEN_3911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4962 = 10'hea == _T_15 ? _ram_T_129[287:0] : _GEN_3912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4963 = 10'heb == _T_15 ? _ram_T_129[287:0] : _GEN_3913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4964 = 10'hec == _T_15 ? _ram_T_129[287:0] : _GEN_3914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4965 = 10'hed == _T_15 ? _ram_T_129[287:0] : _GEN_3915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4966 = 10'hee == _T_15 ? _ram_T_129[287:0] : _GEN_3916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4967 = 10'hef == _T_15 ? _ram_T_129[287:0] : _GEN_3917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4968 = 10'hf0 == _T_15 ? _ram_T_129[287:0] : _GEN_3918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4969 = 10'hf1 == _T_15 ? _ram_T_129[287:0] : _GEN_3919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4970 = 10'hf2 == _T_15 ? _ram_T_129[287:0] : _GEN_3920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4971 = 10'hf3 == _T_15 ? _ram_T_129[287:0] : _GEN_3921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4972 = 10'hf4 == _T_15 ? _ram_T_129[287:0] : _GEN_3922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4973 = 10'hf5 == _T_15 ? _ram_T_129[287:0] : _GEN_3923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4974 = 10'hf6 == _T_15 ? _ram_T_129[287:0] : _GEN_3924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4975 = 10'hf7 == _T_15 ? _ram_T_129[287:0] : _GEN_3925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4976 = 10'hf8 == _T_15 ? _ram_T_129[287:0] : _GEN_3926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4977 = 10'hf9 == _T_15 ? _ram_T_129[287:0] : _GEN_3927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4978 = 10'hfa == _T_15 ? _ram_T_129[287:0] : _GEN_3928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4979 = 10'hfb == _T_15 ? _ram_T_129[287:0] : _GEN_3929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4980 = 10'hfc == _T_15 ? _ram_T_129[287:0] : _GEN_3930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4981 = 10'hfd == _T_15 ? _ram_T_129[287:0] : _GEN_3931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4982 = 10'hfe == _T_15 ? _ram_T_129[287:0] : _GEN_3932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4983 = 10'hff == _T_15 ? _ram_T_129[287:0] : _GEN_3933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4984 = 10'h100 == _T_15 ? _ram_T_129[287:0] : _GEN_3934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4985 = 10'h101 == _T_15 ? _ram_T_129[287:0] : _GEN_3935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4986 = 10'h102 == _T_15 ? _ram_T_129[287:0] : _GEN_3936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4987 = 10'h103 == _T_15 ? _ram_T_129[287:0] : _GEN_3937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4988 = 10'h104 == _T_15 ? _ram_T_129[287:0] : _GEN_3938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4989 = 10'h105 == _T_15 ? _ram_T_129[287:0] : _GEN_3939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4990 = 10'h106 == _T_15 ? _ram_T_129[287:0] : _GEN_3940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4991 = 10'h107 == _T_15 ? _ram_T_129[287:0] : _GEN_3941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4992 = 10'h108 == _T_15 ? _ram_T_129[287:0] : _GEN_3942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4993 = 10'h109 == _T_15 ? _ram_T_129[287:0] : _GEN_3943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4994 = 10'h10a == _T_15 ? _ram_T_129[287:0] : _GEN_3944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4995 = 10'h10b == _T_15 ? _ram_T_129[287:0] : _GEN_3945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4996 = 10'h10c == _T_15 ? _ram_T_129[287:0] : _GEN_3946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4997 = 10'h10d == _T_15 ? _ram_T_129[287:0] : _GEN_3947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4998 = 10'h10e == _T_15 ? _ram_T_129[287:0] : _GEN_3948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_4999 = 10'h10f == _T_15 ? _ram_T_129[287:0] : _GEN_3949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5000 = 10'h110 == _T_15 ? _ram_T_129[287:0] : _GEN_3950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5001 = 10'h111 == _T_15 ? _ram_T_129[287:0] : _GEN_3951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5002 = 10'h112 == _T_15 ? _ram_T_129[287:0] : _GEN_3952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5003 = 10'h113 == _T_15 ? _ram_T_129[287:0] : _GEN_3953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5004 = 10'h114 == _T_15 ? _ram_T_129[287:0] : _GEN_3954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5005 = 10'h115 == _T_15 ? _ram_T_129[287:0] : _GEN_3955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5006 = 10'h116 == _T_15 ? _ram_T_129[287:0] : _GEN_3956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5007 = 10'h117 == _T_15 ? _ram_T_129[287:0] : _GEN_3957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5008 = 10'h118 == _T_15 ? _ram_T_129[287:0] : _GEN_3958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5009 = 10'h119 == _T_15 ? _ram_T_129[287:0] : _GEN_3959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5010 = 10'h11a == _T_15 ? _ram_T_129[287:0] : _GEN_3960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5011 = 10'h11b == _T_15 ? _ram_T_129[287:0] : _GEN_3961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5012 = 10'h11c == _T_15 ? _ram_T_129[287:0] : _GEN_3962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5013 = 10'h11d == _T_15 ? _ram_T_129[287:0] : _GEN_3963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5014 = 10'h11e == _T_15 ? _ram_T_129[287:0] : _GEN_3964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5015 = 10'h11f == _T_15 ? _ram_T_129[287:0] : _GEN_3965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5016 = 10'h120 == _T_15 ? _ram_T_129[287:0] : _GEN_3966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5017 = 10'h121 == _T_15 ? _ram_T_129[287:0] : _GEN_3967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5018 = 10'h122 == _T_15 ? _ram_T_129[287:0] : _GEN_3968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5019 = 10'h123 == _T_15 ? _ram_T_129[287:0] : _GEN_3969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5020 = 10'h124 == _T_15 ? _ram_T_129[287:0] : _GEN_3970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5021 = 10'h125 == _T_15 ? _ram_T_129[287:0] : _GEN_3971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5022 = 10'h126 == _T_15 ? _ram_T_129[287:0] : _GEN_3972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5023 = 10'h127 == _T_15 ? _ram_T_129[287:0] : _GEN_3973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5024 = 10'h128 == _T_15 ? _ram_T_129[287:0] : _GEN_3974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5025 = 10'h129 == _T_15 ? _ram_T_129[287:0] : _GEN_3975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5026 = 10'h12a == _T_15 ? _ram_T_129[287:0] : _GEN_3976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5027 = 10'h12b == _T_15 ? _ram_T_129[287:0] : _GEN_3977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5028 = 10'h12c == _T_15 ? _ram_T_129[287:0] : _GEN_3978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5029 = 10'h12d == _T_15 ? _ram_T_129[287:0] : _GEN_3979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5030 = 10'h12e == _T_15 ? _ram_T_129[287:0] : _GEN_3980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5031 = 10'h12f == _T_15 ? _ram_T_129[287:0] : _GEN_3981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5032 = 10'h130 == _T_15 ? _ram_T_129[287:0] : _GEN_3982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5033 = 10'h131 == _T_15 ? _ram_T_129[287:0] : _GEN_3983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5034 = 10'h132 == _T_15 ? _ram_T_129[287:0] : _GEN_3984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5035 = 10'h133 == _T_15 ? _ram_T_129[287:0] : _GEN_3985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5036 = 10'h134 == _T_15 ? _ram_T_129[287:0] : _GEN_3986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5037 = 10'h135 == _T_15 ? _ram_T_129[287:0] : _GEN_3987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5038 = 10'h136 == _T_15 ? _ram_T_129[287:0] : _GEN_3988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5039 = 10'h137 == _T_15 ? _ram_T_129[287:0] : _GEN_3989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5040 = 10'h138 == _T_15 ? _ram_T_129[287:0] : _GEN_3990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5041 = 10'h139 == _T_15 ? _ram_T_129[287:0] : _GEN_3991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5042 = 10'h13a == _T_15 ? _ram_T_129[287:0] : _GEN_3992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5043 = 10'h13b == _T_15 ? _ram_T_129[287:0] : _GEN_3993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5044 = 10'h13c == _T_15 ? _ram_T_129[287:0] : _GEN_3994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5045 = 10'h13d == _T_15 ? _ram_T_129[287:0] : _GEN_3995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5046 = 10'h13e == _T_15 ? _ram_T_129[287:0] : _GEN_3996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5047 = 10'h13f == _T_15 ? _ram_T_129[287:0] : _GEN_3997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5048 = 10'h140 == _T_15 ? _ram_T_129[287:0] : _GEN_3998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5049 = 10'h141 == _T_15 ? _ram_T_129[287:0] : _GEN_3999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5050 = 10'h142 == _T_15 ? _ram_T_129[287:0] : _GEN_4000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5051 = 10'h143 == _T_15 ? _ram_T_129[287:0] : _GEN_4001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5052 = 10'h144 == _T_15 ? _ram_T_129[287:0] : _GEN_4002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5053 = 10'h145 == _T_15 ? _ram_T_129[287:0] : _GEN_4003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5054 = 10'h146 == _T_15 ? _ram_T_129[287:0] : _GEN_4004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5055 = 10'h147 == _T_15 ? _ram_T_129[287:0] : _GEN_4005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5056 = 10'h148 == _T_15 ? _ram_T_129[287:0] : _GEN_4006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5057 = 10'h149 == _T_15 ? _ram_T_129[287:0] : _GEN_4007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5058 = 10'h14a == _T_15 ? _ram_T_129[287:0] : _GEN_4008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5059 = 10'h14b == _T_15 ? _ram_T_129[287:0] : _GEN_4009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5060 = 10'h14c == _T_15 ? _ram_T_129[287:0] : _GEN_4010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5061 = 10'h14d == _T_15 ? _ram_T_129[287:0] : _GEN_4011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5062 = 10'h14e == _T_15 ? _ram_T_129[287:0] : _GEN_4012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5063 = 10'h14f == _T_15 ? _ram_T_129[287:0] : _GEN_4013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5064 = 10'h150 == _T_15 ? _ram_T_129[287:0] : _GEN_4014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5065 = 10'h151 == _T_15 ? _ram_T_129[287:0] : _GEN_4015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5066 = 10'h152 == _T_15 ? _ram_T_129[287:0] : _GEN_4016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5067 = 10'h153 == _T_15 ? _ram_T_129[287:0] : _GEN_4017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5068 = 10'h154 == _T_15 ? _ram_T_129[287:0] : _GEN_4018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5069 = 10'h155 == _T_15 ? _ram_T_129[287:0] : _GEN_4019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5070 = 10'h156 == _T_15 ? _ram_T_129[287:0] : _GEN_4020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5071 = 10'h157 == _T_15 ? _ram_T_129[287:0] : _GEN_4021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5072 = 10'h158 == _T_15 ? _ram_T_129[287:0] : _GEN_4022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5073 = 10'h159 == _T_15 ? _ram_T_129[287:0] : _GEN_4023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5074 = 10'h15a == _T_15 ? _ram_T_129[287:0] : _GEN_4024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5075 = 10'h15b == _T_15 ? _ram_T_129[287:0] : _GEN_4025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5076 = 10'h15c == _T_15 ? _ram_T_129[287:0] : _GEN_4026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5077 = 10'h15d == _T_15 ? _ram_T_129[287:0] : _GEN_4027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5078 = 10'h15e == _T_15 ? _ram_T_129[287:0] : _GEN_4028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5079 = 10'h15f == _T_15 ? _ram_T_129[287:0] : _GEN_4029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5080 = 10'h160 == _T_15 ? _ram_T_129[287:0] : _GEN_4030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5081 = 10'h161 == _T_15 ? _ram_T_129[287:0] : _GEN_4031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5082 = 10'h162 == _T_15 ? _ram_T_129[287:0] : _GEN_4032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5083 = 10'h163 == _T_15 ? _ram_T_129[287:0] : _GEN_4033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5084 = 10'h164 == _T_15 ? _ram_T_129[287:0] : _GEN_4034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5085 = 10'h165 == _T_15 ? _ram_T_129[287:0] : _GEN_4035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5086 = 10'h166 == _T_15 ? _ram_T_129[287:0] : _GEN_4036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5087 = 10'h167 == _T_15 ? _ram_T_129[287:0] : _GEN_4037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5088 = 10'h168 == _T_15 ? _ram_T_129[287:0] : _GEN_4038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5089 = 10'h169 == _T_15 ? _ram_T_129[287:0] : _GEN_4039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5090 = 10'h16a == _T_15 ? _ram_T_129[287:0] : _GEN_4040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5091 = 10'h16b == _T_15 ? _ram_T_129[287:0] : _GEN_4041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5092 = 10'h16c == _T_15 ? _ram_T_129[287:0] : _GEN_4042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5093 = 10'h16d == _T_15 ? _ram_T_129[287:0] : _GEN_4043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5094 = 10'h16e == _T_15 ? _ram_T_129[287:0] : _GEN_4044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5095 = 10'h16f == _T_15 ? _ram_T_129[287:0] : _GEN_4045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5096 = 10'h170 == _T_15 ? _ram_T_129[287:0] : _GEN_4046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5097 = 10'h171 == _T_15 ? _ram_T_129[287:0] : _GEN_4047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5098 = 10'h172 == _T_15 ? _ram_T_129[287:0] : _GEN_4048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5099 = 10'h173 == _T_15 ? _ram_T_129[287:0] : _GEN_4049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5100 = 10'h174 == _T_15 ? _ram_T_129[287:0] : _GEN_4050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5101 = 10'h175 == _T_15 ? _ram_T_129[287:0] : _GEN_4051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5102 = 10'h176 == _T_15 ? _ram_T_129[287:0] : _GEN_4052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5103 = 10'h177 == _T_15 ? _ram_T_129[287:0] : _GEN_4053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5104 = 10'h178 == _T_15 ? _ram_T_129[287:0] : _GEN_4054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5105 = 10'h179 == _T_15 ? _ram_T_129[287:0] : _GEN_4055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5106 = 10'h17a == _T_15 ? _ram_T_129[287:0] : _GEN_4056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5107 = 10'h17b == _T_15 ? _ram_T_129[287:0] : _GEN_4057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5108 = 10'h17c == _T_15 ? _ram_T_129[287:0] : _GEN_4058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5109 = 10'h17d == _T_15 ? _ram_T_129[287:0] : _GEN_4059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5110 = 10'h17e == _T_15 ? _ram_T_129[287:0] : _GEN_4060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5111 = 10'h17f == _T_15 ? _ram_T_129[287:0] : _GEN_4061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5112 = 10'h180 == _T_15 ? _ram_T_129[287:0] : _GEN_4062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5113 = 10'h181 == _T_15 ? _ram_T_129[287:0] : _GEN_4063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5114 = 10'h182 == _T_15 ? _ram_T_129[287:0] : _GEN_4064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5115 = 10'h183 == _T_15 ? _ram_T_129[287:0] : _GEN_4065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5116 = 10'h184 == _T_15 ? _ram_T_129[287:0] : _GEN_4066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5117 = 10'h185 == _T_15 ? _ram_T_129[287:0] : _GEN_4067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5118 = 10'h186 == _T_15 ? _ram_T_129[287:0] : _GEN_4068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5119 = 10'h187 == _T_15 ? _ram_T_129[287:0] : _GEN_4069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5120 = 10'h188 == _T_15 ? _ram_T_129[287:0] : _GEN_4070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5121 = 10'h189 == _T_15 ? _ram_T_129[287:0] : _GEN_4071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5122 = 10'h18a == _T_15 ? _ram_T_129[287:0] : _GEN_4072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5123 = 10'h18b == _T_15 ? _ram_T_129[287:0] : _GEN_4073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5124 = 10'h18c == _T_15 ? _ram_T_129[287:0] : _GEN_4074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5125 = 10'h18d == _T_15 ? _ram_T_129[287:0] : _GEN_4075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5126 = 10'h18e == _T_15 ? _ram_T_129[287:0] : _GEN_4076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5127 = 10'h18f == _T_15 ? _ram_T_129[287:0] : _GEN_4077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5128 = 10'h190 == _T_15 ? _ram_T_129[287:0] : _GEN_4078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5129 = 10'h191 == _T_15 ? _ram_T_129[287:0] : _GEN_4079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5130 = 10'h192 == _T_15 ? _ram_T_129[287:0] : _GEN_4080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5131 = 10'h193 == _T_15 ? _ram_T_129[287:0] : _GEN_4081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5132 = 10'h194 == _T_15 ? _ram_T_129[287:0] : _GEN_4082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5133 = 10'h195 == _T_15 ? _ram_T_129[287:0] : _GEN_4083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5134 = 10'h196 == _T_15 ? _ram_T_129[287:0] : _GEN_4084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5135 = 10'h197 == _T_15 ? _ram_T_129[287:0] : _GEN_4085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5136 = 10'h198 == _T_15 ? _ram_T_129[287:0] : _GEN_4086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5137 = 10'h199 == _T_15 ? _ram_T_129[287:0] : _GEN_4087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5138 = 10'h19a == _T_15 ? _ram_T_129[287:0] : _GEN_4088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5139 = 10'h19b == _T_15 ? _ram_T_129[287:0] : _GEN_4089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5140 = 10'h19c == _T_15 ? _ram_T_129[287:0] : _GEN_4090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5141 = 10'h19d == _T_15 ? _ram_T_129[287:0] : _GEN_4091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5142 = 10'h19e == _T_15 ? _ram_T_129[287:0] : _GEN_4092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5143 = 10'h19f == _T_15 ? _ram_T_129[287:0] : _GEN_4093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5144 = 10'h1a0 == _T_15 ? _ram_T_129[287:0] : _GEN_4094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5145 = 10'h1a1 == _T_15 ? _ram_T_129[287:0] : _GEN_4095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5146 = 10'h1a2 == _T_15 ? _ram_T_129[287:0] : _GEN_4096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5147 = 10'h1a3 == _T_15 ? _ram_T_129[287:0] : _GEN_4097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5148 = 10'h1a4 == _T_15 ? _ram_T_129[287:0] : _GEN_4098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5149 = 10'h1a5 == _T_15 ? _ram_T_129[287:0] : _GEN_4099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5150 = 10'h1a6 == _T_15 ? _ram_T_129[287:0] : _GEN_4100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5151 = 10'h1a7 == _T_15 ? _ram_T_129[287:0] : _GEN_4101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5152 = 10'h1a8 == _T_15 ? _ram_T_129[287:0] : _GEN_4102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5153 = 10'h1a9 == _T_15 ? _ram_T_129[287:0] : _GEN_4103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5154 = 10'h1aa == _T_15 ? _ram_T_129[287:0] : _GEN_4104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5155 = 10'h1ab == _T_15 ? _ram_T_129[287:0] : _GEN_4105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5156 = 10'h1ac == _T_15 ? _ram_T_129[287:0] : _GEN_4106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5157 = 10'h1ad == _T_15 ? _ram_T_129[287:0] : _GEN_4107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5158 = 10'h1ae == _T_15 ? _ram_T_129[287:0] : _GEN_4108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5159 = 10'h1af == _T_15 ? _ram_T_129[287:0] : _GEN_4109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5160 = 10'h1b0 == _T_15 ? _ram_T_129[287:0] : _GEN_4110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5161 = 10'h1b1 == _T_15 ? _ram_T_129[287:0] : _GEN_4111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5162 = 10'h1b2 == _T_15 ? _ram_T_129[287:0] : _GEN_4112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5163 = 10'h1b3 == _T_15 ? _ram_T_129[287:0] : _GEN_4113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5164 = 10'h1b4 == _T_15 ? _ram_T_129[287:0] : _GEN_4114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5165 = 10'h1b5 == _T_15 ? _ram_T_129[287:0] : _GEN_4115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5166 = 10'h1b6 == _T_15 ? _ram_T_129[287:0] : _GEN_4116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5167 = 10'h1b7 == _T_15 ? _ram_T_129[287:0] : _GEN_4117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5168 = 10'h1b8 == _T_15 ? _ram_T_129[287:0] : _GEN_4118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5169 = 10'h1b9 == _T_15 ? _ram_T_129[287:0] : _GEN_4119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5170 = 10'h1ba == _T_15 ? _ram_T_129[287:0] : _GEN_4120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5171 = 10'h1bb == _T_15 ? _ram_T_129[287:0] : _GEN_4121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5172 = 10'h1bc == _T_15 ? _ram_T_129[287:0] : _GEN_4122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5173 = 10'h1bd == _T_15 ? _ram_T_129[287:0] : _GEN_4123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5174 = 10'h1be == _T_15 ? _ram_T_129[287:0] : _GEN_4124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5175 = 10'h1bf == _T_15 ? _ram_T_129[287:0] : _GEN_4125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5176 = 10'h1c0 == _T_15 ? _ram_T_129[287:0] : _GEN_4126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5177 = 10'h1c1 == _T_15 ? _ram_T_129[287:0] : _GEN_4127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5178 = 10'h1c2 == _T_15 ? _ram_T_129[287:0] : _GEN_4128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5179 = 10'h1c3 == _T_15 ? _ram_T_129[287:0] : _GEN_4129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5180 = 10'h1c4 == _T_15 ? _ram_T_129[287:0] : _GEN_4130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5181 = 10'h1c5 == _T_15 ? _ram_T_129[287:0] : _GEN_4131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5182 = 10'h1c6 == _T_15 ? _ram_T_129[287:0] : _GEN_4132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5183 = 10'h1c7 == _T_15 ? _ram_T_129[287:0] : _GEN_4133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5184 = 10'h1c8 == _T_15 ? _ram_T_129[287:0] : _GEN_4134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5185 = 10'h1c9 == _T_15 ? _ram_T_129[287:0] : _GEN_4135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5186 = 10'h1ca == _T_15 ? _ram_T_129[287:0] : _GEN_4136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5187 = 10'h1cb == _T_15 ? _ram_T_129[287:0] : _GEN_4137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5188 = 10'h1cc == _T_15 ? _ram_T_129[287:0] : _GEN_4138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5189 = 10'h1cd == _T_15 ? _ram_T_129[287:0] : _GEN_4139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5190 = 10'h1ce == _T_15 ? _ram_T_129[287:0] : _GEN_4140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5191 = 10'h1cf == _T_15 ? _ram_T_129[287:0] : _GEN_4141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5192 = 10'h1d0 == _T_15 ? _ram_T_129[287:0] : _GEN_4142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5193 = 10'h1d1 == _T_15 ? _ram_T_129[287:0] : _GEN_4143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5194 = 10'h1d2 == _T_15 ? _ram_T_129[287:0] : _GEN_4144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5195 = 10'h1d3 == _T_15 ? _ram_T_129[287:0] : _GEN_4145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5196 = 10'h1d4 == _T_15 ? _ram_T_129[287:0] : _GEN_4146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5197 = 10'h1d5 == _T_15 ? _ram_T_129[287:0] : _GEN_4147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5198 = 10'h1d6 == _T_15 ? _ram_T_129[287:0] : _GEN_4148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5199 = 10'h1d7 == _T_15 ? _ram_T_129[287:0] : _GEN_4149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5200 = 10'h1d8 == _T_15 ? _ram_T_129[287:0] : _GEN_4150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5201 = 10'h1d9 == _T_15 ? _ram_T_129[287:0] : _GEN_4151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5202 = 10'h1da == _T_15 ? _ram_T_129[287:0] : _GEN_4152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5203 = 10'h1db == _T_15 ? _ram_T_129[287:0] : _GEN_4153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5204 = 10'h1dc == _T_15 ? _ram_T_129[287:0] : _GEN_4154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5205 = 10'h1dd == _T_15 ? _ram_T_129[287:0] : _GEN_4155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5206 = 10'h1de == _T_15 ? _ram_T_129[287:0] : _GEN_4156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5207 = 10'h1df == _T_15 ? _ram_T_129[287:0] : _GEN_4157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5208 = 10'h1e0 == _T_15 ? _ram_T_129[287:0] : _GEN_4158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5209 = 10'h1e1 == _T_15 ? _ram_T_129[287:0] : _GEN_4159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5210 = 10'h1e2 == _T_15 ? _ram_T_129[287:0] : _GEN_4160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5211 = 10'h1e3 == _T_15 ? _ram_T_129[287:0] : _GEN_4161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5212 = 10'h1e4 == _T_15 ? _ram_T_129[287:0] : _GEN_4162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5213 = 10'h1e5 == _T_15 ? _ram_T_129[287:0] : _GEN_4163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5214 = 10'h1e6 == _T_15 ? _ram_T_129[287:0] : _GEN_4164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5215 = 10'h1e7 == _T_15 ? _ram_T_129[287:0] : _GEN_4165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5216 = 10'h1e8 == _T_15 ? _ram_T_129[287:0] : _GEN_4166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5217 = 10'h1e9 == _T_15 ? _ram_T_129[287:0] : _GEN_4167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5218 = 10'h1ea == _T_15 ? _ram_T_129[287:0] : _GEN_4168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5219 = 10'h1eb == _T_15 ? _ram_T_129[287:0] : _GEN_4169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5220 = 10'h1ec == _T_15 ? _ram_T_129[287:0] : _GEN_4170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5221 = 10'h1ed == _T_15 ? _ram_T_129[287:0] : _GEN_4171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5222 = 10'h1ee == _T_15 ? _ram_T_129[287:0] : _GEN_4172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5223 = 10'h1ef == _T_15 ? _ram_T_129[287:0] : _GEN_4173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5224 = 10'h1f0 == _T_15 ? _ram_T_129[287:0] : _GEN_4174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5225 = 10'h1f1 == _T_15 ? _ram_T_129[287:0] : _GEN_4175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5226 = 10'h1f2 == _T_15 ? _ram_T_129[287:0] : _GEN_4176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5227 = 10'h1f3 == _T_15 ? _ram_T_129[287:0] : _GEN_4177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5228 = 10'h1f4 == _T_15 ? _ram_T_129[287:0] : _GEN_4178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5229 = 10'h1f5 == _T_15 ? _ram_T_129[287:0] : _GEN_4179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5230 = 10'h1f6 == _T_15 ? _ram_T_129[287:0] : _GEN_4180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5231 = 10'h1f7 == _T_15 ? _ram_T_129[287:0] : _GEN_4181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5232 = 10'h1f8 == _T_15 ? _ram_T_129[287:0] : _GEN_4182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5233 = 10'h1f9 == _T_15 ? _ram_T_129[287:0] : _GEN_4183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5234 = 10'h1fa == _T_15 ? _ram_T_129[287:0] : _GEN_4184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5235 = 10'h1fb == _T_15 ? _ram_T_129[287:0] : _GEN_4185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5236 = 10'h1fc == _T_15 ? _ram_T_129[287:0] : _GEN_4186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5237 = 10'h1fd == _T_15 ? _ram_T_129[287:0] : _GEN_4187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5238 = 10'h1fe == _T_15 ? _ram_T_129[287:0] : _GEN_4188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5239 = 10'h1ff == _T_15 ? _ram_T_129[287:0] : _GEN_4189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5240 = 10'h200 == _T_15 ? _ram_T_129[287:0] : _GEN_4190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5241 = 10'h201 == _T_15 ? _ram_T_129[287:0] : _GEN_4191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5242 = 10'h202 == _T_15 ? _ram_T_129[287:0] : _GEN_4192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5243 = 10'h203 == _T_15 ? _ram_T_129[287:0] : _GEN_4193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5244 = 10'h204 == _T_15 ? _ram_T_129[287:0] : _GEN_4194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5245 = 10'h205 == _T_15 ? _ram_T_129[287:0] : _GEN_4195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5246 = 10'h206 == _T_15 ? _ram_T_129[287:0] : _GEN_4196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5247 = 10'h207 == _T_15 ? _ram_T_129[287:0] : _GEN_4197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5248 = 10'h208 == _T_15 ? _ram_T_129[287:0] : _GEN_4198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5249 = 10'h209 == _T_15 ? _ram_T_129[287:0] : _GEN_4199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5250 = 10'h20a == _T_15 ? _ram_T_129[287:0] : _GEN_4200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5251 = 10'h20b == _T_15 ? _ram_T_129[287:0] : _GEN_4201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5252 = 10'h20c == _T_15 ? _ram_T_129[287:0] : _GEN_4202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_17 = h + 10'h5; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_5 = vga_mem_ram_MPORT_45_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_5 = vga_mem_ram_MPORT_46_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_5 = vga_mem_ram_MPORT_47_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_5 = vga_mem_ram_MPORT_48_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_5 = vga_mem_ram_MPORT_49_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_5 = vga_mem_ram_MPORT_50_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_5 = vga_mem_ram_MPORT_51_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_5 = vga_mem_ram_MPORT_52_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_5 = vga_mem_ram_MPORT_53_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_150 = {278'h0,ram_hi_hi_hi_lo_5,ram_hi_hi_lo_5,ram_hi_lo_hi_5,ram_hi_lo_lo_5,ram_lo_hi_hi_hi_5,
    ram_lo_hi_hi_lo_5,ram_lo_hi_lo_5,ram_lo_lo_hi_5,ram_lo_lo_lo_5}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19070 = {{8191'd0}, _ram_T_150}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_154 = _GEN_19070 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_5254 = 10'h1 == _T_17 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5255 = 10'h2 == _T_17 ? ram_2 : _GEN_5254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5256 = 10'h3 == _T_17 ? ram_3 : _GEN_5255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5257 = 10'h4 == _T_17 ? ram_4 : _GEN_5256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5258 = 10'h5 == _T_17 ? ram_5 : _GEN_5257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5259 = 10'h6 == _T_17 ? ram_6 : _GEN_5258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5260 = 10'h7 == _T_17 ? ram_7 : _GEN_5259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5261 = 10'h8 == _T_17 ? ram_8 : _GEN_5260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5262 = 10'h9 == _T_17 ? ram_9 : _GEN_5261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5263 = 10'ha == _T_17 ? ram_10 : _GEN_5262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5264 = 10'hb == _T_17 ? ram_11 : _GEN_5263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5265 = 10'hc == _T_17 ? ram_12 : _GEN_5264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5266 = 10'hd == _T_17 ? ram_13 : _GEN_5265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5267 = 10'he == _T_17 ? ram_14 : _GEN_5266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5268 = 10'hf == _T_17 ? ram_15 : _GEN_5267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5269 = 10'h10 == _T_17 ? ram_16 : _GEN_5268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5270 = 10'h11 == _T_17 ? ram_17 : _GEN_5269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5271 = 10'h12 == _T_17 ? ram_18 : _GEN_5270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5272 = 10'h13 == _T_17 ? ram_19 : _GEN_5271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5273 = 10'h14 == _T_17 ? ram_20 : _GEN_5272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5274 = 10'h15 == _T_17 ? ram_21 : _GEN_5273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5275 = 10'h16 == _T_17 ? ram_22 : _GEN_5274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5276 = 10'h17 == _T_17 ? ram_23 : _GEN_5275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5277 = 10'h18 == _T_17 ? ram_24 : _GEN_5276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5278 = 10'h19 == _T_17 ? ram_25 : _GEN_5277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5279 = 10'h1a == _T_17 ? ram_26 : _GEN_5278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5280 = 10'h1b == _T_17 ? ram_27 : _GEN_5279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5281 = 10'h1c == _T_17 ? ram_28 : _GEN_5280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5282 = 10'h1d == _T_17 ? ram_29 : _GEN_5281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5283 = 10'h1e == _T_17 ? ram_30 : _GEN_5282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5284 = 10'h1f == _T_17 ? ram_31 : _GEN_5283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5285 = 10'h20 == _T_17 ? ram_32 : _GEN_5284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5286 = 10'h21 == _T_17 ? ram_33 : _GEN_5285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5287 = 10'h22 == _T_17 ? ram_34 : _GEN_5286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5288 = 10'h23 == _T_17 ? ram_35 : _GEN_5287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5289 = 10'h24 == _T_17 ? ram_36 : _GEN_5288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5290 = 10'h25 == _T_17 ? ram_37 : _GEN_5289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5291 = 10'h26 == _T_17 ? ram_38 : _GEN_5290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5292 = 10'h27 == _T_17 ? ram_39 : _GEN_5291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5293 = 10'h28 == _T_17 ? ram_40 : _GEN_5292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5294 = 10'h29 == _T_17 ? ram_41 : _GEN_5293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5295 = 10'h2a == _T_17 ? ram_42 : _GEN_5294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5296 = 10'h2b == _T_17 ? ram_43 : _GEN_5295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5297 = 10'h2c == _T_17 ? ram_44 : _GEN_5296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5298 = 10'h2d == _T_17 ? ram_45 : _GEN_5297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5299 = 10'h2e == _T_17 ? ram_46 : _GEN_5298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5300 = 10'h2f == _T_17 ? ram_47 : _GEN_5299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5301 = 10'h30 == _T_17 ? ram_48 : _GEN_5300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5302 = 10'h31 == _T_17 ? ram_49 : _GEN_5301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5303 = 10'h32 == _T_17 ? ram_50 : _GEN_5302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5304 = 10'h33 == _T_17 ? ram_51 : _GEN_5303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5305 = 10'h34 == _T_17 ? ram_52 : _GEN_5304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5306 = 10'h35 == _T_17 ? ram_53 : _GEN_5305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5307 = 10'h36 == _T_17 ? ram_54 : _GEN_5306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5308 = 10'h37 == _T_17 ? ram_55 : _GEN_5307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5309 = 10'h38 == _T_17 ? ram_56 : _GEN_5308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5310 = 10'h39 == _T_17 ? ram_57 : _GEN_5309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5311 = 10'h3a == _T_17 ? ram_58 : _GEN_5310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5312 = 10'h3b == _T_17 ? ram_59 : _GEN_5311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5313 = 10'h3c == _T_17 ? ram_60 : _GEN_5312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5314 = 10'h3d == _T_17 ? ram_61 : _GEN_5313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5315 = 10'h3e == _T_17 ? ram_62 : _GEN_5314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5316 = 10'h3f == _T_17 ? ram_63 : _GEN_5315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5317 = 10'h40 == _T_17 ? ram_64 : _GEN_5316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5318 = 10'h41 == _T_17 ? ram_65 : _GEN_5317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5319 = 10'h42 == _T_17 ? ram_66 : _GEN_5318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5320 = 10'h43 == _T_17 ? ram_67 : _GEN_5319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5321 = 10'h44 == _T_17 ? ram_68 : _GEN_5320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5322 = 10'h45 == _T_17 ? ram_69 : _GEN_5321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5323 = 10'h46 == _T_17 ? ram_70 : _GEN_5322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5324 = 10'h47 == _T_17 ? ram_71 : _GEN_5323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5325 = 10'h48 == _T_17 ? ram_72 : _GEN_5324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5326 = 10'h49 == _T_17 ? ram_73 : _GEN_5325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5327 = 10'h4a == _T_17 ? ram_74 : _GEN_5326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5328 = 10'h4b == _T_17 ? ram_75 : _GEN_5327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5329 = 10'h4c == _T_17 ? ram_76 : _GEN_5328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5330 = 10'h4d == _T_17 ? ram_77 : _GEN_5329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5331 = 10'h4e == _T_17 ? ram_78 : _GEN_5330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5332 = 10'h4f == _T_17 ? ram_79 : _GEN_5331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5333 = 10'h50 == _T_17 ? ram_80 : _GEN_5332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5334 = 10'h51 == _T_17 ? ram_81 : _GEN_5333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5335 = 10'h52 == _T_17 ? ram_82 : _GEN_5334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5336 = 10'h53 == _T_17 ? ram_83 : _GEN_5335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5337 = 10'h54 == _T_17 ? ram_84 : _GEN_5336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5338 = 10'h55 == _T_17 ? ram_85 : _GEN_5337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5339 = 10'h56 == _T_17 ? ram_86 : _GEN_5338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5340 = 10'h57 == _T_17 ? ram_87 : _GEN_5339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5341 = 10'h58 == _T_17 ? ram_88 : _GEN_5340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5342 = 10'h59 == _T_17 ? ram_89 : _GEN_5341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5343 = 10'h5a == _T_17 ? ram_90 : _GEN_5342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5344 = 10'h5b == _T_17 ? ram_91 : _GEN_5343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5345 = 10'h5c == _T_17 ? ram_92 : _GEN_5344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5346 = 10'h5d == _T_17 ? ram_93 : _GEN_5345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5347 = 10'h5e == _T_17 ? ram_94 : _GEN_5346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5348 = 10'h5f == _T_17 ? ram_95 : _GEN_5347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5349 = 10'h60 == _T_17 ? ram_96 : _GEN_5348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5350 = 10'h61 == _T_17 ? ram_97 : _GEN_5349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5351 = 10'h62 == _T_17 ? ram_98 : _GEN_5350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5352 = 10'h63 == _T_17 ? ram_99 : _GEN_5351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5353 = 10'h64 == _T_17 ? ram_100 : _GEN_5352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5354 = 10'h65 == _T_17 ? ram_101 : _GEN_5353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5355 = 10'h66 == _T_17 ? ram_102 : _GEN_5354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5356 = 10'h67 == _T_17 ? ram_103 : _GEN_5355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5357 = 10'h68 == _T_17 ? ram_104 : _GEN_5356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5358 = 10'h69 == _T_17 ? ram_105 : _GEN_5357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5359 = 10'h6a == _T_17 ? ram_106 : _GEN_5358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5360 = 10'h6b == _T_17 ? ram_107 : _GEN_5359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5361 = 10'h6c == _T_17 ? ram_108 : _GEN_5360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5362 = 10'h6d == _T_17 ? ram_109 : _GEN_5361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5363 = 10'h6e == _T_17 ? ram_110 : _GEN_5362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5364 = 10'h6f == _T_17 ? ram_111 : _GEN_5363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5365 = 10'h70 == _T_17 ? ram_112 : _GEN_5364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5366 = 10'h71 == _T_17 ? ram_113 : _GEN_5365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5367 = 10'h72 == _T_17 ? ram_114 : _GEN_5366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5368 = 10'h73 == _T_17 ? ram_115 : _GEN_5367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5369 = 10'h74 == _T_17 ? ram_116 : _GEN_5368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5370 = 10'h75 == _T_17 ? ram_117 : _GEN_5369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5371 = 10'h76 == _T_17 ? ram_118 : _GEN_5370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5372 = 10'h77 == _T_17 ? ram_119 : _GEN_5371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5373 = 10'h78 == _T_17 ? ram_120 : _GEN_5372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5374 = 10'h79 == _T_17 ? ram_121 : _GEN_5373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5375 = 10'h7a == _T_17 ? ram_122 : _GEN_5374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5376 = 10'h7b == _T_17 ? ram_123 : _GEN_5375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5377 = 10'h7c == _T_17 ? ram_124 : _GEN_5376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5378 = 10'h7d == _T_17 ? ram_125 : _GEN_5377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5379 = 10'h7e == _T_17 ? ram_126 : _GEN_5378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5380 = 10'h7f == _T_17 ? ram_127 : _GEN_5379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5381 = 10'h80 == _T_17 ? ram_128 : _GEN_5380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5382 = 10'h81 == _T_17 ? ram_129 : _GEN_5381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5383 = 10'h82 == _T_17 ? ram_130 : _GEN_5382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5384 = 10'h83 == _T_17 ? ram_131 : _GEN_5383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5385 = 10'h84 == _T_17 ? ram_132 : _GEN_5384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5386 = 10'h85 == _T_17 ? ram_133 : _GEN_5385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5387 = 10'h86 == _T_17 ? ram_134 : _GEN_5386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5388 = 10'h87 == _T_17 ? ram_135 : _GEN_5387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5389 = 10'h88 == _T_17 ? ram_136 : _GEN_5388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5390 = 10'h89 == _T_17 ? ram_137 : _GEN_5389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5391 = 10'h8a == _T_17 ? ram_138 : _GEN_5390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5392 = 10'h8b == _T_17 ? ram_139 : _GEN_5391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5393 = 10'h8c == _T_17 ? ram_140 : _GEN_5392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5394 = 10'h8d == _T_17 ? ram_141 : _GEN_5393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5395 = 10'h8e == _T_17 ? ram_142 : _GEN_5394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5396 = 10'h8f == _T_17 ? ram_143 : _GEN_5395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5397 = 10'h90 == _T_17 ? ram_144 : _GEN_5396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5398 = 10'h91 == _T_17 ? ram_145 : _GEN_5397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5399 = 10'h92 == _T_17 ? ram_146 : _GEN_5398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5400 = 10'h93 == _T_17 ? ram_147 : _GEN_5399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5401 = 10'h94 == _T_17 ? ram_148 : _GEN_5400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5402 = 10'h95 == _T_17 ? ram_149 : _GEN_5401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5403 = 10'h96 == _T_17 ? ram_150 : _GEN_5402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5404 = 10'h97 == _T_17 ? ram_151 : _GEN_5403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5405 = 10'h98 == _T_17 ? ram_152 : _GEN_5404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5406 = 10'h99 == _T_17 ? ram_153 : _GEN_5405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5407 = 10'h9a == _T_17 ? ram_154 : _GEN_5406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5408 = 10'h9b == _T_17 ? ram_155 : _GEN_5407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5409 = 10'h9c == _T_17 ? ram_156 : _GEN_5408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5410 = 10'h9d == _T_17 ? ram_157 : _GEN_5409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5411 = 10'h9e == _T_17 ? ram_158 : _GEN_5410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5412 = 10'h9f == _T_17 ? ram_159 : _GEN_5411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5413 = 10'ha0 == _T_17 ? ram_160 : _GEN_5412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5414 = 10'ha1 == _T_17 ? ram_161 : _GEN_5413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5415 = 10'ha2 == _T_17 ? ram_162 : _GEN_5414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5416 = 10'ha3 == _T_17 ? ram_163 : _GEN_5415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5417 = 10'ha4 == _T_17 ? ram_164 : _GEN_5416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5418 = 10'ha5 == _T_17 ? ram_165 : _GEN_5417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5419 = 10'ha6 == _T_17 ? ram_166 : _GEN_5418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5420 = 10'ha7 == _T_17 ? ram_167 : _GEN_5419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5421 = 10'ha8 == _T_17 ? ram_168 : _GEN_5420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5422 = 10'ha9 == _T_17 ? ram_169 : _GEN_5421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5423 = 10'haa == _T_17 ? ram_170 : _GEN_5422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5424 = 10'hab == _T_17 ? ram_171 : _GEN_5423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5425 = 10'hac == _T_17 ? ram_172 : _GEN_5424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5426 = 10'had == _T_17 ? ram_173 : _GEN_5425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5427 = 10'hae == _T_17 ? ram_174 : _GEN_5426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5428 = 10'haf == _T_17 ? ram_175 : _GEN_5427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5429 = 10'hb0 == _T_17 ? ram_176 : _GEN_5428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5430 = 10'hb1 == _T_17 ? ram_177 : _GEN_5429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5431 = 10'hb2 == _T_17 ? ram_178 : _GEN_5430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5432 = 10'hb3 == _T_17 ? ram_179 : _GEN_5431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5433 = 10'hb4 == _T_17 ? ram_180 : _GEN_5432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5434 = 10'hb5 == _T_17 ? ram_181 : _GEN_5433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5435 = 10'hb6 == _T_17 ? ram_182 : _GEN_5434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5436 = 10'hb7 == _T_17 ? ram_183 : _GEN_5435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5437 = 10'hb8 == _T_17 ? ram_184 : _GEN_5436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5438 = 10'hb9 == _T_17 ? ram_185 : _GEN_5437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5439 = 10'hba == _T_17 ? ram_186 : _GEN_5438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5440 = 10'hbb == _T_17 ? ram_187 : _GEN_5439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5441 = 10'hbc == _T_17 ? ram_188 : _GEN_5440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5442 = 10'hbd == _T_17 ? ram_189 : _GEN_5441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5443 = 10'hbe == _T_17 ? ram_190 : _GEN_5442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5444 = 10'hbf == _T_17 ? ram_191 : _GEN_5443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5445 = 10'hc0 == _T_17 ? ram_192 : _GEN_5444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5446 = 10'hc1 == _T_17 ? ram_193 : _GEN_5445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5447 = 10'hc2 == _T_17 ? ram_194 : _GEN_5446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5448 = 10'hc3 == _T_17 ? ram_195 : _GEN_5447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5449 = 10'hc4 == _T_17 ? ram_196 : _GEN_5448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5450 = 10'hc5 == _T_17 ? ram_197 : _GEN_5449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5451 = 10'hc6 == _T_17 ? ram_198 : _GEN_5450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5452 = 10'hc7 == _T_17 ? ram_199 : _GEN_5451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5453 = 10'hc8 == _T_17 ? ram_200 : _GEN_5452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5454 = 10'hc9 == _T_17 ? ram_201 : _GEN_5453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5455 = 10'hca == _T_17 ? ram_202 : _GEN_5454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5456 = 10'hcb == _T_17 ? ram_203 : _GEN_5455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5457 = 10'hcc == _T_17 ? ram_204 : _GEN_5456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5458 = 10'hcd == _T_17 ? ram_205 : _GEN_5457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5459 = 10'hce == _T_17 ? ram_206 : _GEN_5458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5460 = 10'hcf == _T_17 ? ram_207 : _GEN_5459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5461 = 10'hd0 == _T_17 ? ram_208 : _GEN_5460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5462 = 10'hd1 == _T_17 ? ram_209 : _GEN_5461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5463 = 10'hd2 == _T_17 ? ram_210 : _GEN_5462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5464 = 10'hd3 == _T_17 ? ram_211 : _GEN_5463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5465 = 10'hd4 == _T_17 ? ram_212 : _GEN_5464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5466 = 10'hd5 == _T_17 ? ram_213 : _GEN_5465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5467 = 10'hd6 == _T_17 ? ram_214 : _GEN_5466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5468 = 10'hd7 == _T_17 ? ram_215 : _GEN_5467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5469 = 10'hd8 == _T_17 ? ram_216 : _GEN_5468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5470 = 10'hd9 == _T_17 ? ram_217 : _GEN_5469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5471 = 10'hda == _T_17 ? ram_218 : _GEN_5470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5472 = 10'hdb == _T_17 ? ram_219 : _GEN_5471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5473 = 10'hdc == _T_17 ? ram_220 : _GEN_5472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5474 = 10'hdd == _T_17 ? ram_221 : _GEN_5473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5475 = 10'hde == _T_17 ? ram_222 : _GEN_5474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5476 = 10'hdf == _T_17 ? ram_223 : _GEN_5475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5477 = 10'he0 == _T_17 ? ram_224 : _GEN_5476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5478 = 10'he1 == _T_17 ? ram_225 : _GEN_5477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5479 = 10'he2 == _T_17 ? ram_226 : _GEN_5478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5480 = 10'he3 == _T_17 ? ram_227 : _GEN_5479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5481 = 10'he4 == _T_17 ? ram_228 : _GEN_5480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5482 = 10'he5 == _T_17 ? ram_229 : _GEN_5481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5483 = 10'he6 == _T_17 ? ram_230 : _GEN_5482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5484 = 10'he7 == _T_17 ? ram_231 : _GEN_5483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5485 = 10'he8 == _T_17 ? ram_232 : _GEN_5484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5486 = 10'he9 == _T_17 ? ram_233 : _GEN_5485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5487 = 10'hea == _T_17 ? ram_234 : _GEN_5486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5488 = 10'heb == _T_17 ? ram_235 : _GEN_5487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5489 = 10'hec == _T_17 ? ram_236 : _GEN_5488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5490 = 10'hed == _T_17 ? ram_237 : _GEN_5489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5491 = 10'hee == _T_17 ? ram_238 : _GEN_5490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5492 = 10'hef == _T_17 ? ram_239 : _GEN_5491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5493 = 10'hf0 == _T_17 ? ram_240 : _GEN_5492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5494 = 10'hf1 == _T_17 ? ram_241 : _GEN_5493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5495 = 10'hf2 == _T_17 ? ram_242 : _GEN_5494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5496 = 10'hf3 == _T_17 ? ram_243 : _GEN_5495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5497 = 10'hf4 == _T_17 ? ram_244 : _GEN_5496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5498 = 10'hf5 == _T_17 ? ram_245 : _GEN_5497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5499 = 10'hf6 == _T_17 ? ram_246 : _GEN_5498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5500 = 10'hf7 == _T_17 ? ram_247 : _GEN_5499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5501 = 10'hf8 == _T_17 ? ram_248 : _GEN_5500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5502 = 10'hf9 == _T_17 ? ram_249 : _GEN_5501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5503 = 10'hfa == _T_17 ? ram_250 : _GEN_5502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5504 = 10'hfb == _T_17 ? ram_251 : _GEN_5503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5505 = 10'hfc == _T_17 ? ram_252 : _GEN_5504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5506 = 10'hfd == _T_17 ? ram_253 : _GEN_5505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5507 = 10'hfe == _T_17 ? ram_254 : _GEN_5506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5508 = 10'hff == _T_17 ? ram_255 : _GEN_5507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5509 = 10'h100 == _T_17 ? ram_256 : _GEN_5508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5510 = 10'h101 == _T_17 ? ram_257 : _GEN_5509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5511 = 10'h102 == _T_17 ? ram_258 : _GEN_5510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5512 = 10'h103 == _T_17 ? ram_259 : _GEN_5511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5513 = 10'h104 == _T_17 ? ram_260 : _GEN_5512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5514 = 10'h105 == _T_17 ? ram_261 : _GEN_5513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5515 = 10'h106 == _T_17 ? ram_262 : _GEN_5514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5516 = 10'h107 == _T_17 ? ram_263 : _GEN_5515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5517 = 10'h108 == _T_17 ? ram_264 : _GEN_5516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5518 = 10'h109 == _T_17 ? ram_265 : _GEN_5517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5519 = 10'h10a == _T_17 ? ram_266 : _GEN_5518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5520 = 10'h10b == _T_17 ? ram_267 : _GEN_5519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5521 = 10'h10c == _T_17 ? ram_268 : _GEN_5520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5522 = 10'h10d == _T_17 ? ram_269 : _GEN_5521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5523 = 10'h10e == _T_17 ? ram_270 : _GEN_5522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5524 = 10'h10f == _T_17 ? ram_271 : _GEN_5523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5525 = 10'h110 == _T_17 ? ram_272 : _GEN_5524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5526 = 10'h111 == _T_17 ? ram_273 : _GEN_5525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5527 = 10'h112 == _T_17 ? ram_274 : _GEN_5526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5528 = 10'h113 == _T_17 ? ram_275 : _GEN_5527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5529 = 10'h114 == _T_17 ? ram_276 : _GEN_5528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5530 = 10'h115 == _T_17 ? ram_277 : _GEN_5529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5531 = 10'h116 == _T_17 ? ram_278 : _GEN_5530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5532 = 10'h117 == _T_17 ? ram_279 : _GEN_5531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5533 = 10'h118 == _T_17 ? ram_280 : _GEN_5532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5534 = 10'h119 == _T_17 ? ram_281 : _GEN_5533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5535 = 10'h11a == _T_17 ? ram_282 : _GEN_5534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5536 = 10'h11b == _T_17 ? ram_283 : _GEN_5535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5537 = 10'h11c == _T_17 ? ram_284 : _GEN_5536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5538 = 10'h11d == _T_17 ? ram_285 : _GEN_5537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5539 = 10'h11e == _T_17 ? ram_286 : _GEN_5538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5540 = 10'h11f == _T_17 ? ram_287 : _GEN_5539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5541 = 10'h120 == _T_17 ? ram_288 : _GEN_5540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5542 = 10'h121 == _T_17 ? ram_289 : _GEN_5541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5543 = 10'h122 == _T_17 ? ram_290 : _GEN_5542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5544 = 10'h123 == _T_17 ? ram_291 : _GEN_5543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5545 = 10'h124 == _T_17 ? ram_292 : _GEN_5544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5546 = 10'h125 == _T_17 ? ram_293 : _GEN_5545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5547 = 10'h126 == _T_17 ? ram_294 : _GEN_5546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5548 = 10'h127 == _T_17 ? ram_295 : _GEN_5547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5549 = 10'h128 == _T_17 ? ram_296 : _GEN_5548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5550 = 10'h129 == _T_17 ? ram_297 : _GEN_5549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5551 = 10'h12a == _T_17 ? ram_298 : _GEN_5550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5552 = 10'h12b == _T_17 ? ram_299 : _GEN_5551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5553 = 10'h12c == _T_17 ? ram_300 : _GEN_5552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5554 = 10'h12d == _T_17 ? ram_301 : _GEN_5553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5555 = 10'h12e == _T_17 ? ram_302 : _GEN_5554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5556 = 10'h12f == _T_17 ? ram_303 : _GEN_5555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5557 = 10'h130 == _T_17 ? ram_304 : _GEN_5556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5558 = 10'h131 == _T_17 ? ram_305 : _GEN_5557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5559 = 10'h132 == _T_17 ? ram_306 : _GEN_5558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5560 = 10'h133 == _T_17 ? ram_307 : _GEN_5559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5561 = 10'h134 == _T_17 ? ram_308 : _GEN_5560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5562 = 10'h135 == _T_17 ? ram_309 : _GEN_5561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5563 = 10'h136 == _T_17 ? ram_310 : _GEN_5562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5564 = 10'h137 == _T_17 ? ram_311 : _GEN_5563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5565 = 10'h138 == _T_17 ? ram_312 : _GEN_5564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5566 = 10'h139 == _T_17 ? ram_313 : _GEN_5565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5567 = 10'h13a == _T_17 ? ram_314 : _GEN_5566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5568 = 10'h13b == _T_17 ? ram_315 : _GEN_5567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5569 = 10'h13c == _T_17 ? ram_316 : _GEN_5568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5570 = 10'h13d == _T_17 ? ram_317 : _GEN_5569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5571 = 10'h13e == _T_17 ? ram_318 : _GEN_5570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5572 = 10'h13f == _T_17 ? ram_319 : _GEN_5571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5573 = 10'h140 == _T_17 ? ram_320 : _GEN_5572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5574 = 10'h141 == _T_17 ? ram_321 : _GEN_5573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5575 = 10'h142 == _T_17 ? ram_322 : _GEN_5574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5576 = 10'h143 == _T_17 ? ram_323 : _GEN_5575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5577 = 10'h144 == _T_17 ? ram_324 : _GEN_5576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5578 = 10'h145 == _T_17 ? ram_325 : _GEN_5577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5579 = 10'h146 == _T_17 ? ram_326 : _GEN_5578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5580 = 10'h147 == _T_17 ? ram_327 : _GEN_5579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5581 = 10'h148 == _T_17 ? ram_328 : _GEN_5580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5582 = 10'h149 == _T_17 ? ram_329 : _GEN_5581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5583 = 10'h14a == _T_17 ? ram_330 : _GEN_5582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5584 = 10'h14b == _T_17 ? ram_331 : _GEN_5583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5585 = 10'h14c == _T_17 ? ram_332 : _GEN_5584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5586 = 10'h14d == _T_17 ? ram_333 : _GEN_5585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5587 = 10'h14e == _T_17 ? ram_334 : _GEN_5586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5588 = 10'h14f == _T_17 ? ram_335 : _GEN_5587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5589 = 10'h150 == _T_17 ? ram_336 : _GEN_5588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5590 = 10'h151 == _T_17 ? ram_337 : _GEN_5589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5591 = 10'h152 == _T_17 ? ram_338 : _GEN_5590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5592 = 10'h153 == _T_17 ? ram_339 : _GEN_5591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5593 = 10'h154 == _T_17 ? ram_340 : _GEN_5592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5594 = 10'h155 == _T_17 ? ram_341 : _GEN_5593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5595 = 10'h156 == _T_17 ? ram_342 : _GEN_5594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5596 = 10'h157 == _T_17 ? ram_343 : _GEN_5595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5597 = 10'h158 == _T_17 ? ram_344 : _GEN_5596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5598 = 10'h159 == _T_17 ? ram_345 : _GEN_5597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5599 = 10'h15a == _T_17 ? ram_346 : _GEN_5598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5600 = 10'h15b == _T_17 ? ram_347 : _GEN_5599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5601 = 10'h15c == _T_17 ? ram_348 : _GEN_5600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5602 = 10'h15d == _T_17 ? ram_349 : _GEN_5601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5603 = 10'h15e == _T_17 ? ram_350 : _GEN_5602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5604 = 10'h15f == _T_17 ? ram_351 : _GEN_5603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5605 = 10'h160 == _T_17 ? ram_352 : _GEN_5604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5606 = 10'h161 == _T_17 ? ram_353 : _GEN_5605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5607 = 10'h162 == _T_17 ? ram_354 : _GEN_5606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5608 = 10'h163 == _T_17 ? ram_355 : _GEN_5607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5609 = 10'h164 == _T_17 ? ram_356 : _GEN_5608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5610 = 10'h165 == _T_17 ? ram_357 : _GEN_5609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5611 = 10'h166 == _T_17 ? ram_358 : _GEN_5610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5612 = 10'h167 == _T_17 ? ram_359 : _GEN_5611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5613 = 10'h168 == _T_17 ? ram_360 : _GEN_5612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5614 = 10'h169 == _T_17 ? ram_361 : _GEN_5613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5615 = 10'h16a == _T_17 ? ram_362 : _GEN_5614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5616 = 10'h16b == _T_17 ? ram_363 : _GEN_5615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5617 = 10'h16c == _T_17 ? ram_364 : _GEN_5616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5618 = 10'h16d == _T_17 ? ram_365 : _GEN_5617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5619 = 10'h16e == _T_17 ? ram_366 : _GEN_5618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5620 = 10'h16f == _T_17 ? ram_367 : _GEN_5619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5621 = 10'h170 == _T_17 ? ram_368 : _GEN_5620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5622 = 10'h171 == _T_17 ? ram_369 : _GEN_5621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5623 = 10'h172 == _T_17 ? ram_370 : _GEN_5622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5624 = 10'h173 == _T_17 ? ram_371 : _GEN_5623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5625 = 10'h174 == _T_17 ? ram_372 : _GEN_5624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5626 = 10'h175 == _T_17 ? ram_373 : _GEN_5625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5627 = 10'h176 == _T_17 ? ram_374 : _GEN_5626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5628 = 10'h177 == _T_17 ? ram_375 : _GEN_5627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5629 = 10'h178 == _T_17 ? ram_376 : _GEN_5628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5630 = 10'h179 == _T_17 ? ram_377 : _GEN_5629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5631 = 10'h17a == _T_17 ? ram_378 : _GEN_5630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5632 = 10'h17b == _T_17 ? ram_379 : _GEN_5631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5633 = 10'h17c == _T_17 ? ram_380 : _GEN_5632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5634 = 10'h17d == _T_17 ? ram_381 : _GEN_5633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5635 = 10'h17e == _T_17 ? ram_382 : _GEN_5634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5636 = 10'h17f == _T_17 ? ram_383 : _GEN_5635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5637 = 10'h180 == _T_17 ? ram_384 : _GEN_5636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5638 = 10'h181 == _T_17 ? ram_385 : _GEN_5637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5639 = 10'h182 == _T_17 ? ram_386 : _GEN_5638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5640 = 10'h183 == _T_17 ? ram_387 : _GEN_5639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5641 = 10'h184 == _T_17 ? ram_388 : _GEN_5640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5642 = 10'h185 == _T_17 ? ram_389 : _GEN_5641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5643 = 10'h186 == _T_17 ? ram_390 : _GEN_5642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5644 = 10'h187 == _T_17 ? ram_391 : _GEN_5643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5645 = 10'h188 == _T_17 ? ram_392 : _GEN_5644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5646 = 10'h189 == _T_17 ? ram_393 : _GEN_5645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5647 = 10'h18a == _T_17 ? ram_394 : _GEN_5646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5648 = 10'h18b == _T_17 ? ram_395 : _GEN_5647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5649 = 10'h18c == _T_17 ? ram_396 : _GEN_5648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5650 = 10'h18d == _T_17 ? ram_397 : _GEN_5649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5651 = 10'h18e == _T_17 ? ram_398 : _GEN_5650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5652 = 10'h18f == _T_17 ? ram_399 : _GEN_5651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5653 = 10'h190 == _T_17 ? ram_400 : _GEN_5652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5654 = 10'h191 == _T_17 ? ram_401 : _GEN_5653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5655 = 10'h192 == _T_17 ? ram_402 : _GEN_5654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5656 = 10'h193 == _T_17 ? ram_403 : _GEN_5655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5657 = 10'h194 == _T_17 ? ram_404 : _GEN_5656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5658 = 10'h195 == _T_17 ? ram_405 : _GEN_5657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5659 = 10'h196 == _T_17 ? ram_406 : _GEN_5658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5660 = 10'h197 == _T_17 ? ram_407 : _GEN_5659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5661 = 10'h198 == _T_17 ? ram_408 : _GEN_5660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5662 = 10'h199 == _T_17 ? ram_409 : _GEN_5661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5663 = 10'h19a == _T_17 ? ram_410 : _GEN_5662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5664 = 10'h19b == _T_17 ? ram_411 : _GEN_5663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5665 = 10'h19c == _T_17 ? ram_412 : _GEN_5664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5666 = 10'h19d == _T_17 ? ram_413 : _GEN_5665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5667 = 10'h19e == _T_17 ? ram_414 : _GEN_5666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5668 = 10'h19f == _T_17 ? ram_415 : _GEN_5667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5669 = 10'h1a0 == _T_17 ? ram_416 : _GEN_5668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5670 = 10'h1a1 == _T_17 ? ram_417 : _GEN_5669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5671 = 10'h1a2 == _T_17 ? ram_418 : _GEN_5670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5672 = 10'h1a3 == _T_17 ? ram_419 : _GEN_5671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5673 = 10'h1a4 == _T_17 ? ram_420 : _GEN_5672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5674 = 10'h1a5 == _T_17 ? ram_421 : _GEN_5673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5675 = 10'h1a6 == _T_17 ? ram_422 : _GEN_5674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5676 = 10'h1a7 == _T_17 ? ram_423 : _GEN_5675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5677 = 10'h1a8 == _T_17 ? ram_424 : _GEN_5676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5678 = 10'h1a9 == _T_17 ? ram_425 : _GEN_5677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5679 = 10'h1aa == _T_17 ? ram_426 : _GEN_5678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5680 = 10'h1ab == _T_17 ? ram_427 : _GEN_5679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5681 = 10'h1ac == _T_17 ? ram_428 : _GEN_5680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5682 = 10'h1ad == _T_17 ? ram_429 : _GEN_5681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5683 = 10'h1ae == _T_17 ? ram_430 : _GEN_5682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5684 = 10'h1af == _T_17 ? ram_431 : _GEN_5683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5685 = 10'h1b0 == _T_17 ? ram_432 : _GEN_5684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5686 = 10'h1b1 == _T_17 ? ram_433 : _GEN_5685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5687 = 10'h1b2 == _T_17 ? ram_434 : _GEN_5686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5688 = 10'h1b3 == _T_17 ? ram_435 : _GEN_5687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5689 = 10'h1b4 == _T_17 ? ram_436 : _GEN_5688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5690 = 10'h1b5 == _T_17 ? ram_437 : _GEN_5689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5691 = 10'h1b6 == _T_17 ? ram_438 : _GEN_5690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5692 = 10'h1b7 == _T_17 ? ram_439 : _GEN_5691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5693 = 10'h1b8 == _T_17 ? ram_440 : _GEN_5692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5694 = 10'h1b9 == _T_17 ? ram_441 : _GEN_5693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5695 = 10'h1ba == _T_17 ? ram_442 : _GEN_5694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5696 = 10'h1bb == _T_17 ? ram_443 : _GEN_5695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5697 = 10'h1bc == _T_17 ? ram_444 : _GEN_5696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5698 = 10'h1bd == _T_17 ? ram_445 : _GEN_5697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5699 = 10'h1be == _T_17 ? ram_446 : _GEN_5698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5700 = 10'h1bf == _T_17 ? ram_447 : _GEN_5699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5701 = 10'h1c0 == _T_17 ? ram_448 : _GEN_5700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5702 = 10'h1c1 == _T_17 ? ram_449 : _GEN_5701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5703 = 10'h1c2 == _T_17 ? ram_450 : _GEN_5702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5704 = 10'h1c3 == _T_17 ? ram_451 : _GEN_5703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5705 = 10'h1c4 == _T_17 ? ram_452 : _GEN_5704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5706 = 10'h1c5 == _T_17 ? ram_453 : _GEN_5705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5707 = 10'h1c6 == _T_17 ? ram_454 : _GEN_5706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5708 = 10'h1c7 == _T_17 ? ram_455 : _GEN_5707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5709 = 10'h1c8 == _T_17 ? ram_456 : _GEN_5708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5710 = 10'h1c9 == _T_17 ? ram_457 : _GEN_5709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5711 = 10'h1ca == _T_17 ? ram_458 : _GEN_5710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5712 = 10'h1cb == _T_17 ? ram_459 : _GEN_5711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5713 = 10'h1cc == _T_17 ? ram_460 : _GEN_5712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5714 = 10'h1cd == _T_17 ? ram_461 : _GEN_5713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5715 = 10'h1ce == _T_17 ? ram_462 : _GEN_5714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5716 = 10'h1cf == _T_17 ? ram_463 : _GEN_5715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5717 = 10'h1d0 == _T_17 ? ram_464 : _GEN_5716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5718 = 10'h1d1 == _T_17 ? ram_465 : _GEN_5717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5719 = 10'h1d2 == _T_17 ? ram_466 : _GEN_5718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5720 = 10'h1d3 == _T_17 ? ram_467 : _GEN_5719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5721 = 10'h1d4 == _T_17 ? ram_468 : _GEN_5720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5722 = 10'h1d5 == _T_17 ? ram_469 : _GEN_5721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5723 = 10'h1d6 == _T_17 ? ram_470 : _GEN_5722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5724 = 10'h1d7 == _T_17 ? ram_471 : _GEN_5723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5725 = 10'h1d8 == _T_17 ? ram_472 : _GEN_5724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5726 = 10'h1d9 == _T_17 ? ram_473 : _GEN_5725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5727 = 10'h1da == _T_17 ? ram_474 : _GEN_5726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5728 = 10'h1db == _T_17 ? ram_475 : _GEN_5727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5729 = 10'h1dc == _T_17 ? ram_476 : _GEN_5728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5730 = 10'h1dd == _T_17 ? ram_477 : _GEN_5729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5731 = 10'h1de == _T_17 ? ram_478 : _GEN_5730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5732 = 10'h1df == _T_17 ? ram_479 : _GEN_5731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5733 = 10'h1e0 == _T_17 ? ram_480 : _GEN_5732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5734 = 10'h1e1 == _T_17 ? ram_481 : _GEN_5733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5735 = 10'h1e2 == _T_17 ? ram_482 : _GEN_5734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5736 = 10'h1e3 == _T_17 ? ram_483 : _GEN_5735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5737 = 10'h1e4 == _T_17 ? ram_484 : _GEN_5736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5738 = 10'h1e5 == _T_17 ? ram_485 : _GEN_5737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5739 = 10'h1e6 == _T_17 ? ram_486 : _GEN_5738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5740 = 10'h1e7 == _T_17 ? ram_487 : _GEN_5739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5741 = 10'h1e8 == _T_17 ? ram_488 : _GEN_5740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5742 = 10'h1e9 == _T_17 ? ram_489 : _GEN_5741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5743 = 10'h1ea == _T_17 ? ram_490 : _GEN_5742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5744 = 10'h1eb == _T_17 ? ram_491 : _GEN_5743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5745 = 10'h1ec == _T_17 ? ram_492 : _GEN_5744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5746 = 10'h1ed == _T_17 ? ram_493 : _GEN_5745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5747 = 10'h1ee == _T_17 ? ram_494 : _GEN_5746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5748 = 10'h1ef == _T_17 ? ram_495 : _GEN_5747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5749 = 10'h1f0 == _T_17 ? ram_496 : _GEN_5748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5750 = 10'h1f1 == _T_17 ? ram_497 : _GEN_5749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5751 = 10'h1f2 == _T_17 ? ram_498 : _GEN_5750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5752 = 10'h1f3 == _T_17 ? ram_499 : _GEN_5751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5753 = 10'h1f4 == _T_17 ? ram_500 : _GEN_5752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5754 = 10'h1f5 == _T_17 ? ram_501 : _GEN_5753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5755 = 10'h1f6 == _T_17 ? ram_502 : _GEN_5754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5756 = 10'h1f7 == _T_17 ? ram_503 : _GEN_5755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5757 = 10'h1f8 == _T_17 ? ram_504 : _GEN_5756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5758 = 10'h1f9 == _T_17 ? ram_505 : _GEN_5757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5759 = 10'h1fa == _T_17 ? ram_506 : _GEN_5758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5760 = 10'h1fb == _T_17 ? ram_507 : _GEN_5759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5761 = 10'h1fc == _T_17 ? ram_508 : _GEN_5760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5762 = 10'h1fd == _T_17 ? ram_509 : _GEN_5761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5763 = 10'h1fe == _T_17 ? ram_510 : _GEN_5762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5764 = 10'h1ff == _T_17 ? ram_511 : _GEN_5763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5765 = 10'h200 == _T_17 ? ram_512 : _GEN_5764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5766 = 10'h201 == _T_17 ? ram_513 : _GEN_5765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5767 = 10'h202 == _T_17 ? ram_514 : _GEN_5766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5768 = 10'h203 == _T_17 ? ram_515 : _GEN_5767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5769 = 10'h204 == _T_17 ? ram_516 : _GEN_5768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5770 = 10'h205 == _T_17 ? ram_517 : _GEN_5769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5771 = 10'h206 == _T_17 ? ram_518 : _GEN_5770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5772 = 10'h207 == _T_17 ? ram_519 : _GEN_5771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5773 = 10'h208 == _T_17 ? ram_520 : _GEN_5772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5774 = 10'h209 == _T_17 ? ram_521 : _GEN_5773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5775 = 10'h20a == _T_17 ? ram_522 : _GEN_5774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5776 = 10'h20b == _T_17 ? ram_523 : _GEN_5775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_5777 = 10'h20c == _T_17 ? ram_524 : _GEN_5776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19071 = {{8190'd0}, _GEN_5777}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_155 = _GEN_19071 ^ _ram_T_154; // @[vga.scala 64:41]
  wire [287:0] _GEN_5778 = 10'h0 == _T_17 ? _ram_T_155[287:0] : _GEN_4728; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5779 = 10'h1 == _T_17 ? _ram_T_155[287:0] : _GEN_4729; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5780 = 10'h2 == _T_17 ? _ram_T_155[287:0] : _GEN_4730; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5781 = 10'h3 == _T_17 ? _ram_T_155[287:0] : _GEN_4731; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5782 = 10'h4 == _T_17 ? _ram_T_155[287:0] : _GEN_4732; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5783 = 10'h5 == _T_17 ? _ram_T_155[287:0] : _GEN_4733; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5784 = 10'h6 == _T_17 ? _ram_T_155[287:0] : _GEN_4734; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5785 = 10'h7 == _T_17 ? _ram_T_155[287:0] : _GEN_4735; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5786 = 10'h8 == _T_17 ? _ram_T_155[287:0] : _GEN_4736; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5787 = 10'h9 == _T_17 ? _ram_T_155[287:0] : _GEN_4737; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5788 = 10'ha == _T_17 ? _ram_T_155[287:0] : _GEN_4738; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5789 = 10'hb == _T_17 ? _ram_T_155[287:0] : _GEN_4739; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5790 = 10'hc == _T_17 ? _ram_T_155[287:0] : _GEN_4740; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5791 = 10'hd == _T_17 ? _ram_T_155[287:0] : _GEN_4741; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5792 = 10'he == _T_17 ? _ram_T_155[287:0] : _GEN_4742; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5793 = 10'hf == _T_17 ? _ram_T_155[287:0] : _GEN_4743; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5794 = 10'h10 == _T_17 ? _ram_T_155[287:0] : _GEN_4744; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5795 = 10'h11 == _T_17 ? _ram_T_155[287:0] : _GEN_4745; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5796 = 10'h12 == _T_17 ? _ram_T_155[287:0] : _GEN_4746; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5797 = 10'h13 == _T_17 ? _ram_T_155[287:0] : _GEN_4747; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5798 = 10'h14 == _T_17 ? _ram_T_155[287:0] : _GEN_4748; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5799 = 10'h15 == _T_17 ? _ram_T_155[287:0] : _GEN_4749; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5800 = 10'h16 == _T_17 ? _ram_T_155[287:0] : _GEN_4750; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5801 = 10'h17 == _T_17 ? _ram_T_155[287:0] : _GEN_4751; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5802 = 10'h18 == _T_17 ? _ram_T_155[287:0] : _GEN_4752; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5803 = 10'h19 == _T_17 ? _ram_T_155[287:0] : _GEN_4753; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5804 = 10'h1a == _T_17 ? _ram_T_155[287:0] : _GEN_4754; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5805 = 10'h1b == _T_17 ? _ram_T_155[287:0] : _GEN_4755; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5806 = 10'h1c == _T_17 ? _ram_T_155[287:0] : _GEN_4756; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5807 = 10'h1d == _T_17 ? _ram_T_155[287:0] : _GEN_4757; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5808 = 10'h1e == _T_17 ? _ram_T_155[287:0] : _GEN_4758; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5809 = 10'h1f == _T_17 ? _ram_T_155[287:0] : _GEN_4759; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5810 = 10'h20 == _T_17 ? _ram_T_155[287:0] : _GEN_4760; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5811 = 10'h21 == _T_17 ? _ram_T_155[287:0] : _GEN_4761; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5812 = 10'h22 == _T_17 ? _ram_T_155[287:0] : _GEN_4762; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5813 = 10'h23 == _T_17 ? _ram_T_155[287:0] : _GEN_4763; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5814 = 10'h24 == _T_17 ? _ram_T_155[287:0] : _GEN_4764; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5815 = 10'h25 == _T_17 ? _ram_T_155[287:0] : _GEN_4765; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5816 = 10'h26 == _T_17 ? _ram_T_155[287:0] : _GEN_4766; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5817 = 10'h27 == _T_17 ? _ram_T_155[287:0] : _GEN_4767; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5818 = 10'h28 == _T_17 ? _ram_T_155[287:0] : _GEN_4768; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5819 = 10'h29 == _T_17 ? _ram_T_155[287:0] : _GEN_4769; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5820 = 10'h2a == _T_17 ? _ram_T_155[287:0] : _GEN_4770; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5821 = 10'h2b == _T_17 ? _ram_T_155[287:0] : _GEN_4771; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5822 = 10'h2c == _T_17 ? _ram_T_155[287:0] : _GEN_4772; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5823 = 10'h2d == _T_17 ? _ram_T_155[287:0] : _GEN_4773; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5824 = 10'h2e == _T_17 ? _ram_T_155[287:0] : _GEN_4774; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5825 = 10'h2f == _T_17 ? _ram_T_155[287:0] : _GEN_4775; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5826 = 10'h30 == _T_17 ? _ram_T_155[287:0] : _GEN_4776; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5827 = 10'h31 == _T_17 ? _ram_T_155[287:0] : _GEN_4777; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5828 = 10'h32 == _T_17 ? _ram_T_155[287:0] : _GEN_4778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5829 = 10'h33 == _T_17 ? _ram_T_155[287:0] : _GEN_4779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5830 = 10'h34 == _T_17 ? _ram_T_155[287:0] : _GEN_4780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5831 = 10'h35 == _T_17 ? _ram_T_155[287:0] : _GEN_4781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5832 = 10'h36 == _T_17 ? _ram_T_155[287:0] : _GEN_4782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5833 = 10'h37 == _T_17 ? _ram_T_155[287:0] : _GEN_4783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5834 = 10'h38 == _T_17 ? _ram_T_155[287:0] : _GEN_4784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5835 = 10'h39 == _T_17 ? _ram_T_155[287:0] : _GEN_4785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5836 = 10'h3a == _T_17 ? _ram_T_155[287:0] : _GEN_4786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5837 = 10'h3b == _T_17 ? _ram_T_155[287:0] : _GEN_4787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5838 = 10'h3c == _T_17 ? _ram_T_155[287:0] : _GEN_4788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5839 = 10'h3d == _T_17 ? _ram_T_155[287:0] : _GEN_4789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5840 = 10'h3e == _T_17 ? _ram_T_155[287:0] : _GEN_4790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5841 = 10'h3f == _T_17 ? _ram_T_155[287:0] : _GEN_4791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5842 = 10'h40 == _T_17 ? _ram_T_155[287:0] : _GEN_4792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5843 = 10'h41 == _T_17 ? _ram_T_155[287:0] : _GEN_4793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5844 = 10'h42 == _T_17 ? _ram_T_155[287:0] : _GEN_4794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5845 = 10'h43 == _T_17 ? _ram_T_155[287:0] : _GEN_4795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5846 = 10'h44 == _T_17 ? _ram_T_155[287:0] : _GEN_4796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5847 = 10'h45 == _T_17 ? _ram_T_155[287:0] : _GEN_4797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5848 = 10'h46 == _T_17 ? _ram_T_155[287:0] : _GEN_4798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5849 = 10'h47 == _T_17 ? _ram_T_155[287:0] : _GEN_4799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5850 = 10'h48 == _T_17 ? _ram_T_155[287:0] : _GEN_4800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5851 = 10'h49 == _T_17 ? _ram_T_155[287:0] : _GEN_4801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5852 = 10'h4a == _T_17 ? _ram_T_155[287:0] : _GEN_4802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5853 = 10'h4b == _T_17 ? _ram_T_155[287:0] : _GEN_4803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5854 = 10'h4c == _T_17 ? _ram_T_155[287:0] : _GEN_4804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5855 = 10'h4d == _T_17 ? _ram_T_155[287:0] : _GEN_4805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5856 = 10'h4e == _T_17 ? _ram_T_155[287:0] : _GEN_4806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5857 = 10'h4f == _T_17 ? _ram_T_155[287:0] : _GEN_4807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5858 = 10'h50 == _T_17 ? _ram_T_155[287:0] : _GEN_4808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5859 = 10'h51 == _T_17 ? _ram_T_155[287:0] : _GEN_4809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5860 = 10'h52 == _T_17 ? _ram_T_155[287:0] : _GEN_4810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5861 = 10'h53 == _T_17 ? _ram_T_155[287:0] : _GEN_4811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5862 = 10'h54 == _T_17 ? _ram_T_155[287:0] : _GEN_4812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5863 = 10'h55 == _T_17 ? _ram_T_155[287:0] : _GEN_4813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5864 = 10'h56 == _T_17 ? _ram_T_155[287:0] : _GEN_4814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5865 = 10'h57 == _T_17 ? _ram_T_155[287:0] : _GEN_4815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5866 = 10'h58 == _T_17 ? _ram_T_155[287:0] : _GEN_4816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5867 = 10'h59 == _T_17 ? _ram_T_155[287:0] : _GEN_4817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5868 = 10'h5a == _T_17 ? _ram_T_155[287:0] : _GEN_4818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5869 = 10'h5b == _T_17 ? _ram_T_155[287:0] : _GEN_4819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5870 = 10'h5c == _T_17 ? _ram_T_155[287:0] : _GEN_4820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5871 = 10'h5d == _T_17 ? _ram_T_155[287:0] : _GEN_4821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5872 = 10'h5e == _T_17 ? _ram_T_155[287:0] : _GEN_4822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5873 = 10'h5f == _T_17 ? _ram_T_155[287:0] : _GEN_4823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5874 = 10'h60 == _T_17 ? _ram_T_155[287:0] : _GEN_4824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5875 = 10'h61 == _T_17 ? _ram_T_155[287:0] : _GEN_4825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5876 = 10'h62 == _T_17 ? _ram_T_155[287:0] : _GEN_4826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5877 = 10'h63 == _T_17 ? _ram_T_155[287:0] : _GEN_4827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5878 = 10'h64 == _T_17 ? _ram_T_155[287:0] : _GEN_4828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5879 = 10'h65 == _T_17 ? _ram_T_155[287:0] : _GEN_4829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5880 = 10'h66 == _T_17 ? _ram_T_155[287:0] : _GEN_4830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5881 = 10'h67 == _T_17 ? _ram_T_155[287:0] : _GEN_4831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5882 = 10'h68 == _T_17 ? _ram_T_155[287:0] : _GEN_4832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5883 = 10'h69 == _T_17 ? _ram_T_155[287:0] : _GEN_4833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5884 = 10'h6a == _T_17 ? _ram_T_155[287:0] : _GEN_4834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5885 = 10'h6b == _T_17 ? _ram_T_155[287:0] : _GEN_4835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5886 = 10'h6c == _T_17 ? _ram_T_155[287:0] : _GEN_4836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5887 = 10'h6d == _T_17 ? _ram_T_155[287:0] : _GEN_4837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5888 = 10'h6e == _T_17 ? _ram_T_155[287:0] : _GEN_4838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5889 = 10'h6f == _T_17 ? _ram_T_155[287:0] : _GEN_4839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5890 = 10'h70 == _T_17 ? _ram_T_155[287:0] : _GEN_4840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5891 = 10'h71 == _T_17 ? _ram_T_155[287:0] : _GEN_4841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5892 = 10'h72 == _T_17 ? _ram_T_155[287:0] : _GEN_4842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5893 = 10'h73 == _T_17 ? _ram_T_155[287:0] : _GEN_4843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5894 = 10'h74 == _T_17 ? _ram_T_155[287:0] : _GEN_4844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5895 = 10'h75 == _T_17 ? _ram_T_155[287:0] : _GEN_4845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5896 = 10'h76 == _T_17 ? _ram_T_155[287:0] : _GEN_4846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5897 = 10'h77 == _T_17 ? _ram_T_155[287:0] : _GEN_4847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5898 = 10'h78 == _T_17 ? _ram_T_155[287:0] : _GEN_4848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5899 = 10'h79 == _T_17 ? _ram_T_155[287:0] : _GEN_4849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5900 = 10'h7a == _T_17 ? _ram_T_155[287:0] : _GEN_4850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5901 = 10'h7b == _T_17 ? _ram_T_155[287:0] : _GEN_4851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5902 = 10'h7c == _T_17 ? _ram_T_155[287:0] : _GEN_4852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5903 = 10'h7d == _T_17 ? _ram_T_155[287:0] : _GEN_4853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5904 = 10'h7e == _T_17 ? _ram_T_155[287:0] : _GEN_4854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5905 = 10'h7f == _T_17 ? _ram_T_155[287:0] : _GEN_4855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5906 = 10'h80 == _T_17 ? _ram_T_155[287:0] : _GEN_4856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5907 = 10'h81 == _T_17 ? _ram_T_155[287:0] : _GEN_4857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5908 = 10'h82 == _T_17 ? _ram_T_155[287:0] : _GEN_4858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5909 = 10'h83 == _T_17 ? _ram_T_155[287:0] : _GEN_4859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5910 = 10'h84 == _T_17 ? _ram_T_155[287:0] : _GEN_4860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5911 = 10'h85 == _T_17 ? _ram_T_155[287:0] : _GEN_4861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5912 = 10'h86 == _T_17 ? _ram_T_155[287:0] : _GEN_4862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5913 = 10'h87 == _T_17 ? _ram_T_155[287:0] : _GEN_4863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5914 = 10'h88 == _T_17 ? _ram_T_155[287:0] : _GEN_4864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5915 = 10'h89 == _T_17 ? _ram_T_155[287:0] : _GEN_4865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5916 = 10'h8a == _T_17 ? _ram_T_155[287:0] : _GEN_4866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5917 = 10'h8b == _T_17 ? _ram_T_155[287:0] : _GEN_4867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5918 = 10'h8c == _T_17 ? _ram_T_155[287:0] : _GEN_4868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5919 = 10'h8d == _T_17 ? _ram_T_155[287:0] : _GEN_4869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5920 = 10'h8e == _T_17 ? _ram_T_155[287:0] : _GEN_4870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5921 = 10'h8f == _T_17 ? _ram_T_155[287:0] : _GEN_4871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5922 = 10'h90 == _T_17 ? _ram_T_155[287:0] : _GEN_4872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5923 = 10'h91 == _T_17 ? _ram_T_155[287:0] : _GEN_4873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5924 = 10'h92 == _T_17 ? _ram_T_155[287:0] : _GEN_4874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5925 = 10'h93 == _T_17 ? _ram_T_155[287:0] : _GEN_4875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5926 = 10'h94 == _T_17 ? _ram_T_155[287:0] : _GEN_4876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5927 = 10'h95 == _T_17 ? _ram_T_155[287:0] : _GEN_4877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5928 = 10'h96 == _T_17 ? _ram_T_155[287:0] : _GEN_4878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5929 = 10'h97 == _T_17 ? _ram_T_155[287:0] : _GEN_4879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5930 = 10'h98 == _T_17 ? _ram_T_155[287:0] : _GEN_4880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5931 = 10'h99 == _T_17 ? _ram_T_155[287:0] : _GEN_4881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5932 = 10'h9a == _T_17 ? _ram_T_155[287:0] : _GEN_4882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5933 = 10'h9b == _T_17 ? _ram_T_155[287:0] : _GEN_4883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5934 = 10'h9c == _T_17 ? _ram_T_155[287:0] : _GEN_4884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5935 = 10'h9d == _T_17 ? _ram_T_155[287:0] : _GEN_4885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5936 = 10'h9e == _T_17 ? _ram_T_155[287:0] : _GEN_4886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5937 = 10'h9f == _T_17 ? _ram_T_155[287:0] : _GEN_4887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5938 = 10'ha0 == _T_17 ? _ram_T_155[287:0] : _GEN_4888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5939 = 10'ha1 == _T_17 ? _ram_T_155[287:0] : _GEN_4889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5940 = 10'ha2 == _T_17 ? _ram_T_155[287:0] : _GEN_4890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5941 = 10'ha3 == _T_17 ? _ram_T_155[287:0] : _GEN_4891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5942 = 10'ha4 == _T_17 ? _ram_T_155[287:0] : _GEN_4892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5943 = 10'ha5 == _T_17 ? _ram_T_155[287:0] : _GEN_4893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5944 = 10'ha6 == _T_17 ? _ram_T_155[287:0] : _GEN_4894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5945 = 10'ha7 == _T_17 ? _ram_T_155[287:0] : _GEN_4895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5946 = 10'ha8 == _T_17 ? _ram_T_155[287:0] : _GEN_4896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5947 = 10'ha9 == _T_17 ? _ram_T_155[287:0] : _GEN_4897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5948 = 10'haa == _T_17 ? _ram_T_155[287:0] : _GEN_4898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5949 = 10'hab == _T_17 ? _ram_T_155[287:0] : _GEN_4899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5950 = 10'hac == _T_17 ? _ram_T_155[287:0] : _GEN_4900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5951 = 10'had == _T_17 ? _ram_T_155[287:0] : _GEN_4901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5952 = 10'hae == _T_17 ? _ram_T_155[287:0] : _GEN_4902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5953 = 10'haf == _T_17 ? _ram_T_155[287:0] : _GEN_4903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5954 = 10'hb0 == _T_17 ? _ram_T_155[287:0] : _GEN_4904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5955 = 10'hb1 == _T_17 ? _ram_T_155[287:0] : _GEN_4905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5956 = 10'hb2 == _T_17 ? _ram_T_155[287:0] : _GEN_4906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5957 = 10'hb3 == _T_17 ? _ram_T_155[287:0] : _GEN_4907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5958 = 10'hb4 == _T_17 ? _ram_T_155[287:0] : _GEN_4908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5959 = 10'hb5 == _T_17 ? _ram_T_155[287:0] : _GEN_4909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5960 = 10'hb6 == _T_17 ? _ram_T_155[287:0] : _GEN_4910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5961 = 10'hb7 == _T_17 ? _ram_T_155[287:0] : _GEN_4911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5962 = 10'hb8 == _T_17 ? _ram_T_155[287:0] : _GEN_4912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5963 = 10'hb9 == _T_17 ? _ram_T_155[287:0] : _GEN_4913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5964 = 10'hba == _T_17 ? _ram_T_155[287:0] : _GEN_4914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5965 = 10'hbb == _T_17 ? _ram_T_155[287:0] : _GEN_4915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5966 = 10'hbc == _T_17 ? _ram_T_155[287:0] : _GEN_4916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5967 = 10'hbd == _T_17 ? _ram_T_155[287:0] : _GEN_4917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5968 = 10'hbe == _T_17 ? _ram_T_155[287:0] : _GEN_4918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5969 = 10'hbf == _T_17 ? _ram_T_155[287:0] : _GEN_4919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5970 = 10'hc0 == _T_17 ? _ram_T_155[287:0] : _GEN_4920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5971 = 10'hc1 == _T_17 ? _ram_T_155[287:0] : _GEN_4921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5972 = 10'hc2 == _T_17 ? _ram_T_155[287:0] : _GEN_4922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5973 = 10'hc3 == _T_17 ? _ram_T_155[287:0] : _GEN_4923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5974 = 10'hc4 == _T_17 ? _ram_T_155[287:0] : _GEN_4924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5975 = 10'hc5 == _T_17 ? _ram_T_155[287:0] : _GEN_4925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5976 = 10'hc6 == _T_17 ? _ram_T_155[287:0] : _GEN_4926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5977 = 10'hc7 == _T_17 ? _ram_T_155[287:0] : _GEN_4927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5978 = 10'hc8 == _T_17 ? _ram_T_155[287:0] : _GEN_4928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5979 = 10'hc9 == _T_17 ? _ram_T_155[287:0] : _GEN_4929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5980 = 10'hca == _T_17 ? _ram_T_155[287:0] : _GEN_4930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5981 = 10'hcb == _T_17 ? _ram_T_155[287:0] : _GEN_4931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5982 = 10'hcc == _T_17 ? _ram_T_155[287:0] : _GEN_4932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5983 = 10'hcd == _T_17 ? _ram_T_155[287:0] : _GEN_4933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5984 = 10'hce == _T_17 ? _ram_T_155[287:0] : _GEN_4934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5985 = 10'hcf == _T_17 ? _ram_T_155[287:0] : _GEN_4935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5986 = 10'hd0 == _T_17 ? _ram_T_155[287:0] : _GEN_4936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5987 = 10'hd1 == _T_17 ? _ram_T_155[287:0] : _GEN_4937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5988 = 10'hd2 == _T_17 ? _ram_T_155[287:0] : _GEN_4938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5989 = 10'hd3 == _T_17 ? _ram_T_155[287:0] : _GEN_4939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5990 = 10'hd4 == _T_17 ? _ram_T_155[287:0] : _GEN_4940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5991 = 10'hd5 == _T_17 ? _ram_T_155[287:0] : _GEN_4941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5992 = 10'hd6 == _T_17 ? _ram_T_155[287:0] : _GEN_4942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5993 = 10'hd7 == _T_17 ? _ram_T_155[287:0] : _GEN_4943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5994 = 10'hd8 == _T_17 ? _ram_T_155[287:0] : _GEN_4944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5995 = 10'hd9 == _T_17 ? _ram_T_155[287:0] : _GEN_4945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5996 = 10'hda == _T_17 ? _ram_T_155[287:0] : _GEN_4946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5997 = 10'hdb == _T_17 ? _ram_T_155[287:0] : _GEN_4947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5998 = 10'hdc == _T_17 ? _ram_T_155[287:0] : _GEN_4948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_5999 = 10'hdd == _T_17 ? _ram_T_155[287:0] : _GEN_4949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6000 = 10'hde == _T_17 ? _ram_T_155[287:0] : _GEN_4950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6001 = 10'hdf == _T_17 ? _ram_T_155[287:0] : _GEN_4951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6002 = 10'he0 == _T_17 ? _ram_T_155[287:0] : _GEN_4952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6003 = 10'he1 == _T_17 ? _ram_T_155[287:0] : _GEN_4953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6004 = 10'he2 == _T_17 ? _ram_T_155[287:0] : _GEN_4954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6005 = 10'he3 == _T_17 ? _ram_T_155[287:0] : _GEN_4955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6006 = 10'he4 == _T_17 ? _ram_T_155[287:0] : _GEN_4956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6007 = 10'he5 == _T_17 ? _ram_T_155[287:0] : _GEN_4957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6008 = 10'he6 == _T_17 ? _ram_T_155[287:0] : _GEN_4958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6009 = 10'he7 == _T_17 ? _ram_T_155[287:0] : _GEN_4959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6010 = 10'he8 == _T_17 ? _ram_T_155[287:0] : _GEN_4960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6011 = 10'he9 == _T_17 ? _ram_T_155[287:0] : _GEN_4961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6012 = 10'hea == _T_17 ? _ram_T_155[287:0] : _GEN_4962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6013 = 10'heb == _T_17 ? _ram_T_155[287:0] : _GEN_4963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6014 = 10'hec == _T_17 ? _ram_T_155[287:0] : _GEN_4964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6015 = 10'hed == _T_17 ? _ram_T_155[287:0] : _GEN_4965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6016 = 10'hee == _T_17 ? _ram_T_155[287:0] : _GEN_4966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6017 = 10'hef == _T_17 ? _ram_T_155[287:0] : _GEN_4967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6018 = 10'hf0 == _T_17 ? _ram_T_155[287:0] : _GEN_4968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6019 = 10'hf1 == _T_17 ? _ram_T_155[287:0] : _GEN_4969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6020 = 10'hf2 == _T_17 ? _ram_T_155[287:0] : _GEN_4970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6021 = 10'hf3 == _T_17 ? _ram_T_155[287:0] : _GEN_4971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6022 = 10'hf4 == _T_17 ? _ram_T_155[287:0] : _GEN_4972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6023 = 10'hf5 == _T_17 ? _ram_T_155[287:0] : _GEN_4973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6024 = 10'hf6 == _T_17 ? _ram_T_155[287:0] : _GEN_4974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6025 = 10'hf7 == _T_17 ? _ram_T_155[287:0] : _GEN_4975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6026 = 10'hf8 == _T_17 ? _ram_T_155[287:0] : _GEN_4976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6027 = 10'hf9 == _T_17 ? _ram_T_155[287:0] : _GEN_4977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6028 = 10'hfa == _T_17 ? _ram_T_155[287:0] : _GEN_4978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6029 = 10'hfb == _T_17 ? _ram_T_155[287:0] : _GEN_4979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6030 = 10'hfc == _T_17 ? _ram_T_155[287:0] : _GEN_4980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6031 = 10'hfd == _T_17 ? _ram_T_155[287:0] : _GEN_4981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6032 = 10'hfe == _T_17 ? _ram_T_155[287:0] : _GEN_4982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6033 = 10'hff == _T_17 ? _ram_T_155[287:0] : _GEN_4983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6034 = 10'h100 == _T_17 ? _ram_T_155[287:0] : _GEN_4984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6035 = 10'h101 == _T_17 ? _ram_T_155[287:0] : _GEN_4985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6036 = 10'h102 == _T_17 ? _ram_T_155[287:0] : _GEN_4986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6037 = 10'h103 == _T_17 ? _ram_T_155[287:0] : _GEN_4987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6038 = 10'h104 == _T_17 ? _ram_T_155[287:0] : _GEN_4988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6039 = 10'h105 == _T_17 ? _ram_T_155[287:0] : _GEN_4989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6040 = 10'h106 == _T_17 ? _ram_T_155[287:0] : _GEN_4990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6041 = 10'h107 == _T_17 ? _ram_T_155[287:0] : _GEN_4991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6042 = 10'h108 == _T_17 ? _ram_T_155[287:0] : _GEN_4992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6043 = 10'h109 == _T_17 ? _ram_T_155[287:0] : _GEN_4993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6044 = 10'h10a == _T_17 ? _ram_T_155[287:0] : _GEN_4994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6045 = 10'h10b == _T_17 ? _ram_T_155[287:0] : _GEN_4995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6046 = 10'h10c == _T_17 ? _ram_T_155[287:0] : _GEN_4996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6047 = 10'h10d == _T_17 ? _ram_T_155[287:0] : _GEN_4997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6048 = 10'h10e == _T_17 ? _ram_T_155[287:0] : _GEN_4998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6049 = 10'h10f == _T_17 ? _ram_T_155[287:0] : _GEN_4999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6050 = 10'h110 == _T_17 ? _ram_T_155[287:0] : _GEN_5000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6051 = 10'h111 == _T_17 ? _ram_T_155[287:0] : _GEN_5001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6052 = 10'h112 == _T_17 ? _ram_T_155[287:0] : _GEN_5002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6053 = 10'h113 == _T_17 ? _ram_T_155[287:0] : _GEN_5003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6054 = 10'h114 == _T_17 ? _ram_T_155[287:0] : _GEN_5004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6055 = 10'h115 == _T_17 ? _ram_T_155[287:0] : _GEN_5005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6056 = 10'h116 == _T_17 ? _ram_T_155[287:0] : _GEN_5006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6057 = 10'h117 == _T_17 ? _ram_T_155[287:0] : _GEN_5007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6058 = 10'h118 == _T_17 ? _ram_T_155[287:0] : _GEN_5008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6059 = 10'h119 == _T_17 ? _ram_T_155[287:0] : _GEN_5009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6060 = 10'h11a == _T_17 ? _ram_T_155[287:0] : _GEN_5010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6061 = 10'h11b == _T_17 ? _ram_T_155[287:0] : _GEN_5011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6062 = 10'h11c == _T_17 ? _ram_T_155[287:0] : _GEN_5012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6063 = 10'h11d == _T_17 ? _ram_T_155[287:0] : _GEN_5013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6064 = 10'h11e == _T_17 ? _ram_T_155[287:0] : _GEN_5014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6065 = 10'h11f == _T_17 ? _ram_T_155[287:0] : _GEN_5015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6066 = 10'h120 == _T_17 ? _ram_T_155[287:0] : _GEN_5016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6067 = 10'h121 == _T_17 ? _ram_T_155[287:0] : _GEN_5017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6068 = 10'h122 == _T_17 ? _ram_T_155[287:0] : _GEN_5018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6069 = 10'h123 == _T_17 ? _ram_T_155[287:0] : _GEN_5019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6070 = 10'h124 == _T_17 ? _ram_T_155[287:0] : _GEN_5020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6071 = 10'h125 == _T_17 ? _ram_T_155[287:0] : _GEN_5021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6072 = 10'h126 == _T_17 ? _ram_T_155[287:0] : _GEN_5022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6073 = 10'h127 == _T_17 ? _ram_T_155[287:0] : _GEN_5023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6074 = 10'h128 == _T_17 ? _ram_T_155[287:0] : _GEN_5024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6075 = 10'h129 == _T_17 ? _ram_T_155[287:0] : _GEN_5025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6076 = 10'h12a == _T_17 ? _ram_T_155[287:0] : _GEN_5026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6077 = 10'h12b == _T_17 ? _ram_T_155[287:0] : _GEN_5027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6078 = 10'h12c == _T_17 ? _ram_T_155[287:0] : _GEN_5028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6079 = 10'h12d == _T_17 ? _ram_T_155[287:0] : _GEN_5029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6080 = 10'h12e == _T_17 ? _ram_T_155[287:0] : _GEN_5030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6081 = 10'h12f == _T_17 ? _ram_T_155[287:0] : _GEN_5031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6082 = 10'h130 == _T_17 ? _ram_T_155[287:0] : _GEN_5032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6083 = 10'h131 == _T_17 ? _ram_T_155[287:0] : _GEN_5033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6084 = 10'h132 == _T_17 ? _ram_T_155[287:0] : _GEN_5034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6085 = 10'h133 == _T_17 ? _ram_T_155[287:0] : _GEN_5035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6086 = 10'h134 == _T_17 ? _ram_T_155[287:0] : _GEN_5036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6087 = 10'h135 == _T_17 ? _ram_T_155[287:0] : _GEN_5037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6088 = 10'h136 == _T_17 ? _ram_T_155[287:0] : _GEN_5038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6089 = 10'h137 == _T_17 ? _ram_T_155[287:0] : _GEN_5039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6090 = 10'h138 == _T_17 ? _ram_T_155[287:0] : _GEN_5040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6091 = 10'h139 == _T_17 ? _ram_T_155[287:0] : _GEN_5041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6092 = 10'h13a == _T_17 ? _ram_T_155[287:0] : _GEN_5042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6093 = 10'h13b == _T_17 ? _ram_T_155[287:0] : _GEN_5043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6094 = 10'h13c == _T_17 ? _ram_T_155[287:0] : _GEN_5044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6095 = 10'h13d == _T_17 ? _ram_T_155[287:0] : _GEN_5045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6096 = 10'h13e == _T_17 ? _ram_T_155[287:0] : _GEN_5046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6097 = 10'h13f == _T_17 ? _ram_T_155[287:0] : _GEN_5047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6098 = 10'h140 == _T_17 ? _ram_T_155[287:0] : _GEN_5048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6099 = 10'h141 == _T_17 ? _ram_T_155[287:0] : _GEN_5049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6100 = 10'h142 == _T_17 ? _ram_T_155[287:0] : _GEN_5050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6101 = 10'h143 == _T_17 ? _ram_T_155[287:0] : _GEN_5051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6102 = 10'h144 == _T_17 ? _ram_T_155[287:0] : _GEN_5052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6103 = 10'h145 == _T_17 ? _ram_T_155[287:0] : _GEN_5053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6104 = 10'h146 == _T_17 ? _ram_T_155[287:0] : _GEN_5054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6105 = 10'h147 == _T_17 ? _ram_T_155[287:0] : _GEN_5055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6106 = 10'h148 == _T_17 ? _ram_T_155[287:0] : _GEN_5056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6107 = 10'h149 == _T_17 ? _ram_T_155[287:0] : _GEN_5057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6108 = 10'h14a == _T_17 ? _ram_T_155[287:0] : _GEN_5058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6109 = 10'h14b == _T_17 ? _ram_T_155[287:0] : _GEN_5059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6110 = 10'h14c == _T_17 ? _ram_T_155[287:0] : _GEN_5060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6111 = 10'h14d == _T_17 ? _ram_T_155[287:0] : _GEN_5061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6112 = 10'h14e == _T_17 ? _ram_T_155[287:0] : _GEN_5062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6113 = 10'h14f == _T_17 ? _ram_T_155[287:0] : _GEN_5063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6114 = 10'h150 == _T_17 ? _ram_T_155[287:0] : _GEN_5064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6115 = 10'h151 == _T_17 ? _ram_T_155[287:0] : _GEN_5065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6116 = 10'h152 == _T_17 ? _ram_T_155[287:0] : _GEN_5066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6117 = 10'h153 == _T_17 ? _ram_T_155[287:0] : _GEN_5067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6118 = 10'h154 == _T_17 ? _ram_T_155[287:0] : _GEN_5068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6119 = 10'h155 == _T_17 ? _ram_T_155[287:0] : _GEN_5069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6120 = 10'h156 == _T_17 ? _ram_T_155[287:0] : _GEN_5070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6121 = 10'h157 == _T_17 ? _ram_T_155[287:0] : _GEN_5071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6122 = 10'h158 == _T_17 ? _ram_T_155[287:0] : _GEN_5072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6123 = 10'h159 == _T_17 ? _ram_T_155[287:0] : _GEN_5073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6124 = 10'h15a == _T_17 ? _ram_T_155[287:0] : _GEN_5074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6125 = 10'h15b == _T_17 ? _ram_T_155[287:0] : _GEN_5075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6126 = 10'h15c == _T_17 ? _ram_T_155[287:0] : _GEN_5076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6127 = 10'h15d == _T_17 ? _ram_T_155[287:0] : _GEN_5077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6128 = 10'h15e == _T_17 ? _ram_T_155[287:0] : _GEN_5078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6129 = 10'h15f == _T_17 ? _ram_T_155[287:0] : _GEN_5079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6130 = 10'h160 == _T_17 ? _ram_T_155[287:0] : _GEN_5080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6131 = 10'h161 == _T_17 ? _ram_T_155[287:0] : _GEN_5081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6132 = 10'h162 == _T_17 ? _ram_T_155[287:0] : _GEN_5082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6133 = 10'h163 == _T_17 ? _ram_T_155[287:0] : _GEN_5083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6134 = 10'h164 == _T_17 ? _ram_T_155[287:0] : _GEN_5084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6135 = 10'h165 == _T_17 ? _ram_T_155[287:0] : _GEN_5085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6136 = 10'h166 == _T_17 ? _ram_T_155[287:0] : _GEN_5086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6137 = 10'h167 == _T_17 ? _ram_T_155[287:0] : _GEN_5087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6138 = 10'h168 == _T_17 ? _ram_T_155[287:0] : _GEN_5088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6139 = 10'h169 == _T_17 ? _ram_T_155[287:0] : _GEN_5089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6140 = 10'h16a == _T_17 ? _ram_T_155[287:0] : _GEN_5090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6141 = 10'h16b == _T_17 ? _ram_T_155[287:0] : _GEN_5091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6142 = 10'h16c == _T_17 ? _ram_T_155[287:0] : _GEN_5092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6143 = 10'h16d == _T_17 ? _ram_T_155[287:0] : _GEN_5093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6144 = 10'h16e == _T_17 ? _ram_T_155[287:0] : _GEN_5094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6145 = 10'h16f == _T_17 ? _ram_T_155[287:0] : _GEN_5095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6146 = 10'h170 == _T_17 ? _ram_T_155[287:0] : _GEN_5096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6147 = 10'h171 == _T_17 ? _ram_T_155[287:0] : _GEN_5097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6148 = 10'h172 == _T_17 ? _ram_T_155[287:0] : _GEN_5098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6149 = 10'h173 == _T_17 ? _ram_T_155[287:0] : _GEN_5099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6150 = 10'h174 == _T_17 ? _ram_T_155[287:0] : _GEN_5100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6151 = 10'h175 == _T_17 ? _ram_T_155[287:0] : _GEN_5101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6152 = 10'h176 == _T_17 ? _ram_T_155[287:0] : _GEN_5102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6153 = 10'h177 == _T_17 ? _ram_T_155[287:0] : _GEN_5103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6154 = 10'h178 == _T_17 ? _ram_T_155[287:0] : _GEN_5104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6155 = 10'h179 == _T_17 ? _ram_T_155[287:0] : _GEN_5105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6156 = 10'h17a == _T_17 ? _ram_T_155[287:0] : _GEN_5106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6157 = 10'h17b == _T_17 ? _ram_T_155[287:0] : _GEN_5107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6158 = 10'h17c == _T_17 ? _ram_T_155[287:0] : _GEN_5108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6159 = 10'h17d == _T_17 ? _ram_T_155[287:0] : _GEN_5109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6160 = 10'h17e == _T_17 ? _ram_T_155[287:0] : _GEN_5110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6161 = 10'h17f == _T_17 ? _ram_T_155[287:0] : _GEN_5111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6162 = 10'h180 == _T_17 ? _ram_T_155[287:0] : _GEN_5112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6163 = 10'h181 == _T_17 ? _ram_T_155[287:0] : _GEN_5113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6164 = 10'h182 == _T_17 ? _ram_T_155[287:0] : _GEN_5114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6165 = 10'h183 == _T_17 ? _ram_T_155[287:0] : _GEN_5115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6166 = 10'h184 == _T_17 ? _ram_T_155[287:0] : _GEN_5116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6167 = 10'h185 == _T_17 ? _ram_T_155[287:0] : _GEN_5117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6168 = 10'h186 == _T_17 ? _ram_T_155[287:0] : _GEN_5118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6169 = 10'h187 == _T_17 ? _ram_T_155[287:0] : _GEN_5119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6170 = 10'h188 == _T_17 ? _ram_T_155[287:0] : _GEN_5120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6171 = 10'h189 == _T_17 ? _ram_T_155[287:0] : _GEN_5121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6172 = 10'h18a == _T_17 ? _ram_T_155[287:0] : _GEN_5122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6173 = 10'h18b == _T_17 ? _ram_T_155[287:0] : _GEN_5123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6174 = 10'h18c == _T_17 ? _ram_T_155[287:0] : _GEN_5124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6175 = 10'h18d == _T_17 ? _ram_T_155[287:0] : _GEN_5125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6176 = 10'h18e == _T_17 ? _ram_T_155[287:0] : _GEN_5126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6177 = 10'h18f == _T_17 ? _ram_T_155[287:0] : _GEN_5127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6178 = 10'h190 == _T_17 ? _ram_T_155[287:0] : _GEN_5128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6179 = 10'h191 == _T_17 ? _ram_T_155[287:0] : _GEN_5129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6180 = 10'h192 == _T_17 ? _ram_T_155[287:0] : _GEN_5130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6181 = 10'h193 == _T_17 ? _ram_T_155[287:0] : _GEN_5131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6182 = 10'h194 == _T_17 ? _ram_T_155[287:0] : _GEN_5132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6183 = 10'h195 == _T_17 ? _ram_T_155[287:0] : _GEN_5133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6184 = 10'h196 == _T_17 ? _ram_T_155[287:0] : _GEN_5134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6185 = 10'h197 == _T_17 ? _ram_T_155[287:0] : _GEN_5135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6186 = 10'h198 == _T_17 ? _ram_T_155[287:0] : _GEN_5136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6187 = 10'h199 == _T_17 ? _ram_T_155[287:0] : _GEN_5137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6188 = 10'h19a == _T_17 ? _ram_T_155[287:0] : _GEN_5138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6189 = 10'h19b == _T_17 ? _ram_T_155[287:0] : _GEN_5139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6190 = 10'h19c == _T_17 ? _ram_T_155[287:0] : _GEN_5140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6191 = 10'h19d == _T_17 ? _ram_T_155[287:0] : _GEN_5141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6192 = 10'h19e == _T_17 ? _ram_T_155[287:0] : _GEN_5142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6193 = 10'h19f == _T_17 ? _ram_T_155[287:0] : _GEN_5143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6194 = 10'h1a0 == _T_17 ? _ram_T_155[287:0] : _GEN_5144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6195 = 10'h1a1 == _T_17 ? _ram_T_155[287:0] : _GEN_5145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6196 = 10'h1a2 == _T_17 ? _ram_T_155[287:0] : _GEN_5146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6197 = 10'h1a3 == _T_17 ? _ram_T_155[287:0] : _GEN_5147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6198 = 10'h1a4 == _T_17 ? _ram_T_155[287:0] : _GEN_5148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6199 = 10'h1a5 == _T_17 ? _ram_T_155[287:0] : _GEN_5149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6200 = 10'h1a6 == _T_17 ? _ram_T_155[287:0] : _GEN_5150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6201 = 10'h1a7 == _T_17 ? _ram_T_155[287:0] : _GEN_5151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6202 = 10'h1a8 == _T_17 ? _ram_T_155[287:0] : _GEN_5152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6203 = 10'h1a9 == _T_17 ? _ram_T_155[287:0] : _GEN_5153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6204 = 10'h1aa == _T_17 ? _ram_T_155[287:0] : _GEN_5154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6205 = 10'h1ab == _T_17 ? _ram_T_155[287:0] : _GEN_5155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6206 = 10'h1ac == _T_17 ? _ram_T_155[287:0] : _GEN_5156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6207 = 10'h1ad == _T_17 ? _ram_T_155[287:0] : _GEN_5157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6208 = 10'h1ae == _T_17 ? _ram_T_155[287:0] : _GEN_5158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6209 = 10'h1af == _T_17 ? _ram_T_155[287:0] : _GEN_5159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6210 = 10'h1b0 == _T_17 ? _ram_T_155[287:0] : _GEN_5160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6211 = 10'h1b1 == _T_17 ? _ram_T_155[287:0] : _GEN_5161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6212 = 10'h1b2 == _T_17 ? _ram_T_155[287:0] : _GEN_5162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6213 = 10'h1b3 == _T_17 ? _ram_T_155[287:0] : _GEN_5163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6214 = 10'h1b4 == _T_17 ? _ram_T_155[287:0] : _GEN_5164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6215 = 10'h1b5 == _T_17 ? _ram_T_155[287:0] : _GEN_5165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6216 = 10'h1b6 == _T_17 ? _ram_T_155[287:0] : _GEN_5166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6217 = 10'h1b7 == _T_17 ? _ram_T_155[287:0] : _GEN_5167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6218 = 10'h1b8 == _T_17 ? _ram_T_155[287:0] : _GEN_5168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6219 = 10'h1b9 == _T_17 ? _ram_T_155[287:0] : _GEN_5169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6220 = 10'h1ba == _T_17 ? _ram_T_155[287:0] : _GEN_5170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6221 = 10'h1bb == _T_17 ? _ram_T_155[287:0] : _GEN_5171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6222 = 10'h1bc == _T_17 ? _ram_T_155[287:0] : _GEN_5172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6223 = 10'h1bd == _T_17 ? _ram_T_155[287:0] : _GEN_5173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6224 = 10'h1be == _T_17 ? _ram_T_155[287:0] : _GEN_5174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6225 = 10'h1bf == _T_17 ? _ram_T_155[287:0] : _GEN_5175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6226 = 10'h1c0 == _T_17 ? _ram_T_155[287:0] : _GEN_5176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6227 = 10'h1c1 == _T_17 ? _ram_T_155[287:0] : _GEN_5177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6228 = 10'h1c2 == _T_17 ? _ram_T_155[287:0] : _GEN_5178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6229 = 10'h1c3 == _T_17 ? _ram_T_155[287:0] : _GEN_5179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6230 = 10'h1c4 == _T_17 ? _ram_T_155[287:0] : _GEN_5180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6231 = 10'h1c5 == _T_17 ? _ram_T_155[287:0] : _GEN_5181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6232 = 10'h1c6 == _T_17 ? _ram_T_155[287:0] : _GEN_5182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6233 = 10'h1c7 == _T_17 ? _ram_T_155[287:0] : _GEN_5183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6234 = 10'h1c8 == _T_17 ? _ram_T_155[287:0] : _GEN_5184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6235 = 10'h1c9 == _T_17 ? _ram_T_155[287:0] : _GEN_5185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6236 = 10'h1ca == _T_17 ? _ram_T_155[287:0] : _GEN_5186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6237 = 10'h1cb == _T_17 ? _ram_T_155[287:0] : _GEN_5187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6238 = 10'h1cc == _T_17 ? _ram_T_155[287:0] : _GEN_5188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6239 = 10'h1cd == _T_17 ? _ram_T_155[287:0] : _GEN_5189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6240 = 10'h1ce == _T_17 ? _ram_T_155[287:0] : _GEN_5190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6241 = 10'h1cf == _T_17 ? _ram_T_155[287:0] : _GEN_5191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6242 = 10'h1d0 == _T_17 ? _ram_T_155[287:0] : _GEN_5192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6243 = 10'h1d1 == _T_17 ? _ram_T_155[287:0] : _GEN_5193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6244 = 10'h1d2 == _T_17 ? _ram_T_155[287:0] : _GEN_5194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6245 = 10'h1d3 == _T_17 ? _ram_T_155[287:0] : _GEN_5195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6246 = 10'h1d4 == _T_17 ? _ram_T_155[287:0] : _GEN_5196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6247 = 10'h1d5 == _T_17 ? _ram_T_155[287:0] : _GEN_5197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6248 = 10'h1d6 == _T_17 ? _ram_T_155[287:0] : _GEN_5198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6249 = 10'h1d7 == _T_17 ? _ram_T_155[287:0] : _GEN_5199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6250 = 10'h1d8 == _T_17 ? _ram_T_155[287:0] : _GEN_5200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6251 = 10'h1d9 == _T_17 ? _ram_T_155[287:0] : _GEN_5201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6252 = 10'h1da == _T_17 ? _ram_T_155[287:0] : _GEN_5202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6253 = 10'h1db == _T_17 ? _ram_T_155[287:0] : _GEN_5203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6254 = 10'h1dc == _T_17 ? _ram_T_155[287:0] : _GEN_5204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6255 = 10'h1dd == _T_17 ? _ram_T_155[287:0] : _GEN_5205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6256 = 10'h1de == _T_17 ? _ram_T_155[287:0] : _GEN_5206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6257 = 10'h1df == _T_17 ? _ram_T_155[287:0] : _GEN_5207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6258 = 10'h1e0 == _T_17 ? _ram_T_155[287:0] : _GEN_5208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6259 = 10'h1e1 == _T_17 ? _ram_T_155[287:0] : _GEN_5209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6260 = 10'h1e2 == _T_17 ? _ram_T_155[287:0] : _GEN_5210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6261 = 10'h1e3 == _T_17 ? _ram_T_155[287:0] : _GEN_5211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6262 = 10'h1e4 == _T_17 ? _ram_T_155[287:0] : _GEN_5212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6263 = 10'h1e5 == _T_17 ? _ram_T_155[287:0] : _GEN_5213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6264 = 10'h1e6 == _T_17 ? _ram_T_155[287:0] : _GEN_5214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6265 = 10'h1e7 == _T_17 ? _ram_T_155[287:0] : _GEN_5215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6266 = 10'h1e8 == _T_17 ? _ram_T_155[287:0] : _GEN_5216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6267 = 10'h1e9 == _T_17 ? _ram_T_155[287:0] : _GEN_5217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6268 = 10'h1ea == _T_17 ? _ram_T_155[287:0] : _GEN_5218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6269 = 10'h1eb == _T_17 ? _ram_T_155[287:0] : _GEN_5219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6270 = 10'h1ec == _T_17 ? _ram_T_155[287:0] : _GEN_5220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6271 = 10'h1ed == _T_17 ? _ram_T_155[287:0] : _GEN_5221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6272 = 10'h1ee == _T_17 ? _ram_T_155[287:0] : _GEN_5222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6273 = 10'h1ef == _T_17 ? _ram_T_155[287:0] : _GEN_5223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6274 = 10'h1f0 == _T_17 ? _ram_T_155[287:0] : _GEN_5224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6275 = 10'h1f1 == _T_17 ? _ram_T_155[287:0] : _GEN_5225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6276 = 10'h1f2 == _T_17 ? _ram_T_155[287:0] : _GEN_5226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6277 = 10'h1f3 == _T_17 ? _ram_T_155[287:0] : _GEN_5227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6278 = 10'h1f4 == _T_17 ? _ram_T_155[287:0] : _GEN_5228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6279 = 10'h1f5 == _T_17 ? _ram_T_155[287:0] : _GEN_5229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6280 = 10'h1f6 == _T_17 ? _ram_T_155[287:0] : _GEN_5230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6281 = 10'h1f7 == _T_17 ? _ram_T_155[287:0] : _GEN_5231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6282 = 10'h1f8 == _T_17 ? _ram_T_155[287:0] : _GEN_5232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6283 = 10'h1f9 == _T_17 ? _ram_T_155[287:0] : _GEN_5233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6284 = 10'h1fa == _T_17 ? _ram_T_155[287:0] : _GEN_5234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6285 = 10'h1fb == _T_17 ? _ram_T_155[287:0] : _GEN_5235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6286 = 10'h1fc == _T_17 ? _ram_T_155[287:0] : _GEN_5236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6287 = 10'h1fd == _T_17 ? _ram_T_155[287:0] : _GEN_5237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6288 = 10'h1fe == _T_17 ? _ram_T_155[287:0] : _GEN_5238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6289 = 10'h1ff == _T_17 ? _ram_T_155[287:0] : _GEN_5239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6290 = 10'h200 == _T_17 ? _ram_T_155[287:0] : _GEN_5240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6291 = 10'h201 == _T_17 ? _ram_T_155[287:0] : _GEN_5241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6292 = 10'h202 == _T_17 ? _ram_T_155[287:0] : _GEN_5242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6293 = 10'h203 == _T_17 ? _ram_T_155[287:0] : _GEN_5243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6294 = 10'h204 == _T_17 ? _ram_T_155[287:0] : _GEN_5244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6295 = 10'h205 == _T_17 ? _ram_T_155[287:0] : _GEN_5245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6296 = 10'h206 == _T_17 ? _ram_T_155[287:0] : _GEN_5246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6297 = 10'h207 == _T_17 ? _ram_T_155[287:0] : _GEN_5247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6298 = 10'h208 == _T_17 ? _ram_T_155[287:0] : _GEN_5248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6299 = 10'h209 == _T_17 ? _ram_T_155[287:0] : _GEN_5249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6300 = 10'h20a == _T_17 ? _ram_T_155[287:0] : _GEN_5250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6301 = 10'h20b == _T_17 ? _ram_T_155[287:0] : _GEN_5251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6302 = 10'h20c == _T_17 ? _ram_T_155[287:0] : _GEN_5252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_19 = h + 10'h6; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_6 = vga_mem_ram_MPORT_54_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_6 = vga_mem_ram_MPORT_55_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_6 = vga_mem_ram_MPORT_56_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_6 = vga_mem_ram_MPORT_57_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_6 = vga_mem_ram_MPORT_58_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_6 = vga_mem_ram_MPORT_59_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_6 = vga_mem_ram_MPORT_60_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_6 = vga_mem_ram_MPORT_61_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_6 = vga_mem_ram_MPORT_62_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_176 = {278'h0,ram_hi_hi_hi_lo_6,ram_hi_hi_lo_6,ram_hi_lo_hi_6,ram_hi_lo_lo_6,ram_lo_hi_hi_hi_6,
    ram_lo_hi_hi_lo_6,ram_lo_hi_lo_6,ram_lo_lo_hi_6,ram_lo_lo_lo_6}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19072 = {{8191'd0}, _ram_T_176}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_180 = _GEN_19072 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_6304 = 10'h1 == _T_19 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6305 = 10'h2 == _T_19 ? ram_2 : _GEN_6304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6306 = 10'h3 == _T_19 ? ram_3 : _GEN_6305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6307 = 10'h4 == _T_19 ? ram_4 : _GEN_6306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6308 = 10'h5 == _T_19 ? ram_5 : _GEN_6307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6309 = 10'h6 == _T_19 ? ram_6 : _GEN_6308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6310 = 10'h7 == _T_19 ? ram_7 : _GEN_6309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6311 = 10'h8 == _T_19 ? ram_8 : _GEN_6310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6312 = 10'h9 == _T_19 ? ram_9 : _GEN_6311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6313 = 10'ha == _T_19 ? ram_10 : _GEN_6312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6314 = 10'hb == _T_19 ? ram_11 : _GEN_6313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6315 = 10'hc == _T_19 ? ram_12 : _GEN_6314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6316 = 10'hd == _T_19 ? ram_13 : _GEN_6315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6317 = 10'he == _T_19 ? ram_14 : _GEN_6316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6318 = 10'hf == _T_19 ? ram_15 : _GEN_6317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6319 = 10'h10 == _T_19 ? ram_16 : _GEN_6318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6320 = 10'h11 == _T_19 ? ram_17 : _GEN_6319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6321 = 10'h12 == _T_19 ? ram_18 : _GEN_6320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6322 = 10'h13 == _T_19 ? ram_19 : _GEN_6321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6323 = 10'h14 == _T_19 ? ram_20 : _GEN_6322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6324 = 10'h15 == _T_19 ? ram_21 : _GEN_6323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6325 = 10'h16 == _T_19 ? ram_22 : _GEN_6324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6326 = 10'h17 == _T_19 ? ram_23 : _GEN_6325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6327 = 10'h18 == _T_19 ? ram_24 : _GEN_6326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6328 = 10'h19 == _T_19 ? ram_25 : _GEN_6327; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6329 = 10'h1a == _T_19 ? ram_26 : _GEN_6328; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6330 = 10'h1b == _T_19 ? ram_27 : _GEN_6329; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6331 = 10'h1c == _T_19 ? ram_28 : _GEN_6330; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6332 = 10'h1d == _T_19 ? ram_29 : _GEN_6331; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6333 = 10'h1e == _T_19 ? ram_30 : _GEN_6332; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6334 = 10'h1f == _T_19 ? ram_31 : _GEN_6333; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6335 = 10'h20 == _T_19 ? ram_32 : _GEN_6334; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6336 = 10'h21 == _T_19 ? ram_33 : _GEN_6335; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6337 = 10'h22 == _T_19 ? ram_34 : _GEN_6336; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6338 = 10'h23 == _T_19 ? ram_35 : _GEN_6337; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6339 = 10'h24 == _T_19 ? ram_36 : _GEN_6338; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6340 = 10'h25 == _T_19 ? ram_37 : _GEN_6339; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6341 = 10'h26 == _T_19 ? ram_38 : _GEN_6340; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6342 = 10'h27 == _T_19 ? ram_39 : _GEN_6341; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6343 = 10'h28 == _T_19 ? ram_40 : _GEN_6342; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6344 = 10'h29 == _T_19 ? ram_41 : _GEN_6343; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6345 = 10'h2a == _T_19 ? ram_42 : _GEN_6344; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6346 = 10'h2b == _T_19 ? ram_43 : _GEN_6345; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6347 = 10'h2c == _T_19 ? ram_44 : _GEN_6346; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6348 = 10'h2d == _T_19 ? ram_45 : _GEN_6347; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6349 = 10'h2e == _T_19 ? ram_46 : _GEN_6348; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6350 = 10'h2f == _T_19 ? ram_47 : _GEN_6349; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6351 = 10'h30 == _T_19 ? ram_48 : _GEN_6350; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6352 = 10'h31 == _T_19 ? ram_49 : _GEN_6351; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6353 = 10'h32 == _T_19 ? ram_50 : _GEN_6352; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6354 = 10'h33 == _T_19 ? ram_51 : _GEN_6353; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6355 = 10'h34 == _T_19 ? ram_52 : _GEN_6354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6356 = 10'h35 == _T_19 ? ram_53 : _GEN_6355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6357 = 10'h36 == _T_19 ? ram_54 : _GEN_6356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6358 = 10'h37 == _T_19 ? ram_55 : _GEN_6357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6359 = 10'h38 == _T_19 ? ram_56 : _GEN_6358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6360 = 10'h39 == _T_19 ? ram_57 : _GEN_6359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6361 = 10'h3a == _T_19 ? ram_58 : _GEN_6360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6362 = 10'h3b == _T_19 ? ram_59 : _GEN_6361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6363 = 10'h3c == _T_19 ? ram_60 : _GEN_6362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6364 = 10'h3d == _T_19 ? ram_61 : _GEN_6363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6365 = 10'h3e == _T_19 ? ram_62 : _GEN_6364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6366 = 10'h3f == _T_19 ? ram_63 : _GEN_6365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6367 = 10'h40 == _T_19 ? ram_64 : _GEN_6366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6368 = 10'h41 == _T_19 ? ram_65 : _GEN_6367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6369 = 10'h42 == _T_19 ? ram_66 : _GEN_6368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6370 = 10'h43 == _T_19 ? ram_67 : _GEN_6369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6371 = 10'h44 == _T_19 ? ram_68 : _GEN_6370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6372 = 10'h45 == _T_19 ? ram_69 : _GEN_6371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6373 = 10'h46 == _T_19 ? ram_70 : _GEN_6372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6374 = 10'h47 == _T_19 ? ram_71 : _GEN_6373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6375 = 10'h48 == _T_19 ? ram_72 : _GEN_6374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6376 = 10'h49 == _T_19 ? ram_73 : _GEN_6375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6377 = 10'h4a == _T_19 ? ram_74 : _GEN_6376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6378 = 10'h4b == _T_19 ? ram_75 : _GEN_6377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6379 = 10'h4c == _T_19 ? ram_76 : _GEN_6378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6380 = 10'h4d == _T_19 ? ram_77 : _GEN_6379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6381 = 10'h4e == _T_19 ? ram_78 : _GEN_6380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6382 = 10'h4f == _T_19 ? ram_79 : _GEN_6381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6383 = 10'h50 == _T_19 ? ram_80 : _GEN_6382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6384 = 10'h51 == _T_19 ? ram_81 : _GEN_6383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6385 = 10'h52 == _T_19 ? ram_82 : _GEN_6384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6386 = 10'h53 == _T_19 ? ram_83 : _GEN_6385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6387 = 10'h54 == _T_19 ? ram_84 : _GEN_6386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6388 = 10'h55 == _T_19 ? ram_85 : _GEN_6387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6389 = 10'h56 == _T_19 ? ram_86 : _GEN_6388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6390 = 10'h57 == _T_19 ? ram_87 : _GEN_6389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6391 = 10'h58 == _T_19 ? ram_88 : _GEN_6390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6392 = 10'h59 == _T_19 ? ram_89 : _GEN_6391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6393 = 10'h5a == _T_19 ? ram_90 : _GEN_6392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6394 = 10'h5b == _T_19 ? ram_91 : _GEN_6393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6395 = 10'h5c == _T_19 ? ram_92 : _GEN_6394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6396 = 10'h5d == _T_19 ? ram_93 : _GEN_6395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6397 = 10'h5e == _T_19 ? ram_94 : _GEN_6396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6398 = 10'h5f == _T_19 ? ram_95 : _GEN_6397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6399 = 10'h60 == _T_19 ? ram_96 : _GEN_6398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6400 = 10'h61 == _T_19 ? ram_97 : _GEN_6399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6401 = 10'h62 == _T_19 ? ram_98 : _GEN_6400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6402 = 10'h63 == _T_19 ? ram_99 : _GEN_6401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6403 = 10'h64 == _T_19 ? ram_100 : _GEN_6402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6404 = 10'h65 == _T_19 ? ram_101 : _GEN_6403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6405 = 10'h66 == _T_19 ? ram_102 : _GEN_6404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6406 = 10'h67 == _T_19 ? ram_103 : _GEN_6405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6407 = 10'h68 == _T_19 ? ram_104 : _GEN_6406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6408 = 10'h69 == _T_19 ? ram_105 : _GEN_6407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6409 = 10'h6a == _T_19 ? ram_106 : _GEN_6408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6410 = 10'h6b == _T_19 ? ram_107 : _GEN_6409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6411 = 10'h6c == _T_19 ? ram_108 : _GEN_6410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6412 = 10'h6d == _T_19 ? ram_109 : _GEN_6411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6413 = 10'h6e == _T_19 ? ram_110 : _GEN_6412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6414 = 10'h6f == _T_19 ? ram_111 : _GEN_6413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6415 = 10'h70 == _T_19 ? ram_112 : _GEN_6414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6416 = 10'h71 == _T_19 ? ram_113 : _GEN_6415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6417 = 10'h72 == _T_19 ? ram_114 : _GEN_6416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6418 = 10'h73 == _T_19 ? ram_115 : _GEN_6417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6419 = 10'h74 == _T_19 ? ram_116 : _GEN_6418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6420 = 10'h75 == _T_19 ? ram_117 : _GEN_6419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6421 = 10'h76 == _T_19 ? ram_118 : _GEN_6420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6422 = 10'h77 == _T_19 ? ram_119 : _GEN_6421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6423 = 10'h78 == _T_19 ? ram_120 : _GEN_6422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6424 = 10'h79 == _T_19 ? ram_121 : _GEN_6423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6425 = 10'h7a == _T_19 ? ram_122 : _GEN_6424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6426 = 10'h7b == _T_19 ? ram_123 : _GEN_6425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6427 = 10'h7c == _T_19 ? ram_124 : _GEN_6426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6428 = 10'h7d == _T_19 ? ram_125 : _GEN_6427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6429 = 10'h7e == _T_19 ? ram_126 : _GEN_6428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6430 = 10'h7f == _T_19 ? ram_127 : _GEN_6429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6431 = 10'h80 == _T_19 ? ram_128 : _GEN_6430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6432 = 10'h81 == _T_19 ? ram_129 : _GEN_6431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6433 = 10'h82 == _T_19 ? ram_130 : _GEN_6432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6434 = 10'h83 == _T_19 ? ram_131 : _GEN_6433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6435 = 10'h84 == _T_19 ? ram_132 : _GEN_6434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6436 = 10'h85 == _T_19 ? ram_133 : _GEN_6435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6437 = 10'h86 == _T_19 ? ram_134 : _GEN_6436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6438 = 10'h87 == _T_19 ? ram_135 : _GEN_6437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6439 = 10'h88 == _T_19 ? ram_136 : _GEN_6438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6440 = 10'h89 == _T_19 ? ram_137 : _GEN_6439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6441 = 10'h8a == _T_19 ? ram_138 : _GEN_6440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6442 = 10'h8b == _T_19 ? ram_139 : _GEN_6441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6443 = 10'h8c == _T_19 ? ram_140 : _GEN_6442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6444 = 10'h8d == _T_19 ? ram_141 : _GEN_6443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6445 = 10'h8e == _T_19 ? ram_142 : _GEN_6444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6446 = 10'h8f == _T_19 ? ram_143 : _GEN_6445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6447 = 10'h90 == _T_19 ? ram_144 : _GEN_6446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6448 = 10'h91 == _T_19 ? ram_145 : _GEN_6447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6449 = 10'h92 == _T_19 ? ram_146 : _GEN_6448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6450 = 10'h93 == _T_19 ? ram_147 : _GEN_6449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6451 = 10'h94 == _T_19 ? ram_148 : _GEN_6450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6452 = 10'h95 == _T_19 ? ram_149 : _GEN_6451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6453 = 10'h96 == _T_19 ? ram_150 : _GEN_6452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6454 = 10'h97 == _T_19 ? ram_151 : _GEN_6453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6455 = 10'h98 == _T_19 ? ram_152 : _GEN_6454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6456 = 10'h99 == _T_19 ? ram_153 : _GEN_6455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6457 = 10'h9a == _T_19 ? ram_154 : _GEN_6456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6458 = 10'h9b == _T_19 ? ram_155 : _GEN_6457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6459 = 10'h9c == _T_19 ? ram_156 : _GEN_6458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6460 = 10'h9d == _T_19 ? ram_157 : _GEN_6459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6461 = 10'h9e == _T_19 ? ram_158 : _GEN_6460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6462 = 10'h9f == _T_19 ? ram_159 : _GEN_6461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6463 = 10'ha0 == _T_19 ? ram_160 : _GEN_6462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6464 = 10'ha1 == _T_19 ? ram_161 : _GEN_6463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6465 = 10'ha2 == _T_19 ? ram_162 : _GEN_6464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6466 = 10'ha3 == _T_19 ? ram_163 : _GEN_6465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6467 = 10'ha4 == _T_19 ? ram_164 : _GEN_6466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6468 = 10'ha5 == _T_19 ? ram_165 : _GEN_6467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6469 = 10'ha6 == _T_19 ? ram_166 : _GEN_6468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6470 = 10'ha7 == _T_19 ? ram_167 : _GEN_6469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6471 = 10'ha8 == _T_19 ? ram_168 : _GEN_6470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6472 = 10'ha9 == _T_19 ? ram_169 : _GEN_6471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6473 = 10'haa == _T_19 ? ram_170 : _GEN_6472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6474 = 10'hab == _T_19 ? ram_171 : _GEN_6473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6475 = 10'hac == _T_19 ? ram_172 : _GEN_6474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6476 = 10'had == _T_19 ? ram_173 : _GEN_6475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6477 = 10'hae == _T_19 ? ram_174 : _GEN_6476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6478 = 10'haf == _T_19 ? ram_175 : _GEN_6477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6479 = 10'hb0 == _T_19 ? ram_176 : _GEN_6478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6480 = 10'hb1 == _T_19 ? ram_177 : _GEN_6479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6481 = 10'hb2 == _T_19 ? ram_178 : _GEN_6480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6482 = 10'hb3 == _T_19 ? ram_179 : _GEN_6481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6483 = 10'hb4 == _T_19 ? ram_180 : _GEN_6482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6484 = 10'hb5 == _T_19 ? ram_181 : _GEN_6483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6485 = 10'hb6 == _T_19 ? ram_182 : _GEN_6484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6486 = 10'hb7 == _T_19 ? ram_183 : _GEN_6485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6487 = 10'hb8 == _T_19 ? ram_184 : _GEN_6486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6488 = 10'hb9 == _T_19 ? ram_185 : _GEN_6487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6489 = 10'hba == _T_19 ? ram_186 : _GEN_6488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6490 = 10'hbb == _T_19 ? ram_187 : _GEN_6489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6491 = 10'hbc == _T_19 ? ram_188 : _GEN_6490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6492 = 10'hbd == _T_19 ? ram_189 : _GEN_6491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6493 = 10'hbe == _T_19 ? ram_190 : _GEN_6492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6494 = 10'hbf == _T_19 ? ram_191 : _GEN_6493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6495 = 10'hc0 == _T_19 ? ram_192 : _GEN_6494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6496 = 10'hc1 == _T_19 ? ram_193 : _GEN_6495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6497 = 10'hc2 == _T_19 ? ram_194 : _GEN_6496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6498 = 10'hc3 == _T_19 ? ram_195 : _GEN_6497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6499 = 10'hc4 == _T_19 ? ram_196 : _GEN_6498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6500 = 10'hc5 == _T_19 ? ram_197 : _GEN_6499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6501 = 10'hc6 == _T_19 ? ram_198 : _GEN_6500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6502 = 10'hc7 == _T_19 ? ram_199 : _GEN_6501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6503 = 10'hc8 == _T_19 ? ram_200 : _GEN_6502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6504 = 10'hc9 == _T_19 ? ram_201 : _GEN_6503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6505 = 10'hca == _T_19 ? ram_202 : _GEN_6504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6506 = 10'hcb == _T_19 ? ram_203 : _GEN_6505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6507 = 10'hcc == _T_19 ? ram_204 : _GEN_6506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6508 = 10'hcd == _T_19 ? ram_205 : _GEN_6507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6509 = 10'hce == _T_19 ? ram_206 : _GEN_6508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6510 = 10'hcf == _T_19 ? ram_207 : _GEN_6509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6511 = 10'hd0 == _T_19 ? ram_208 : _GEN_6510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6512 = 10'hd1 == _T_19 ? ram_209 : _GEN_6511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6513 = 10'hd2 == _T_19 ? ram_210 : _GEN_6512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6514 = 10'hd3 == _T_19 ? ram_211 : _GEN_6513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6515 = 10'hd4 == _T_19 ? ram_212 : _GEN_6514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6516 = 10'hd5 == _T_19 ? ram_213 : _GEN_6515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6517 = 10'hd6 == _T_19 ? ram_214 : _GEN_6516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6518 = 10'hd7 == _T_19 ? ram_215 : _GEN_6517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6519 = 10'hd8 == _T_19 ? ram_216 : _GEN_6518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6520 = 10'hd9 == _T_19 ? ram_217 : _GEN_6519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6521 = 10'hda == _T_19 ? ram_218 : _GEN_6520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6522 = 10'hdb == _T_19 ? ram_219 : _GEN_6521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6523 = 10'hdc == _T_19 ? ram_220 : _GEN_6522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6524 = 10'hdd == _T_19 ? ram_221 : _GEN_6523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6525 = 10'hde == _T_19 ? ram_222 : _GEN_6524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6526 = 10'hdf == _T_19 ? ram_223 : _GEN_6525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6527 = 10'he0 == _T_19 ? ram_224 : _GEN_6526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6528 = 10'he1 == _T_19 ? ram_225 : _GEN_6527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6529 = 10'he2 == _T_19 ? ram_226 : _GEN_6528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6530 = 10'he3 == _T_19 ? ram_227 : _GEN_6529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6531 = 10'he4 == _T_19 ? ram_228 : _GEN_6530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6532 = 10'he5 == _T_19 ? ram_229 : _GEN_6531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6533 = 10'he6 == _T_19 ? ram_230 : _GEN_6532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6534 = 10'he7 == _T_19 ? ram_231 : _GEN_6533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6535 = 10'he8 == _T_19 ? ram_232 : _GEN_6534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6536 = 10'he9 == _T_19 ? ram_233 : _GEN_6535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6537 = 10'hea == _T_19 ? ram_234 : _GEN_6536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6538 = 10'heb == _T_19 ? ram_235 : _GEN_6537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6539 = 10'hec == _T_19 ? ram_236 : _GEN_6538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6540 = 10'hed == _T_19 ? ram_237 : _GEN_6539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6541 = 10'hee == _T_19 ? ram_238 : _GEN_6540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6542 = 10'hef == _T_19 ? ram_239 : _GEN_6541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6543 = 10'hf0 == _T_19 ? ram_240 : _GEN_6542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6544 = 10'hf1 == _T_19 ? ram_241 : _GEN_6543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6545 = 10'hf2 == _T_19 ? ram_242 : _GEN_6544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6546 = 10'hf3 == _T_19 ? ram_243 : _GEN_6545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6547 = 10'hf4 == _T_19 ? ram_244 : _GEN_6546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6548 = 10'hf5 == _T_19 ? ram_245 : _GEN_6547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6549 = 10'hf6 == _T_19 ? ram_246 : _GEN_6548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6550 = 10'hf7 == _T_19 ? ram_247 : _GEN_6549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6551 = 10'hf8 == _T_19 ? ram_248 : _GEN_6550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6552 = 10'hf9 == _T_19 ? ram_249 : _GEN_6551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6553 = 10'hfa == _T_19 ? ram_250 : _GEN_6552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6554 = 10'hfb == _T_19 ? ram_251 : _GEN_6553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6555 = 10'hfc == _T_19 ? ram_252 : _GEN_6554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6556 = 10'hfd == _T_19 ? ram_253 : _GEN_6555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6557 = 10'hfe == _T_19 ? ram_254 : _GEN_6556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6558 = 10'hff == _T_19 ? ram_255 : _GEN_6557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6559 = 10'h100 == _T_19 ? ram_256 : _GEN_6558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6560 = 10'h101 == _T_19 ? ram_257 : _GEN_6559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6561 = 10'h102 == _T_19 ? ram_258 : _GEN_6560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6562 = 10'h103 == _T_19 ? ram_259 : _GEN_6561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6563 = 10'h104 == _T_19 ? ram_260 : _GEN_6562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6564 = 10'h105 == _T_19 ? ram_261 : _GEN_6563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6565 = 10'h106 == _T_19 ? ram_262 : _GEN_6564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6566 = 10'h107 == _T_19 ? ram_263 : _GEN_6565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6567 = 10'h108 == _T_19 ? ram_264 : _GEN_6566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6568 = 10'h109 == _T_19 ? ram_265 : _GEN_6567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6569 = 10'h10a == _T_19 ? ram_266 : _GEN_6568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6570 = 10'h10b == _T_19 ? ram_267 : _GEN_6569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6571 = 10'h10c == _T_19 ? ram_268 : _GEN_6570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6572 = 10'h10d == _T_19 ? ram_269 : _GEN_6571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6573 = 10'h10e == _T_19 ? ram_270 : _GEN_6572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6574 = 10'h10f == _T_19 ? ram_271 : _GEN_6573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6575 = 10'h110 == _T_19 ? ram_272 : _GEN_6574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6576 = 10'h111 == _T_19 ? ram_273 : _GEN_6575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6577 = 10'h112 == _T_19 ? ram_274 : _GEN_6576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6578 = 10'h113 == _T_19 ? ram_275 : _GEN_6577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6579 = 10'h114 == _T_19 ? ram_276 : _GEN_6578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6580 = 10'h115 == _T_19 ? ram_277 : _GEN_6579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6581 = 10'h116 == _T_19 ? ram_278 : _GEN_6580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6582 = 10'h117 == _T_19 ? ram_279 : _GEN_6581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6583 = 10'h118 == _T_19 ? ram_280 : _GEN_6582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6584 = 10'h119 == _T_19 ? ram_281 : _GEN_6583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6585 = 10'h11a == _T_19 ? ram_282 : _GEN_6584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6586 = 10'h11b == _T_19 ? ram_283 : _GEN_6585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6587 = 10'h11c == _T_19 ? ram_284 : _GEN_6586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6588 = 10'h11d == _T_19 ? ram_285 : _GEN_6587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6589 = 10'h11e == _T_19 ? ram_286 : _GEN_6588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6590 = 10'h11f == _T_19 ? ram_287 : _GEN_6589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6591 = 10'h120 == _T_19 ? ram_288 : _GEN_6590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6592 = 10'h121 == _T_19 ? ram_289 : _GEN_6591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6593 = 10'h122 == _T_19 ? ram_290 : _GEN_6592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6594 = 10'h123 == _T_19 ? ram_291 : _GEN_6593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6595 = 10'h124 == _T_19 ? ram_292 : _GEN_6594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6596 = 10'h125 == _T_19 ? ram_293 : _GEN_6595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6597 = 10'h126 == _T_19 ? ram_294 : _GEN_6596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6598 = 10'h127 == _T_19 ? ram_295 : _GEN_6597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6599 = 10'h128 == _T_19 ? ram_296 : _GEN_6598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6600 = 10'h129 == _T_19 ? ram_297 : _GEN_6599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6601 = 10'h12a == _T_19 ? ram_298 : _GEN_6600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6602 = 10'h12b == _T_19 ? ram_299 : _GEN_6601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6603 = 10'h12c == _T_19 ? ram_300 : _GEN_6602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6604 = 10'h12d == _T_19 ? ram_301 : _GEN_6603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6605 = 10'h12e == _T_19 ? ram_302 : _GEN_6604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6606 = 10'h12f == _T_19 ? ram_303 : _GEN_6605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6607 = 10'h130 == _T_19 ? ram_304 : _GEN_6606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6608 = 10'h131 == _T_19 ? ram_305 : _GEN_6607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6609 = 10'h132 == _T_19 ? ram_306 : _GEN_6608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6610 = 10'h133 == _T_19 ? ram_307 : _GEN_6609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6611 = 10'h134 == _T_19 ? ram_308 : _GEN_6610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6612 = 10'h135 == _T_19 ? ram_309 : _GEN_6611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6613 = 10'h136 == _T_19 ? ram_310 : _GEN_6612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6614 = 10'h137 == _T_19 ? ram_311 : _GEN_6613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6615 = 10'h138 == _T_19 ? ram_312 : _GEN_6614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6616 = 10'h139 == _T_19 ? ram_313 : _GEN_6615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6617 = 10'h13a == _T_19 ? ram_314 : _GEN_6616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6618 = 10'h13b == _T_19 ? ram_315 : _GEN_6617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6619 = 10'h13c == _T_19 ? ram_316 : _GEN_6618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6620 = 10'h13d == _T_19 ? ram_317 : _GEN_6619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6621 = 10'h13e == _T_19 ? ram_318 : _GEN_6620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6622 = 10'h13f == _T_19 ? ram_319 : _GEN_6621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6623 = 10'h140 == _T_19 ? ram_320 : _GEN_6622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6624 = 10'h141 == _T_19 ? ram_321 : _GEN_6623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6625 = 10'h142 == _T_19 ? ram_322 : _GEN_6624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6626 = 10'h143 == _T_19 ? ram_323 : _GEN_6625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6627 = 10'h144 == _T_19 ? ram_324 : _GEN_6626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6628 = 10'h145 == _T_19 ? ram_325 : _GEN_6627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6629 = 10'h146 == _T_19 ? ram_326 : _GEN_6628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6630 = 10'h147 == _T_19 ? ram_327 : _GEN_6629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6631 = 10'h148 == _T_19 ? ram_328 : _GEN_6630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6632 = 10'h149 == _T_19 ? ram_329 : _GEN_6631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6633 = 10'h14a == _T_19 ? ram_330 : _GEN_6632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6634 = 10'h14b == _T_19 ? ram_331 : _GEN_6633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6635 = 10'h14c == _T_19 ? ram_332 : _GEN_6634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6636 = 10'h14d == _T_19 ? ram_333 : _GEN_6635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6637 = 10'h14e == _T_19 ? ram_334 : _GEN_6636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6638 = 10'h14f == _T_19 ? ram_335 : _GEN_6637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6639 = 10'h150 == _T_19 ? ram_336 : _GEN_6638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6640 = 10'h151 == _T_19 ? ram_337 : _GEN_6639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6641 = 10'h152 == _T_19 ? ram_338 : _GEN_6640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6642 = 10'h153 == _T_19 ? ram_339 : _GEN_6641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6643 = 10'h154 == _T_19 ? ram_340 : _GEN_6642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6644 = 10'h155 == _T_19 ? ram_341 : _GEN_6643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6645 = 10'h156 == _T_19 ? ram_342 : _GEN_6644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6646 = 10'h157 == _T_19 ? ram_343 : _GEN_6645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6647 = 10'h158 == _T_19 ? ram_344 : _GEN_6646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6648 = 10'h159 == _T_19 ? ram_345 : _GEN_6647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6649 = 10'h15a == _T_19 ? ram_346 : _GEN_6648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6650 = 10'h15b == _T_19 ? ram_347 : _GEN_6649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6651 = 10'h15c == _T_19 ? ram_348 : _GEN_6650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6652 = 10'h15d == _T_19 ? ram_349 : _GEN_6651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6653 = 10'h15e == _T_19 ? ram_350 : _GEN_6652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6654 = 10'h15f == _T_19 ? ram_351 : _GEN_6653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6655 = 10'h160 == _T_19 ? ram_352 : _GEN_6654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6656 = 10'h161 == _T_19 ? ram_353 : _GEN_6655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6657 = 10'h162 == _T_19 ? ram_354 : _GEN_6656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6658 = 10'h163 == _T_19 ? ram_355 : _GEN_6657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6659 = 10'h164 == _T_19 ? ram_356 : _GEN_6658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6660 = 10'h165 == _T_19 ? ram_357 : _GEN_6659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6661 = 10'h166 == _T_19 ? ram_358 : _GEN_6660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6662 = 10'h167 == _T_19 ? ram_359 : _GEN_6661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6663 = 10'h168 == _T_19 ? ram_360 : _GEN_6662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6664 = 10'h169 == _T_19 ? ram_361 : _GEN_6663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6665 = 10'h16a == _T_19 ? ram_362 : _GEN_6664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6666 = 10'h16b == _T_19 ? ram_363 : _GEN_6665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6667 = 10'h16c == _T_19 ? ram_364 : _GEN_6666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6668 = 10'h16d == _T_19 ? ram_365 : _GEN_6667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6669 = 10'h16e == _T_19 ? ram_366 : _GEN_6668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6670 = 10'h16f == _T_19 ? ram_367 : _GEN_6669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6671 = 10'h170 == _T_19 ? ram_368 : _GEN_6670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6672 = 10'h171 == _T_19 ? ram_369 : _GEN_6671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6673 = 10'h172 == _T_19 ? ram_370 : _GEN_6672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6674 = 10'h173 == _T_19 ? ram_371 : _GEN_6673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6675 = 10'h174 == _T_19 ? ram_372 : _GEN_6674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6676 = 10'h175 == _T_19 ? ram_373 : _GEN_6675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6677 = 10'h176 == _T_19 ? ram_374 : _GEN_6676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6678 = 10'h177 == _T_19 ? ram_375 : _GEN_6677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6679 = 10'h178 == _T_19 ? ram_376 : _GEN_6678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6680 = 10'h179 == _T_19 ? ram_377 : _GEN_6679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6681 = 10'h17a == _T_19 ? ram_378 : _GEN_6680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6682 = 10'h17b == _T_19 ? ram_379 : _GEN_6681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6683 = 10'h17c == _T_19 ? ram_380 : _GEN_6682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6684 = 10'h17d == _T_19 ? ram_381 : _GEN_6683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6685 = 10'h17e == _T_19 ? ram_382 : _GEN_6684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6686 = 10'h17f == _T_19 ? ram_383 : _GEN_6685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6687 = 10'h180 == _T_19 ? ram_384 : _GEN_6686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6688 = 10'h181 == _T_19 ? ram_385 : _GEN_6687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6689 = 10'h182 == _T_19 ? ram_386 : _GEN_6688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6690 = 10'h183 == _T_19 ? ram_387 : _GEN_6689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6691 = 10'h184 == _T_19 ? ram_388 : _GEN_6690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6692 = 10'h185 == _T_19 ? ram_389 : _GEN_6691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6693 = 10'h186 == _T_19 ? ram_390 : _GEN_6692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6694 = 10'h187 == _T_19 ? ram_391 : _GEN_6693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6695 = 10'h188 == _T_19 ? ram_392 : _GEN_6694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6696 = 10'h189 == _T_19 ? ram_393 : _GEN_6695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6697 = 10'h18a == _T_19 ? ram_394 : _GEN_6696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6698 = 10'h18b == _T_19 ? ram_395 : _GEN_6697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6699 = 10'h18c == _T_19 ? ram_396 : _GEN_6698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6700 = 10'h18d == _T_19 ? ram_397 : _GEN_6699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6701 = 10'h18e == _T_19 ? ram_398 : _GEN_6700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6702 = 10'h18f == _T_19 ? ram_399 : _GEN_6701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6703 = 10'h190 == _T_19 ? ram_400 : _GEN_6702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6704 = 10'h191 == _T_19 ? ram_401 : _GEN_6703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6705 = 10'h192 == _T_19 ? ram_402 : _GEN_6704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6706 = 10'h193 == _T_19 ? ram_403 : _GEN_6705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6707 = 10'h194 == _T_19 ? ram_404 : _GEN_6706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6708 = 10'h195 == _T_19 ? ram_405 : _GEN_6707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6709 = 10'h196 == _T_19 ? ram_406 : _GEN_6708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6710 = 10'h197 == _T_19 ? ram_407 : _GEN_6709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6711 = 10'h198 == _T_19 ? ram_408 : _GEN_6710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6712 = 10'h199 == _T_19 ? ram_409 : _GEN_6711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6713 = 10'h19a == _T_19 ? ram_410 : _GEN_6712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6714 = 10'h19b == _T_19 ? ram_411 : _GEN_6713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6715 = 10'h19c == _T_19 ? ram_412 : _GEN_6714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6716 = 10'h19d == _T_19 ? ram_413 : _GEN_6715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6717 = 10'h19e == _T_19 ? ram_414 : _GEN_6716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6718 = 10'h19f == _T_19 ? ram_415 : _GEN_6717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6719 = 10'h1a0 == _T_19 ? ram_416 : _GEN_6718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6720 = 10'h1a1 == _T_19 ? ram_417 : _GEN_6719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6721 = 10'h1a2 == _T_19 ? ram_418 : _GEN_6720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6722 = 10'h1a3 == _T_19 ? ram_419 : _GEN_6721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6723 = 10'h1a4 == _T_19 ? ram_420 : _GEN_6722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6724 = 10'h1a5 == _T_19 ? ram_421 : _GEN_6723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6725 = 10'h1a6 == _T_19 ? ram_422 : _GEN_6724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6726 = 10'h1a7 == _T_19 ? ram_423 : _GEN_6725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6727 = 10'h1a8 == _T_19 ? ram_424 : _GEN_6726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6728 = 10'h1a9 == _T_19 ? ram_425 : _GEN_6727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6729 = 10'h1aa == _T_19 ? ram_426 : _GEN_6728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6730 = 10'h1ab == _T_19 ? ram_427 : _GEN_6729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6731 = 10'h1ac == _T_19 ? ram_428 : _GEN_6730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6732 = 10'h1ad == _T_19 ? ram_429 : _GEN_6731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6733 = 10'h1ae == _T_19 ? ram_430 : _GEN_6732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6734 = 10'h1af == _T_19 ? ram_431 : _GEN_6733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6735 = 10'h1b0 == _T_19 ? ram_432 : _GEN_6734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6736 = 10'h1b1 == _T_19 ? ram_433 : _GEN_6735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6737 = 10'h1b2 == _T_19 ? ram_434 : _GEN_6736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6738 = 10'h1b3 == _T_19 ? ram_435 : _GEN_6737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6739 = 10'h1b4 == _T_19 ? ram_436 : _GEN_6738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6740 = 10'h1b5 == _T_19 ? ram_437 : _GEN_6739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6741 = 10'h1b6 == _T_19 ? ram_438 : _GEN_6740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6742 = 10'h1b7 == _T_19 ? ram_439 : _GEN_6741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6743 = 10'h1b8 == _T_19 ? ram_440 : _GEN_6742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6744 = 10'h1b9 == _T_19 ? ram_441 : _GEN_6743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6745 = 10'h1ba == _T_19 ? ram_442 : _GEN_6744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6746 = 10'h1bb == _T_19 ? ram_443 : _GEN_6745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6747 = 10'h1bc == _T_19 ? ram_444 : _GEN_6746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6748 = 10'h1bd == _T_19 ? ram_445 : _GEN_6747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6749 = 10'h1be == _T_19 ? ram_446 : _GEN_6748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6750 = 10'h1bf == _T_19 ? ram_447 : _GEN_6749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6751 = 10'h1c0 == _T_19 ? ram_448 : _GEN_6750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6752 = 10'h1c1 == _T_19 ? ram_449 : _GEN_6751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6753 = 10'h1c2 == _T_19 ? ram_450 : _GEN_6752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6754 = 10'h1c3 == _T_19 ? ram_451 : _GEN_6753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6755 = 10'h1c4 == _T_19 ? ram_452 : _GEN_6754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6756 = 10'h1c5 == _T_19 ? ram_453 : _GEN_6755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6757 = 10'h1c6 == _T_19 ? ram_454 : _GEN_6756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6758 = 10'h1c7 == _T_19 ? ram_455 : _GEN_6757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6759 = 10'h1c8 == _T_19 ? ram_456 : _GEN_6758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6760 = 10'h1c9 == _T_19 ? ram_457 : _GEN_6759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6761 = 10'h1ca == _T_19 ? ram_458 : _GEN_6760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6762 = 10'h1cb == _T_19 ? ram_459 : _GEN_6761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6763 = 10'h1cc == _T_19 ? ram_460 : _GEN_6762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6764 = 10'h1cd == _T_19 ? ram_461 : _GEN_6763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6765 = 10'h1ce == _T_19 ? ram_462 : _GEN_6764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6766 = 10'h1cf == _T_19 ? ram_463 : _GEN_6765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6767 = 10'h1d0 == _T_19 ? ram_464 : _GEN_6766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6768 = 10'h1d1 == _T_19 ? ram_465 : _GEN_6767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6769 = 10'h1d2 == _T_19 ? ram_466 : _GEN_6768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6770 = 10'h1d3 == _T_19 ? ram_467 : _GEN_6769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6771 = 10'h1d4 == _T_19 ? ram_468 : _GEN_6770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6772 = 10'h1d5 == _T_19 ? ram_469 : _GEN_6771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6773 = 10'h1d6 == _T_19 ? ram_470 : _GEN_6772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6774 = 10'h1d7 == _T_19 ? ram_471 : _GEN_6773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6775 = 10'h1d8 == _T_19 ? ram_472 : _GEN_6774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6776 = 10'h1d9 == _T_19 ? ram_473 : _GEN_6775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6777 = 10'h1da == _T_19 ? ram_474 : _GEN_6776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6778 = 10'h1db == _T_19 ? ram_475 : _GEN_6777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6779 = 10'h1dc == _T_19 ? ram_476 : _GEN_6778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6780 = 10'h1dd == _T_19 ? ram_477 : _GEN_6779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6781 = 10'h1de == _T_19 ? ram_478 : _GEN_6780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6782 = 10'h1df == _T_19 ? ram_479 : _GEN_6781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6783 = 10'h1e0 == _T_19 ? ram_480 : _GEN_6782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6784 = 10'h1e1 == _T_19 ? ram_481 : _GEN_6783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6785 = 10'h1e2 == _T_19 ? ram_482 : _GEN_6784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6786 = 10'h1e3 == _T_19 ? ram_483 : _GEN_6785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6787 = 10'h1e4 == _T_19 ? ram_484 : _GEN_6786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6788 = 10'h1e5 == _T_19 ? ram_485 : _GEN_6787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6789 = 10'h1e6 == _T_19 ? ram_486 : _GEN_6788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6790 = 10'h1e7 == _T_19 ? ram_487 : _GEN_6789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6791 = 10'h1e8 == _T_19 ? ram_488 : _GEN_6790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6792 = 10'h1e9 == _T_19 ? ram_489 : _GEN_6791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6793 = 10'h1ea == _T_19 ? ram_490 : _GEN_6792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6794 = 10'h1eb == _T_19 ? ram_491 : _GEN_6793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6795 = 10'h1ec == _T_19 ? ram_492 : _GEN_6794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6796 = 10'h1ed == _T_19 ? ram_493 : _GEN_6795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6797 = 10'h1ee == _T_19 ? ram_494 : _GEN_6796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6798 = 10'h1ef == _T_19 ? ram_495 : _GEN_6797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6799 = 10'h1f0 == _T_19 ? ram_496 : _GEN_6798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6800 = 10'h1f1 == _T_19 ? ram_497 : _GEN_6799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6801 = 10'h1f2 == _T_19 ? ram_498 : _GEN_6800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6802 = 10'h1f3 == _T_19 ? ram_499 : _GEN_6801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6803 = 10'h1f4 == _T_19 ? ram_500 : _GEN_6802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6804 = 10'h1f5 == _T_19 ? ram_501 : _GEN_6803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6805 = 10'h1f6 == _T_19 ? ram_502 : _GEN_6804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6806 = 10'h1f7 == _T_19 ? ram_503 : _GEN_6805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6807 = 10'h1f8 == _T_19 ? ram_504 : _GEN_6806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6808 = 10'h1f9 == _T_19 ? ram_505 : _GEN_6807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6809 = 10'h1fa == _T_19 ? ram_506 : _GEN_6808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6810 = 10'h1fb == _T_19 ? ram_507 : _GEN_6809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6811 = 10'h1fc == _T_19 ? ram_508 : _GEN_6810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6812 = 10'h1fd == _T_19 ? ram_509 : _GEN_6811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6813 = 10'h1fe == _T_19 ? ram_510 : _GEN_6812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6814 = 10'h1ff == _T_19 ? ram_511 : _GEN_6813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6815 = 10'h200 == _T_19 ? ram_512 : _GEN_6814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6816 = 10'h201 == _T_19 ? ram_513 : _GEN_6815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6817 = 10'h202 == _T_19 ? ram_514 : _GEN_6816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6818 = 10'h203 == _T_19 ? ram_515 : _GEN_6817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6819 = 10'h204 == _T_19 ? ram_516 : _GEN_6818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6820 = 10'h205 == _T_19 ? ram_517 : _GEN_6819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6821 = 10'h206 == _T_19 ? ram_518 : _GEN_6820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6822 = 10'h207 == _T_19 ? ram_519 : _GEN_6821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6823 = 10'h208 == _T_19 ? ram_520 : _GEN_6822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6824 = 10'h209 == _T_19 ? ram_521 : _GEN_6823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6825 = 10'h20a == _T_19 ? ram_522 : _GEN_6824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6826 = 10'h20b == _T_19 ? ram_523 : _GEN_6825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_6827 = 10'h20c == _T_19 ? ram_524 : _GEN_6826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19073 = {{8190'd0}, _GEN_6827}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_181 = _GEN_19073 ^ _ram_T_180; // @[vga.scala 64:41]
  wire [287:0] _GEN_6828 = 10'h0 == _T_19 ? _ram_T_181[287:0] : _GEN_5778; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6829 = 10'h1 == _T_19 ? _ram_T_181[287:0] : _GEN_5779; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6830 = 10'h2 == _T_19 ? _ram_T_181[287:0] : _GEN_5780; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6831 = 10'h3 == _T_19 ? _ram_T_181[287:0] : _GEN_5781; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6832 = 10'h4 == _T_19 ? _ram_T_181[287:0] : _GEN_5782; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6833 = 10'h5 == _T_19 ? _ram_T_181[287:0] : _GEN_5783; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6834 = 10'h6 == _T_19 ? _ram_T_181[287:0] : _GEN_5784; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6835 = 10'h7 == _T_19 ? _ram_T_181[287:0] : _GEN_5785; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6836 = 10'h8 == _T_19 ? _ram_T_181[287:0] : _GEN_5786; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6837 = 10'h9 == _T_19 ? _ram_T_181[287:0] : _GEN_5787; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6838 = 10'ha == _T_19 ? _ram_T_181[287:0] : _GEN_5788; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6839 = 10'hb == _T_19 ? _ram_T_181[287:0] : _GEN_5789; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6840 = 10'hc == _T_19 ? _ram_T_181[287:0] : _GEN_5790; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6841 = 10'hd == _T_19 ? _ram_T_181[287:0] : _GEN_5791; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6842 = 10'he == _T_19 ? _ram_T_181[287:0] : _GEN_5792; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6843 = 10'hf == _T_19 ? _ram_T_181[287:0] : _GEN_5793; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6844 = 10'h10 == _T_19 ? _ram_T_181[287:0] : _GEN_5794; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6845 = 10'h11 == _T_19 ? _ram_T_181[287:0] : _GEN_5795; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6846 = 10'h12 == _T_19 ? _ram_T_181[287:0] : _GEN_5796; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6847 = 10'h13 == _T_19 ? _ram_T_181[287:0] : _GEN_5797; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6848 = 10'h14 == _T_19 ? _ram_T_181[287:0] : _GEN_5798; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6849 = 10'h15 == _T_19 ? _ram_T_181[287:0] : _GEN_5799; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6850 = 10'h16 == _T_19 ? _ram_T_181[287:0] : _GEN_5800; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6851 = 10'h17 == _T_19 ? _ram_T_181[287:0] : _GEN_5801; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6852 = 10'h18 == _T_19 ? _ram_T_181[287:0] : _GEN_5802; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6853 = 10'h19 == _T_19 ? _ram_T_181[287:0] : _GEN_5803; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6854 = 10'h1a == _T_19 ? _ram_T_181[287:0] : _GEN_5804; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6855 = 10'h1b == _T_19 ? _ram_T_181[287:0] : _GEN_5805; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6856 = 10'h1c == _T_19 ? _ram_T_181[287:0] : _GEN_5806; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6857 = 10'h1d == _T_19 ? _ram_T_181[287:0] : _GEN_5807; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6858 = 10'h1e == _T_19 ? _ram_T_181[287:0] : _GEN_5808; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6859 = 10'h1f == _T_19 ? _ram_T_181[287:0] : _GEN_5809; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6860 = 10'h20 == _T_19 ? _ram_T_181[287:0] : _GEN_5810; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6861 = 10'h21 == _T_19 ? _ram_T_181[287:0] : _GEN_5811; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6862 = 10'h22 == _T_19 ? _ram_T_181[287:0] : _GEN_5812; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6863 = 10'h23 == _T_19 ? _ram_T_181[287:0] : _GEN_5813; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6864 = 10'h24 == _T_19 ? _ram_T_181[287:0] : _GEN_5814; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6865 = 10'h25 == _T_19 ? _ram_T_181[287:0] : _GEN_5815; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6866 = 10'h26 == _T_19 ? _ram_T_181[287:0] : _GEN_5816; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6867 = 10'h27 == _T_19 ? _ram_T_181[287:0] : _GEN_5817; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6868 = 10'h28 == _T_19 ? _ram_T_181[287:0] : _GEN_5818; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6869 = 10'h29 == _T_19 ? _ram_T_181[287:0] : _GEN_5819; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6870 = 10'h2a == _T_19 ? _ram_T_181[287:0] : _GEN_5820; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6871 = 10'h2b == _T_19 ? _ram_T_181[287:0] : _GEN_5821; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6872 = 10'h2c == _T_19 ? _ram_T_181[287:0] : _GEN_5822; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6873 = 10'h2d == _T_19 ? _ram_T_181[287:0] : _GEN_5823; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6874 = 10'h2e == _T_19 ? _ram_T_181[287:0] : _GEN_5824; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6875 = 10'h2f == _T_19 ? _ram_T_181[287:0] : _GEN_5825; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6876 = 10'h30 == _T_19 ? _ram_T_181[287:0] : _GEN_5826; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6877 = 10'h31 == _T_19 ? _ram_T_181[287:0] : _GEN_5827; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6878 = 10'h32 == _T_19 ? _ram_T_181[287:0] : _GEN_5828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6879 = 10'h33 == _T_19 ? _ram_T_181[287:0] : _GEN_5829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6880 = 10'h34 == _T_19 ? _ram_T_181[287:0] : _GEN_5830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6881 = 10'h35 == _T_19 ? _ram_T_181[287:0] : _GEN_5831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6882 = 10'h36 == _T_19 ? _ram_T_181[287:0] : _GEN_5832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6883 = 10'h37 == _T_19 ? _ram_T_181[287:0] : _GEN_5833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6884 = 10'h38 == _T_19 ? _ram_T_181[287:0] : _GEN_5834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6885 = 10'h39 == _T_19 ? _ram_T_181[287:0] : _GEN_5835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6886 = 10'h3a == _T_19 ? _ram_T_181[287:0] : _GEN_5836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6887 = 10'h3b == _T_19 ? _ram_T_181[287:0] : _GEN_5837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6888 = 10'h3c == _T_19 ? _ram_T_181[287:0] : _GEN_5838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6889 = 10'h3d == _T_19 ? _ram_T_181[287:0] : _GEN_5839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6890 = 10'h3e == _T_19 ? _ram_T_181[287:0] : _GEN_5840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6891 = 10'h3f == _T_19 ? _ram_T_181[287:0] : _GEN_5841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6892 = 10'h40 == _T_19 ? _ram_T_181[287:0] : _GEN_5842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6893 = 10'h41 == _T_19 ? _ram_T_181[287:0] : _GEN_5843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6894 = 10'h42 == _T_19 ? _ram_T_181[287:0] : _GEN_5844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6895 = 10'h43 == _T_19 ? _ram_T_181[287:0] : _GEN_5845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6896 = 10'h44 == _T_19 ? _ram_T_181[287:0] : _GEN_5846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6897 = 10'h45 == _T_19 ? _ram_T_181[287:0] : _GEN_5847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6898 = 10'h46 == _T_19 ? _ram_T_181[287:0] : _GEN_5848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6899 = 10'h47 == _T_19 ? _ram_T_181[287:0] : _GEN_5849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6900 = 10'h48 == _T_19 ? _ram_T_181[287:0] : _GEN_5850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6901 = 10'h49 == _T_19 ? _ram_T_181[287:0] : _GEN_5851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6902 = 10'h4a == _T_19 ? _ram_T_181[287:0] : _GEN_5852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6903 = 10'h4b == _T_19 ? _ram_T_181[287:0] : _GEN_5853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6904 = 10'h4c == _T_19 ? _ram_T_181[287:0] : _GEN_5854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6905 = 10'h4d == _T_19 ? _ram_T_181[287:0] : _GEN_5855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6906 = 10'h4e == _T_19 ? _ram_T_181[287:0] : _GEN_5856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6907 = 10'h4f == _T_19 ? _ram_T_181[287:0] : _GEN_5857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6908 = 10'h50 == _T_19 ? _ram_T_181[287:0] : _GEN_5858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6909 = 10'h51 == _T_19 ? _ram_T_181[287:0] : _GEN_5859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6910 = 10'h52 == _T_19 ? _ram_T_181[287:0] : _GEN_5860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6911 = 10'h53 == _T_19 ? _ram_T_181[287:0] : _GEN_5861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6912 = 10'h54 == _T_19 ? _ram_T_181[287:0] : _GEN_5862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6913 = 10'h55 == _T_19 ? _ram_T_181[287:0] : _GEN_5863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6914 = 10'h56 == _T_19 ? _ram_T_181[287:0] : _GEN_5864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6915 = 10'h57 == _T_19 ? _ram_T_181[287:0] : _GEN_5865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6916 = 10'h58 == _T_19 ? _ram_T_181[287:0] : _GEN_5866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6917 = 10'h59 == _T_19 ? _ram_T_181[287:0] : _GEN_5867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6918 = 10'h5a == _T_19 ? _ram_T_181[287:0] : _GEN_5868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6919 = 10'h5b == _T_19 ? _ram_T_181[287:0] : _GEN_5869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6920 = 10'h5c == _T_19 ? _ram_T_181[287:0] : _GEN_5870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6921 = 10'h5d == _T_19 ? _ram_T_181[287:0] : _GEN_5871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6922 = 10'h5e == _T_19 ? _ram_T_181[287:0] : _GEN_5872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6923 = 10'h5f == _T_19 ? _ram_T_181[287:0] : _GEN_5873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6924 = 10'h60 == _T_19 ? _ram_T_181[287:0] : _GEN_5874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6925 = 10'h61 == _T_19 ? _ram_T_181[287:0] : _GEN_5875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6926 = 10'h62 == _T_19 ? _ram_T_181[287:0] : _GEN_5876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6927 = 10'h63 == _T_19 ? _ram_T_181[287:0] : _GEN_5877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6928 = 10'h64 == _T_19 ? _ram_T_181[287:0] : _GEN_5878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6929 = 10'h65 == _T_19 ? _ram_T_181[287:0] : _GEN_5879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6930 = 10'h66 == _T_19 ? _ram_T_181[287:0] : _GEN_5880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6931 = 10'h67 == _T_19 ? _ram_T_181[287:0] : _GEN_5881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6932 = 10'h68 == _T_19 ? _ram_T_181[287:0] : _GEN_5882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6933 = 10'h69 == _T_19 ? _ram_T_181[287:0] : _GEN_5883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6934 = 10'h6a == _T_19 ? _ram_T_181[287:0] : _GEN_5884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6935 = 10'h6b == _T_19 ? _ram_T_181[287:0] : _GEN_5885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6936 = 10'h6c == _T_19 ? _ram_T_181[287:0] : _GEN_5886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6937 = 10'h6d == _T_19 ? _ram_T_181[287:0] : _GEN_5887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6938 = 10'h6e == _T_19 ? _ram_T_181[287:0] : _GEN_5888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6939 = 10'h6f == _T_19 ? _ram_T_181[287:0] : _GEN_5889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6940 = 10'h70 == _T_19 ? _ram_T_181[287:0] : _GEN_5890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6941 = 10'h71 == _T_19 ? _ram_T_181[287:0] : _GEN_5891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6942 = 10'h72 == _T_19 ? _ram_T_181[287:0] : _GEN_5892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6943 = 10'h73 == _T_19 ? _ram_T_181[287:0] : _GEN_5893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6944 = 10'h74 == _T_19 ? _ram_T_181[287:0] : _GEN_5894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6945 = 10'h75 == _T_19 ? _ram_T_181[287:0] : _GEN_5895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6946 = 10'h76 == _T_19 ? _ram_T_181[287:0] : _GEN_5896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6947 = 10'h77 == _T_19 ? _ram_T_181[287:0] : _GEN_5897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6948 = 10'h78 == _T_19 ? _ram_T_181[287:0] : _GEN_5898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6949 = 10'h79 == _T_19 ? _ram_T_181[287:0] : _GEN_5899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6950 = 10'h7a == _T_19 ? _ram_T_181[287:0] : _GEN_5900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6951 = 10'h7b == _T_19 ? _ram_T_181[287:0] : _GEN_5901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6952 = 10'h7c == _T_19 ? _ram_T_181[287:0] : _GEN_5902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6953 = 10'h7d == _T_19 ? _ram_T_181[287:0] : _GEN_5903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6954 = 10'h7e == _T_19 ? _ram_T_181[287:0] : _GEN_5904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6955 = 10'h7f == _T_19 ? _ram_T_181[287:0] : _GEN_5905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6956 = 10'h80 == _T_19 ? _ram_T_181[287:0] : _GEN_5906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6957 = 10'h81 == _T_19 ? _ram_T_181[287:0] : _GEN_5907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6958 = 10'h82 == _T_19 ? _ram_T_181[287:0] : _GEN_5908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6959 = 10'h83 == _T_19 ? _ram_T_181[287:0] : _GEN_5909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6960 = 10'h84 == _T_19 ? _ram_T_181[287:0] : _GEN_5910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6961 = 10'h85 == _T_19 ? _ram_T_181[287:0] : _GEN_5911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6962 = 10'h86 == _T_19 ? _ram_T_181[287:0] : _GEN_5912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6963 = 10'h87 == _T_19 ? _ram_T_181[287:0] : _GEN_5913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6964 = 10'h88 == _T_19 ? _ram_T_181[287:0] : _GEN_5914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6965 = 10'h89 == _T_19 ? _ram_T_181[287:0] : _GEN_5915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6966 = 10'h8a == _T_19 ? _ram_T_181[287:0] : _GEN_5916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6967 = 10'h8b == _T_19 ? _ram_T_181[287:0] : _GEN_5917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6968 = 10'h8c == _T_19 ? _ram_T_181[287:0] : _GEN_5918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6969 = 10'h8d == _T_19 ? _ram_T_181[287:0] : _GEN_5919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6970 = 10'h8e == _T_19 ? _ram_T_181[287:0] : _GEN_5920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6971 = 10'h8f == _T_19 ? _ram_T_181[287:0] : _GEN_5921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6972 = 10'h90 == _T_19 ? _ram_T_181[287:0] : _GEN_5922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6973 = 10'h91 == _T_19 ? _ram_T_181[287:0] : _GEN_5923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6974 = 10'h92 == _T_19 ? _ram_T_181[287:0] : _GEN_5924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6975 = 10'h93 == _T_19 ? _ram_T_181[287:0] : _GEN_5925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6976 = 10'h94 == _T_19 ? _ram_T_181[287:0] : _GEN_5926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6977 = 10'h95 == _T_19 ? _ram_T_181[287:0] : _GEN_5927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6978 = 10'h96 == _T_19 ? _ram_T_181[287:0] : _GEN_5928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6979 = 10'h97 == _T_19 ? _ram_T_181[287:0] : _GEN_5929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6980 = 10'h98 == _T_19 ? _ram_T_181[287:0] : _GEN_5930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6981 = 10'h99 == _T_19 ? _ram_T_181[287:0] : _GEN_5931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6982 = 10'h9a == _T_19 ? _ram_T_181[287:0] : _GEN_5932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6983 = 10'h9b == _T_19 ? _ram_T_181[287:0] : _GEN_5933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6984 = 10'h9c == _T_19 ? _ram_T_181[287:0] : _GEN_5934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6985 = 10'h9d == _T_19 ? _ram_T_181[287:0] : _GEN_5935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6986 = 10'h9e == _T_19 ? _ram_T_181[287:0] : _GEN_5936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6987 = 10'h9f == _T_19 ? _ram_T_181[287:0] : _GEN_5937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6988 = 10'ha0 == _T_19 ? _ram_T_181[287:0] : _GEN_5938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6989 = 10'ha1 == _T_19 ? _ram_T_181[287:0] : _GEN_5939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6990 = 10'ha2 == _T_19 ? _ram_T_181[287:0] : _GEN_5940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6991 = 10'ha3 == _T_19 ? _ram_T_181[287:0] : _GEN_5941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6992 = 10'ha4 == _T_19 ? _ram_T_181[287:0] : _GEN_5942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6993 = 10'ha5 == _T_19 ? _ram_T_181[287:0] : _GEN_5943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6994 = 10'ha6 == _T_19 ? _ram_T_181[287:0] : _GEN_5944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6995 = 10'ha7 == _T_19 ? _ram_T_181[287:0] : _GEN_5945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6996 = 10'ha8 == _T_19 ? _ram_T_181[287:0] : _GEN_5946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6997 = 10'ha9 == _T_19 ? _ram_T_181[287:0] : _GEN_5947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6998 = 10'haa == _T_19 ? _ram_T_181[287:0] : _GEN_5948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_6999 = 10'hab == _T_19 ? _ram_T_181[287:0] : _GEN_5949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7000 = 10'hac == _T_19 ? _ram_T_181[287:0] : _GEN_5950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7001 = 10'had == _T_19 ? _ram_T_181[287:0] : _GEN_5951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7002 = 10'hae == _T_19 ? _ram_T_181[287:0] : _GEN_5952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7003 = 10'haf == _T_19 ? _ram_T_181[287:0] : _GEN_5953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7004 = 10'hb0 == _T_19 ? _ram_T_181[287:0] : _GEN_5954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7005 = 10'hb1 == _T_19 ? _ram_T_181[287:0] : _GEN_5955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7006 = 10'hb2 == _T_19 ? _ram_T_181[287:0] : _GEN_5956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7007 = 10'hb3 == _T_19 ? _ram_T_181[287:0] : _GEN_5957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7008 = 10'hb4 == _T_19 ? _ram_T_181[287:0] : _GEN_5958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7009 = 10'hb5 == _T_19 ? _ram_T_181[287:0] : _GEN_5959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7010 = 10'hb6 == _T_19 ? _ram_T_181[287:0] : _GEN_5960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7011 = 10'hb7 == _T_19 ? _ram_T_181[287:0] : _GEN_5961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7012 = 10'hb8 == _T_19 ? _ram_T_181[287:0] : _GEN_5962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7013 = 10'hb9 == _T_19 ? _ram_T_181[287:0] : _GEN_5963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7014 = 10'hba == _T_19 ? _ram_T_181[287:0] : _GEN_5964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7015 = 10'hbb == _T_19 ? _ram_T_181[287:0] : _GEN_5965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7016 = 10'hbc == _T_19 ? _ram_T_181[287:0] : _GEN_5966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7017 = 10'hbd == _T_19 ? _ram_T_181[287:0] : _GEN_5967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7018 = 10'hbe == _T_19 ? _ram_T_181[287:0] : _GEN_5968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7019 = 10'hbf == _T_19 ? _ram_T_181[287:0] : _GEN_5969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7020 = 10'hc0 == _T_19 ? _ram_T_181[287:0] : _GEN_5970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7021 = 10'hc1 == _T_19 ? _ram_T_181[287:0] : _GEN_5971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7022 = 10'hc2 == _T_19 ? _ram_T_181[287:0] : _GEN_5972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7023 = 10'hc3 == _T_19 ? _ram_T_181[287:0] : _GEN_5973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7024 = 10'hc4 == _T_19 ? _ram_T_181[287:0] : _GEN_5974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7025 = 10'hc5 == _T_19 ? _ram_T_181[287:0] : _GEN_5975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7026 = 10'hc6 == _T_19 ? _ram_T_181[287:0] : _GEN_5976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7027 = 10'hc7 == _T_19 ? _ram_T_181[287:0] : _GEN_5977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7028 = 10'hc8 == _T_19 ? _ram_T_181[287:0] : _GEN_5978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7029 = 10'hc9 == _T_19 ? _ram_T_181[287:0] : _GEN_5979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7030 = 10'hca == _T_19 ? _ram_T_181[287:0] : _GEN_5980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7031 = 10'hcb == _T_19 ? _ram_T_181[287:0] : _GEN_5981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7032 = 10'hcc == _T_19 ? _ram_T_181[287:0] : _GEN_5982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7033 = 10'hcd == _T_19 ? _ram_T_181[287:0] : _GEN_5983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7034 = 10'hce == _T_19 ? _ram_T_181[287:0] : _GEN_5984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7035 = 10'hcf == _T_19 ? _ram_T_181[287:0] : _GEN_5985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7036 = 10'hd0 == _T_19 ? _ram_T_181[287:0] : _GEN_5986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7037 = 10'hd1 == _T_19 ? _ram_T_181[287:0] : _GEN_5987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7038 = 10'hd2 == _T_19 ? _ram_T_181[287:0] : _GEN_5988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7039 = 10'hd3 == _T_19 ? _ram_T_181[287:0] : _GEN_5989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7040 = 10'hd4 == _T_19 ? _ram_T_181[287:0] : _GEN_5990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7041 = 10'hd5 == _T_19 ? _ram_T_181[287:0] : _GEN_5991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7042 = 10'hd6 == _T_19 ? _ram_T_181[287:0] : _GEN_5992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7043 = 10'hd7 == _T_19 ? _ram_T_181[287:0] : _GEN_5993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7044 = 10'hd8 == _T_19 ? _ram_T_181[287:0] : _GEN_5994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7045 = 10'hd9 == _T_19 ? _ram_T_181[287:0] : _GEN_5995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7046 = 10'hda == _T_19 ? _ram_T_181[287:0] : _GEN_5996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7047 = 10'hdb == _T_19 ? _ram_T_181[287:0] : _GEN_5997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7048 = 10'hdc == _T_19 ? _ram_T_181[287:0] : _GEN_5998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7049 = 10'hdd == _T_19 ? _ram_T_181[287:0] : _GEN_5999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7050 = 10'hde == _T_19 ? _ram_T_181[287:0] : _GEN_6000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7051 = 10'hdf == _T_19 ? _ram_T_181[287:0] : _GEN_6001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7052 = 10'he0 == _T_19 ? _ram_T_181[287:0] : _GEN_6002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7053 = 10'he1 == _T_19 ? _ram_T_181[287:0] : _GEN_6003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7054 = 10'he2 == _T_19 ? _ram_T_181[287:0] : _GEN_6004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7055 = 10'he3 == _T_19 ? _ram_T_181[287:0] : _GEN_6005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7056 = 10'he4 == _T_19 ? _ram_T_181[287:0] : _GEN_6006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7057 = 10'he5 == _T_19 ? _ram_T_181[287:0] : _GEN_6007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7058 = 10'he6 == _T_19 ? _ram_T_181[287:0] : _GEN_6008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7059 = 10'he7 == _T_19 ? _ram_T_181[287:0] : _GEN_6009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7060 = 10'he8 == _T_19 ? _ram_T_181[287:0] : _GEN_6010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7061 = 10'he9 == _T_19 ? _ram_T_181[287:0] : _GEN_6011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7062 = 10'hea == _T_19 ? _ram_T_181[287:0] : _GEN_6012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7063 = 10'heb == _T_19 ? _ram_T_181[287:0] : _GEN_6013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7064 = 10'hec == _T_19 ? _ram_T_181[287:0] : _GEN_6014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7065 = 10'hed == _T_19 ? _ram_T_181[287:0] : _GEN_6015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7066 = 10'hee == _T_19 ? _ram_T_181[287:0] : _GEN_6016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7067 = 10'hef == _T_19 ? _ram_T_181[287:0] : _GEN_6017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7068 = 10'hf0 == _T_19 ? _ram_T_181[287:0] : _GEN_6018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7069 = 10'hf1 == _T_19 ? _ram_T_181[287:0] : _GEN_6019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7070 = 10'hf2 == _T_19 ? _ram_T_181[287:0] : _GEN_6020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7071 = 10'hf3 == _T_19 ? _ram_T_181[287:0] : _GEN_6021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7072 = 10'hf4 == _T_19 ? _ram_T_181[287:0] : _GEN_6022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7073 = 10'hf5 == _T_19 ? _ram_T_181[287:0] : _GEN_6023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7074 = 10'hf6 == _T_19 ? _ram_T_181[287:0] : _GEN_6024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7075 = 10'hf7 == _T_19 ? _ram_T_181[287:0] : _GEN_6025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7076 = 10'hf8 == _T_19 ? _ram_T_181[287:0] : _GEN_6026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7077 = 10'hf9 == _T_19 ? _ram_T_181[287:0] : _GEN_6027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7078 = 10'hfa == _T_19 ? _ram_T_181[287:0] : _GEN_6028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7079 = 10'hfb == _T_19 ? _ram_T_181[287:0] : _GEN_6029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7080 = 10'hfc == _T_19 ? _ram_T_181[287:0] : _GEN_6030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7081 = 10'hfd == _T_19 ? _ram_T_181[287:0] : _GEN_6031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7082 = 10'hfe == _T_19 ? _ram_T_181[287:0] : _GEN_6032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7083 = 10'hff == _T_19 ? _ram_T_181[287:0] : _GEN_6033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7084 = 10'h100 == _T_19 ? _ram_T_181[287:0] : _GEN_6034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7085 = 10'h101 == _T_19 ? _ram_T_181[287:0] : _GEN_6035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7086 = 10'h102 == _T_19 ? _ram_T_181[287:0] : _GEN_6036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7087 = 10'h103 == _T_19 ? _ram_T_181[287:0] : _GEN_6037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7088 = 10'h104 == _T_19 ? _ram_T_181[287:0] : _GEN_6038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7089 = 10'h105 == _T_19 ? _ram_T_181[287:0] : _GEN_6039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7090 = 10'h106 == _T_19 ? _ram_T_181[287:0] : _GEN_6040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7091 = 10'h107 == _T_19 ? _ram_T_181[287:0] : _GEN_6041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7092 = 10'h108 == _T_19 ? _ram_T_181[287:0] : _GEN_6042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7093 = 10'h109 == _T_19 ? _ram_T_181[287:0] : _GEN_6043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7094 = 10'h10a == _T_19 ? _ram_T_181[287:0] : _GEN_6044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7095 = 10'h10b == _T_19 ? _ram_T_181[287:0] : _GEN_6045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7096 = 10'h10c == _T_19 ? _ram_T_181[287:0] : _GEN_6046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7097 = 10'h10d == _T_19 ? _ram_T_181[287:0] : _GEN_6047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7098 = 10'h10e == _T_19 ? _ram_T_181[287:0] : _GEN_6048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7099 = 10'h10f == _T_19 ? _ram_T_181[287:0] : _GEN_6049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7100 = 10'h110 == _T_19 ? _ram_T_181[287:0] : _GEN_6050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7101 = 10'h111 == _T_19 ? _ram_T_181[287:0] : _GEN_6051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7102 = 10'h112 == _T_19 ? _ram_T_181[287:0] : _GEN_6052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7103 = 10'h113 == _T_19 ? _ram_T_181[287:0] : _GEN_6053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7104 = 10'h114 == _T_19 ? _ram_T_181[287:0] : _GEN_6054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7105 = 10'h115 == _T_19 ? _ram_T_181[287:0] : _GEN_6055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7106 = 10'h116 == _T_19 ? _ram_T_181[287:0] : _GEN_6056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7107 = 10'h117 == _T_19 ? _ram_T_181[287:0] : _GEN_6057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7108 = 10'h118 == _T_19 ? _ram_T_181[287:0] : _GEN_6058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7109 = 10'h119 == _T_19 ? _ram_T_181[287:0] : _GEN_6059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7110 = 10'h11a == _T_19 ? _ram_T_181[287:0] : _GEN_6060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7111 = 10'h11b == _T_19 ? _ram_T_181[287:0] : _GEN_6061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7112 = 10'h11c == _T_19 ? _ram_T_181[287:0] : _GEN_6062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7113 = 10'h11d == _T_19 ? _ram_T_181[287:0] : _GEN_6063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7114 = 10'h11e == _T_19 ? _ram_T_181[287:0] : _GEN_6064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7115 = 10'h11f == _T_19 ? _ram_T_181[287:0] : _GEN_6065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7116 = 10'h120 == _T_19 ? _ram_T_181[287:0] : _GEN_6066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7117 = 10'h121 == _T_19 ? _ram_T_181[287:0] : _GEN_6067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7118 = 10'h122 == _T_19 ? _ram_T_181[287:0] : _GEN_6068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7119 = 10'h123 == _T_19 ? _ram_T_181[287:0] : _GEN_6069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7120 = 10'h124 == _T_19 ? _ram_T_181[287:0] : _GEN_6070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7121 = 10'h125 == _T_19 ? _ram_T_181[287:0] : _GEN_6071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7122 = 10'h126 == _T_19 ? _ram_T_181[287:0] : _GEN_6072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7123 = 10'h127 == _T_19 ? _ram_T_181[287:0] : _GEN_6073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7124 = 10'h128 == _T_19 ? _ram_T_181[287:0] : _GEN_6074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7125 = 10'h129 == _T_19 ? _ram_T_181[287:0] : _GEN_6075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7126 = 10'h12a == _T_19 ? _ram_T_181[287:0] : _GEN_6076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7127 = 10'h12b == _T_19 ? _ram_T_181[287:0] : _GEN_6077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7128 = 10'h12c == _T_19 ? _ram_T_181[287:0] : _GEN_6078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7129 = 10'h12d == _T_19 ? _ram_T_181[287:0] : _GEN_6079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7130 = 10'h12e == _T_19 ? _ram_T_181[287:0] : _GEN_6080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7131 = 10'h12f == _T_19 ? _ram_T_181[287:0] : _GEN_6081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7132 = 10'h130 == _T_19 ? _ram_T_181[287:0] : _GEN_6082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7133 = 10'h131 == _T_19 ? _ram_T_181[287:0] : _GEN_6083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7134 = 10'h132 == _T_19 ? _ram_T_181[287:0] : _GEN_6084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7135 = 10'h133 == _T_19 ? _ram_T_181[287:0] : _GEN_6085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7136 = 10'h134 == _T_19 ? _ram_T_181[287:0] : _GEN_6086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7137 = 10'h135 == _T_19 ? _ram_T_181[287:0] : _GEN_6087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7138 = 10'h136 == _T_19 ? _ram_T_181[287:0] : _GEN_6088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7139 = 10'h137 == _T_19 ? _ram_T_181[287:0] : _GEN_6089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7140 = 10'h138 == _T_19 ? _ram_T_181[287:0] : _GEN_6090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7141 = 10'h139 == _T_19 ? _ram_T_181[287:0] : _GEN_6091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7142 = 10'h13a == _T_19 ? _ram_T_181[287:0] : _GEN_6092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7143 = 10'h13b == _T_19 ? _ram_T_181[287:0] : _GEN_6093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7144 = 10'h13c == _T_19 ? _ram_T_181[287:0] : _GEN_6094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7145 = 10'h13d == _T_19 ? _ram_T_181[287:0] : _GEN_6095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7146 = 10'h13e == _T_19 ? _ram_T_181[287:0] : _GEN_6096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7147 = 10'h13f == _T_19 ? _ram_T_181[287:0] : _GEN_6097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7148 = 10'h140 == _T_19 ? _ram_T_181[287:0] : _GEN_6098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7149 = 10'h141 == _T_19 ? _ram_T_181[287:0] : _GEN_6099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7150 = 10'h142 == _T_19 ? _ram_T_181[287:0] : _GEN_6100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7151 = 10'h143 == _T_19 ? _ram_T_181[287:0] : _GEN_6101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7152 = 10'h144 == _T_19 ? _ram_T_181[287:0] : _GEN_6102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7153 = 10'h145 == _T_19 ? _ram_T_181[287:0] : _GEN_6103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7154 = 10'h146 == _T_19 ? _ram_T_181[287:0] : _GEN_6104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7155 = 10'h147 == _T_19 ? _ram_T_181[287:0] : _GEN_6105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7156 = 10'h148 == _T_19 ? _ram_T_181[287:0] : _GEN_6106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7157 = 10'h149 == _T_19 ? _ram_T_181[287:0] : _GEN_6107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7158 = 10'h14a == _T_19 ? _ram_T_181[287:0] : _GEN_6108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7159 = 10'h14b == _T_19 ? _ram_T_181[287:0] : _GEN_6109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7160 = 10'h14c == _T_19 ? _ram_T_181[287:0] : _GEN_6110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7161 = 10'h14d == _T_19 ? _ram_T_181[287:0] : _GEN_6111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7162 = 10'h14e == _T_19 ? _ram_T_181[287:0] : _GEN_6112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7163 = 10'h14f == _T_19 ? _ram_T_181[287:0] : _GEN_6113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7164 = 10'h150 == _T_19 ? _ram_T_181[287:0] : _GEN_6114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7165 = 10'h151 == _T_19 ? _ram_T_181[287:0] : _GEN_6115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7166 = 10'h152 == _T_19 ? _ram_T_181[287:0] : _GEN_6116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7167 = 10'h153 == _T_19 ? _ram_T_181[287:0] : _GEN_6117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7168 = 10'h154 == _T_19 ? _ram_T_181[287:0] : _GEN_6118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7169 = 10'h155 == _T_19 ? _ram_T_181[287:0] : _GEN_6119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7170 = 10'h156 == _T_19 ? _ram_T_181[287:0] : _GEN_6120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7171 = 10'h157 == _T_19 ? _ram_T_181[287:0] : _GEN_6121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7172 = 10'h158 == _T_19 ? _ram_T_181[287:0] : _GEN_6122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7173 = 10'h159 == _T_19 ? _ram_T_181[287:0] : _GEN_6123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7174 = 10'h15a == _T_19 ? _ram_T_181[287:0] : _GEN_6124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7175 = 10'h15b == _T_19 ? _ram_T_181[287:0] : _GEN_6125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7176 = 10'h15c == _T_19 ? _ram_T_181[287:0] : _GEN_6126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7177 = 10'h15d == _T_19 ? _ram_T_181[287:0] : _GEN_6127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7178 = 10'h15e == _T_19 ? _ram_T_181[287:0] : _GEN_6128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7179 = 10'h15f == _T_19 ? _ram_T_181[287:0] : _GEN_6129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7180 = 10'h160 == _T_19 ? _ram_T_181[287:0] : _GEN_6130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7181 = 10'h161 == _T_19 ? _ram_T_181[287:0] : _GEN_6131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7182 = 10'h162 == _T_19 ? _ram_T_181[287:0] : _GEN_6132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7183 = 10'h163 == _T_19 ? _ram_T_181[287:0] : _GEN_6133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7184 = 10'h164 == _T_19 ? _ram_T_181[287:0] : _GEN_6134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7185 = 10'h165 == _T_19 ? _ram_T_181[287:0] : _GEN_6135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7186 = 10'h166 == _T_19 ? _ram_T_181[287:0] : _GEN_6136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7187 = 10'h167 == _T_19 ? _ram_T_181[287:0] : _GEN_6137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7188 = 10'h168 == _T_19 ? _ram_T_181[287:0] : _GEN_6138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7189 = 10'h169 == _T_19 ? _ram_T_181[287:0] : _GEN_6139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7190 = 10'h16a == _T_19 ? _ram_T_181[287:0] : _GEN_6140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7191 = 10'h16b == _T_19 ? _ram_T_181[287:0] : _GEN_6141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7192 = 10'h16c == _T_19 ? _ram_T_181[287:0] : _GEN_6142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7193 = 10'h16d == _T_19 ? _ram_T_181[287:0] : _GEN_6143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7194 = 10'h16e == _T_19 ? _ram_T_181[287:0] : _GEN_6144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7195 = 10'h16f == _T_19 ? _ram_T_181[287:0] : _GEN_6145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7196 = 10'h170 == _T_19 ? _ram_T_181[287:0] : _GEN_6146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7197 = 10'h171 == _T_19 ? _ram_T_181[287:0] : _GEN_6147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7198 = 10'h172 == _T_19 ? _ram_T_181[287:0] : _GEN_6148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7199 = 10'h173 == _T_19 ? _ram_T_181[287:0] : _GEN_6149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7200 = 10'h174 == _T_19 ? _ram_T_181[287:0] : _GEN_6150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7201 = 10'h175 == _T_19 ? _ram_T_181[287:0] : _GEN_6151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7202 = 10'h176 == _T_19 ? _ram_T_181[287:0] : _GEN_6152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7203 = 10'h177 == _T_19 ? _ram_T_181[287:0] : _GEN_6153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7204 = 10'h178 == _T_19 ? _ram_T_181[287:0] : _GEN_6154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7205 = 10'h179 == _T_19 ? _ram_T_181[287:0] : _GEN_6155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7206 = 10'h17a == _T_19 ? _ram_T_181[287:0] : _GEN_6156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7207 = 10'h17b == _T_19 ? _ram_T_181[287:0] : _GEN_6157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7208 = 10'h17c == _T_19 ? _ram_T_181[287:0] : _GEN_6158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7209 = 10'h17d == _T_19 ? _ram_T_181[287:0] : _GEN_6159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7210 = 10'h17e == _T_19 ? _ram_T_181[287:0] : _GEN_6160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7211 = 10'h17f == _T_19 ? _ram_T_181[287:0] : _GEN_6161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7212 = 10'h180 == _T_19 ? _ram_T_181[287:0] : _GEN_6162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7213 = 10'h181 == _T_19 ? _ram_T_181[287:0] : _GEN_6163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7214 = 10'h182 == _T_19 ? _ram_T_181[287:0] : _GEN_6164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7215 = 10'h183 == _T_19 ? _ram_T_181[287:0] : _GEN_6165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7216 = 10'h184 == _T_19 ? _ram_T_181[287:0] : _GEN_6166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7217 = 10'h185 == _T_19 ? _ram_T_181[287:0] : _GEN_6167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7218 = 10'h186 == _T_19 ? _ram_T_181[287:0] : _GEN_6168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7219 = 10'h187 == _T_19 ? _ram_T_181[287:0] : _GEN_6169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7220 = 10'h188 == _T_19 ? _ram_T_181[287:0] : _GEN_6170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7221 = 10'h189 == _T_19 ? _ram_T_181[287:0] : _GEN_6171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7222 = 10'h18a == _T_19 ? _ram_T_181[287:0] : _GEN_6172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7223 = 10'h18b == _T_19 ? _ram_T_181[287:0] : _GEN_6173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7224 = 10'h18c == _T_19 ? _ram_T_181[287:0] : _GEN_6174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7225 = 10'h18d == _T_19 ? _ram_T_181[287:0] : _GEN_6175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7226 = 10'h18e == _T_19 ? _ram_T_181[287:0] : _GEN_6176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7227 = 10'h18f == _T_19 ? _ram_T_181[287:0] : _GEN_6177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7228 = 10'h190 == _T_19 ? _ram_T_181[287:0] : _GEN_6178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7229 = 10'h191 == _T_19 ? _ram_T_181[287:0] : _GEN_6179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7230 = 10'h192 == _T_19 ? _ram_T_181[287:0] : _GEN_6180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7231 = 10'h193 == _T_19 ? _ram_T_181[287:0] : _GEN_6181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7232 = 10'h194 == _T_19 ? _ram_T_181[287:0] : _GEN_6182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7233 = 10'h195 == _T_19 ? _ram_T_181[287:0] : _GEN_6183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7234 = 10'h196 == _T_19 ? _ram_T_181[287:0] : _GEN_6184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7235 = 10'h197 == _T_19 ? _ram_T_181[287:0] : _GEN_6185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7236 = 10'h198 == _T_19 ? _ram_T_181[287:0] : _GEN_6186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7237 = 10'h199 == _T_19 ? _ram_T_181[287:0] : _GEN_6187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7238 = 10'h19a == _T_19 ? _ram_T_181[287:0] : _GEN_6188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7239 = 10'h19b == _T_19 ? _ram_T_181[287:0] : _GEN_6189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7240 = 10'h19c == _T_19 ? _ram_T_181[287:0] : _GEN_6190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7241 = 10'h19d == _T_19 ? _ram_T_181[287:0] : _GEN_6191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7242 = 10'h19e == _T_19 ? _ram_T_181[287:0] : _GEN_6192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7243 = 10'h19f == _T_19 ? _ram_T_181[287:0] : _GEN_6193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7244 = 10'h1a0 == _T_19 ? _ram_T_181[287:0] : _GEN_6194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7245 = 10'h1a1 == _T_19 ? _ram_T_181[287:0] : _GEN_6195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7246 = 10'h1a2 == _T_19 ? _ram_T_181[287:0] : _GEN_6196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7247 = 10'h1a3 == _T_19 ? _ram_T_181[287:0] : _GEN_6197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7248 = 10'h1a4 == _T_19 ? _ram_T_181[287:0] : _GEN_6198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7249 = 10'h1a5 == _T_19 ? _ram_T_181[287:0] : _GEN_6199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7250 = 10'h1a6 == _T_19 ? _ram_T_181[287:0] : _GEN_6200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7251 = 10'h1a7 == _T_19 ? _ram_T_181[287:0] : _GEN_6201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7252 = 10'h1a8 == _T_19 ? _ram_T_181[287:0] : _GEN_6202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7253 = 10'h1a9 == _T_19 ? _ram_T_181[287:0] : _GEN_6203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7254 = 10'h1aa == _T_19 ? _ram_T_181[287:0] : _GEN_6204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7255 = 10'h1ab == _T_19 ? _ram_T_181[287:0] : _GEN_6205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7256 = 10'h1ac == _T_19 ? _ram_T_181[287:0] : _GEN_6206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7257 = 10'h1ad == _T_19 ? _ram_T_181[287:0] : _GEN_6207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7258 = 10'h1ae == _T_19 ? _ram_T_181[287:0] : _GEN_6208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7259 = 10'h1af == _T_19 ? _ram_T_181[287:0] : _GEN_6209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7260 = 10'h1b0 == _T_19 ? _ram_T_181[287:0] : _GEN_6210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7261 = 10'h1b1 == _T_19 ? _ram_T_181[287:0] : _GEN_6211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7262 = 10'h1b2 == _T_19 ? _ram_T_181[287:0] : _GEN_6212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7263 = 10'h1b3 == _T_19 ? _ram_T_181[287:0] : _GEN_6213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7264 = 10'h1b4 == _T_19 ? _ram_T_181[287:0] : _GEN_6214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7265 = 10'h1b5 == _T_19 ? _ram_T_181[287:0] : _GEN_6215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7266 = 10'h1b6 == _T_19 ? _ram_T_181[287:0] : _GEN_6216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7267 = 10'h1b7 == _T_19 ? _ram_T_181[287:0] : _GEN_6217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7268 = 10'h1b8 == _T_19 ? _ram_T_181[287:0] : _GEN_6218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7269 = 10'h1b9 == _T_19 ? _ram_T_181[287:0] : _GEN_6219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7270 = 10'h1ba == _T_19 ? _ram_T_181[287:0] : _GEN_6220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7271 = 10'h1bb == _T_19 ? _ram_T_181[287:0] : _GEN_6221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7272 = 10'h1bc == _T_19 ? _ram_T_181[287:0] : _GEN_6222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7273 = 10'h1bd == _T_19 ? _ram_T_181[287:0] : _GEN_6223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7274 = 10'h1be == _T_19 ? _ram_T_181[287:0] : _GEN_6224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7275 = 10'h1bf == _T_19 ? _ram_T_181[287:0] : _GEN_6225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7276 = 10'h1c0 == _T_19 ? _ram_T_181[287:0] : _GEN_6226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7277 = 10'h1c1 == _T_19 ? _ram_T_181[287:0] : _GEN_6227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7278 = 10'h1c2 == _T_19 ? _ram_T_181[287:0] : _GEN_6228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7279 = 10'h1c3 == _T_19 ? _ram_T_181[287:0] : _GEN_6229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7280 = 10'h1c4 == _T_19 ? _ram_T_181[287:0] : _GEN_6230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7281 = 10'h1c5 == _T_19 ? _ram_T_181[287:0] : _GEN_6231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7282 = 10'h1c6 == _T_19 ? _ram_T_181[287:0] : _GEN_6232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7283 = 10'h1c7 == _T_19 ? _ram_T_181[287:0] : _GEN_6233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7284 = 10'h1c8 == _T_19 ? _ram_T_181[287:0] : _GEN_6234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7285 = 10'h1c9 == _T_19 ? _ram_T_181[287:0] : _GEN_6235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7286 = 10'h1ca == _T_19 ? _ram_T_181[287:0] : _GEN_6236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7287 = 10'h1cb == _T_19 ? _ram_T_181[287:0] : _GEN_6237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7288 = 10'h1cc == _T_19 ? _ram_T_181[287:0] : _GEN_6238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7289 = 10'h1cd == _T_19 ? _ram_T_181[287:0] : _GEN_6239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7290 = 10'h1ce == _T_19 ? _ram_T_181[287:0] : _GEN_6240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7291 = 10'h1cf == _T_19 ? _ram_T_181[287:0] : _GEN_6241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7292 = 10'h1d0 == _T_19 ? _ram_T_181[287:0] : _GEN_6242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7293 = 10'h1d1 == _T_19 ? _ram_T_181[287:0] : _GEN_6243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7294 = 10'h1d2 == _T_19 ? _ram_T_181[287:0] : _GEN_6244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7295 = 10'h1d3 == _T_19 ? _ram_T_181[287:0] : _GEN_6245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7296 = 10'h1d4 == _T_19 ? _ram_T_181[287:0] : _GEN_6246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7297 = 10'h1d5 == _T_19 ? _ram_T_181[287:0] : _GEN_6247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7298 = 10'h1d6 == _T_19 ? _ram_T_181[287:0] : _GEN_6248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7299 = 10'h1d7 == _T_19 ? _ram_T_181[287:0] : _GEN_6249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7300 = 10'h1d8 == _T_19 ? _ram_T_181[287:0] : _GEN_6250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7301 = 10'h1d9 == _T_19 ? _ram_T_181[287:0] : _GEN_6251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7302 = 10'h1da == _T_19 ? _ram_T_181[287:0] : _GEN_6252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7303 = 10'h1db == _T_19 ? _ram_T_181[287:0] : _GEN_6253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7304 = 10'h1dc == _T_19 ? _ram_T_181[287:0] : _GEN_6254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7305 = 10'h1dd == _T_19 ? _ram_T_181[287:0] : _GEN_6255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7306 = 10'h1de == _T_19 ? _ram_T_181[287:0] : _GEN_6256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7307 = 10'h1df == _T_19 ? _ram_T_181[287:0] : _GEN_6257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7308 = 10'h1e0 == _T_19 ? _ram_T_181[287:0] : _GEN_6258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7309 = 10'h1e1 == _T_19 ? _ram_T_181[287:0] : _GEN_6259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7310 = 10'h1e2 == _T_19 ? _ram_T_181[287:0] : _GEN_6260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7311 = 10'h1e3 == _T_19 ? _ram_T_181[287:0] : _GEN_6261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7312 = 10'h1e4 == _T_19 ? _ram_T_181[287:0] : _GEN_6262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7313 = 10'h1e5 == _T_19 ? _ram_T_181[287:0] : _GEN_6263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7314 = 10'h1e6 == _T_19 ? _ram_T_181[287:0] : _GEN_6264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7315 = 10'h1e7 == _T_19 ? _ram_T_181[287:0] : _GEN_6265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7316 = 10'h1e8 == _T_19 ? _ram_T_181[287:0] : _GEN_6266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7317 = 10'h1e9 == _T_19 ? _ram_T_181[287:0] : _GEN_6267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7318 = 10'h1ea == _T_19 ? _ram_T_181[287:0] : _GEN_6268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7319 = 10'h1eb == _T_19 ? _ram_T_181[287:0] : _GEN_6269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7320 = 10'h1ec == _T_19 ? _ram_T_181[287:0] : _GEN_6270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7321 = 10'h1ed == _T_19 ? _ram_T_181[287:0] : _GEN_6271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7322 = 10'h1ee == _T_19 ? _ram_T_181[287:0] : _GEN_6272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7323 = 10'h1ef == _T_19 ? _ram_T_181[287:0] : _GEN_6273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7324 = 10'h1f0 == _T_19 ? _ram_T_181[287:0] : _GEN_6274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7325 = 10'h1f1 == _T_19 ? _ram_T_181[287:0] : _GEN_6275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7326 = 10'h1f2 == _T_19 ? _ram_T_181[287:0] : _GEN_6276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7327 = 10'h1f3 == _T_19 ? _ram_T_181[287:0] : _GEN_6277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7328 = 10'h1f4 == _T_19 ? _ram_T_181[287:0] : _GEN_6278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7329 = 10'h1f5 == _T_19 ? _ram_T_181[287:0] : _GEN_6279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7330 = 10'h1f6 == _T_19 ? _ram_T_181[287:0] : _GEN_6280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7331 = 10'h1f7 == _T_19 ? _ram_T_181[287:0] : _GEN_6281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7332 = 10'h1f8 == _T_19 ? _ram_T_181[287:0] : _GEN_6282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7333 = 10'h1f9 == _T_19 ? _ram_T_181[287:0] : _GEN_6283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7334 = 10'h1fa == _T_19 ? _ram_T_181[287:0] : _GEN_6284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7335 = 10'h1fb == _T_19 ? _ram_T_181[287:0] : _GEN_6285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7336 = 10'h1fc == _T_19 ? _ram_T_181[287:0] : _GEN_6286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7337 = 10'h1fd == _T_19 ? _ram_T_181[287:0] : _GEN_6287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7338 = 10'h1fe == _T_19 ? _ram_T_181[287:0] : _GEN_6288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7339 = 10'h1ff == _T_19 ? _ram_T_181[287:0] : _GEN_6289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7340 = 10'h200 == _T_19 ? _ram_T_181[287:0] : _GEN_6290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7341 = 10'h201 == _T_19 ? _ram_T_181[287:0] : _GEN_6291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7342 = 10'h202 == _T_19 ? _ram_T_181[287:0] : _GEN_6292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7343 = 10'h203 == _T_19 ? _ram_T_181[287:0] : _GEN_6293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7344 = 10'h204 == _T_19 ? _ram_T_181[287:0] : _GEN_6294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7345 = 10'h205 == _T_19 ? _ram_T_181[287:0] : _GEN_6295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7346 = 10'h206 == _T_19 ? _ram_T_181[287:0] : _GEN_6296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7347 = 10'h207 == _T_19 ? _ram_T_181[287:0] : _GEN_6297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7348 = 10'h208 == _T_19 ? _ram_T_181[287:0] : _GEN_6298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7349 = 10'h209 == _T_19 ? _ram_T_181[287:0] : _GEN_6299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7350 = 10'h20a == _T_19 ? _ram_T_181[287:0] : _GEN_6300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7351 = 10'h20b == _T_19 ? _ram_T_181[287:0] : _GEN_6301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7352 = 10'h20c == _T_19 ? _ram_T_181[287:0] : _GEN_6302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_21 = h + 10'h7; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_7 = vga_mem_ram_MPORT_63_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_7 = vga_mem_ram_MPORT_64_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_7 = vga_mem_ram_MPORT_65_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_7 = vga_mem_ram_MPORT_66_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_7 = vga_mem_ram_MPORT_67_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_7 = vga_mem_ram_MPORT_68_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_7 = vga_mem_ram_MPORT_69_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_7 = vga_mem_ram_MPORT_70_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_7 = vga_mem_ram_MPORT_71_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_202 = {278'h0,ram_hi_hi_hi_lo_7,ram_hi_hi_lo_7,ram_hi_lo_hi_7,ram_hi_lo_lo_7,ram_lo_hi_hi_hi_7,
    ram_lo_hi_hi_lo_7,ram_lo_hi_lo_7,ram_lo_lo_hi_7,ram_lo_lo_lo_7}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19074 = {{8191'd0}, _ram_T_202}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_206 = _GEN_19074 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_7354 = 10'h1 == _T_21 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7355 = 10'h2 == _T_21 ? ram_2 : _GEN_7354; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7356 = 10'h3 == _T_21 ? ram_3 : _GEN_7355; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7357 = 10'h4 == _T_21 ? ram_4 : _GEN_7356; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7358 = 10'h5 == _T_21 ? ram_5 : _GEN_7357; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7359 = 10'h6 == _T_21 ? ram_6 : _GEN_7358; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7360 = 10'h7 == _T_21 ? ram_7 : _GEN_7359; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7361 = 10'h8 == _T_21 ? ram_8 : _GEN_7360; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7362 = 10'h9 == _T_21 ? ram_9 : _GEN_7361; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7363 = 10'ha == _T_21 ? ram_10 : _GEN_7362; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7364 = 10'hb == _T_21 ? ram_11 : _GEN_7363; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7365 = 10'hc == _T_21 ? ram_12 : _GEN_7364; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7366 = 10'hd == _T_21 ? ram_13 : _GEN_7365; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7367 = 10'he == _T_21 ? ram_14 : _GEN_7366; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7368 = 10'hf == _T_21 ? ram_15 : _GEN_7367; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7369 = 10'h10 == _T_21 ? ram_16 : _GEN_7368; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7370 = 10'h11 == _T_21 ? ram_17 : _GEN_7369; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7371 = 10'h12 == _T_21 ? ram_18 : _GEN_7370; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7372 = 10'h13 == _T_21 ? ram_19 : _GEN_7371; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7373 = 10'h14 == _T_21 ? ram_20 : _GEN_7372; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7374 = 10'h15 == _T_21 ? ram_21 : _GEN_7373; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7375 = 10'h16 == _T_21 ? ram_22 : _GEN_7374; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7376 = 10'h17 == _T_21 ? ram_23 : _GEN_7375; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7377 = 10'h18 == _T_21 ? ram_24 : _GEN_7376; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7378 = 10'h19 == _T_21 ? ram_25 : _GEN_7377; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7379 = 10'h1a == _T_21 ? ram_26 : _GEN_7378; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7380 = 10'h1b == _T_21 ? ram_27 : _GEN_7379; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7381 = 10'h1c == _T_21 ? ram_28 : _GEN_7380; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7382 = 10'h1d == _T_21 ? ram_29 : _GEN_7381; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7383 = 10'h1e == _T_21 ? ram_30 : _GEN_7382; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7384 = 10'h1f == _T_21 ? ram_31 : _GEN_7383; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7385 = 10'h20 == _T_21 ? ram_32 : _GEN_7384; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7386 = 10'h21 == _T_21 ? ram_33 : _GEN_7385; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7387 = 10'h22 == _T_21 ? ram_34 : _GEN_7386; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7388 = 10'h23 == _T_21 ? ram_35 : _GEN_7387; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7389 = 10'h24 == _T_21 ? ram_36 : _GEN_7388; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7390 = 10'h25 == _T_21 ? ram_37 : _GEN_7389; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7391 = 10'h26 == _T_21 ? ram_38 : _GEN_7390; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7392 = 10'h27 == _T_21 ? ram_39 : _GEN_7391; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7393 = 10'h28 == _T_21 ? ram_40 : _GEN_7392; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7394 = 10'h29 == _T_21 ? ram_41 : _GEN_7393; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7395 = 10'h2a == _T_21 ? ram_42 : _GEN_7394; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7396 = 10'h2b == _T_21 ? ram_43 : _GEN_7395; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7397 = 10'h2c == _T_21 ? ram_44 : _GEN_7396; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7398 = 10'h2d == _T_21 ? ram_45 : _GEN_7397; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7399 = 10'h2e == _T_21 ? ram_46 : _GEN_7398; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7400 = 10'h2f == _T_21 ? ram_47 : _GEN_7399; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7401 = 10'h30 == _T_21 ? ram_48 : _GEN_7400; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7402 = 10'h31 == _T_21 ? ram_49 : _GEN_7401; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7403 = 10'h32 == _T_21 ? ram_50 : _GEN_7402; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7404 = 10'h33 == _T_21 ? ram_51 : _GEN_7403; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7405 = 10'h34 == _T_21 ? ram_52 : _GEN_7404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7406 = 10'h35 == _T_21 ? ram_53 : _GEN_7405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7407 = 10'h36 == _T_21 ? ram_54 : _GEN_7406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7408 = 10'h37 == _T_21 ? ram_55 : _GEN_7407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7409 = 10'h38 == _T_21 ? ram_56 : _GEN_7408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7410 = 10'h39 == _T_21 ? ram_57 : _GEN_7409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7411 = 10'h3a == _T_21 ? ram_58 : _GEN_7410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7412 = 10'h3b == _T_21 ? ram_59 : _GEN_7411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7413 = 10'h3c == _T_21 ? ram_60 : _GEN_7412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7414 = 10'h3d == _T_21 ? ram_61 : _GEN_7413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7415 = 10'h3e == _T_21 ? ram_62 : _GEN_7414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7416 = 10'h3f == _T_21 ? ram_63 : _GEN_7415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7417 = 10'h40 == _T_21 ? ram_64 : _GEN_7416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7418 = 10'h41 == _T_21 ? ram_65 : _GEN_7417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7419 = 10'h42 == _T_21 ? ram_66 : _GEN_7418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7420 = 10'h43 == _T_21 ? ram_67 : _GEN_7419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7421 = 10'h44 == _T_21 ? ram_68 : _GEN_7420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7422 = 10'h45 == _T_21 ? ram_69 : _GEN_7421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7423 = 10'h46 == _T_21 ? ram_70 : _GEN_7422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7424 = 10'h47 == _T_21 ? ram_71 : _GEN_7423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7425 = 10'h48 == _T_21 ? ram_72 : _GEN_7424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7426 = 10'h49 == _T_21 ? ram_73 : _GEN_7425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7427 = 10'h4a == _T_21 ? ram_74 : _GEN_7426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7428 = 10'h4b == _T_21 ? ram_75 : _GEN_7427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7429 = 10'h4c == _T_21 ? ram_76 : _GEN_7428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7430 = 10'h4d == _T_21 ? ram_77 : _GEN_7429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7431 = 10'h4e == _T_21 ? ram_78 : _GEN_7430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7432 = 10'h4f == _T_21 ? ram_79 : _GEN_7431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7433 = 10'h50 == _T_21 ? ram_80 : _GEN_7432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7434 = 10'h51 == _T_21 ? ram_81 : _GEN_7433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7435 = 10'h52 == _T_21 ? ram_82 : _GEN_7434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7436 = 10'h53 == _T_21 ? ram_83 : _GEN_7435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7437 = 10'h54 == _T_21 ? ram_84 : _GEN_7436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7438 = 10'h55 == _T_21 ? ram_85 : _GEN_7437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7439 = 10'h56 == _T_21 ? ram_86 : _GEN_7438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7440 = 10'h57 == _T_21 ? ram_87 : _GEN_7439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7441 = 10'h58 == _T_21 ? ram_88 : _GEN_7440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7442 = 10'h59 == _T_21 ? ram_89 : _GEN_7441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7443 = 10'h5a == _T_21 ? ram_90 : _GEN_7442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7444 = 10'h5b == _T_21 ? ram_91 : _GEN_7443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7445 = 10'h5c == _T_21 ? ram_92 : _GEN_7444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7446 = 10'h5d == _T_21 ? ram_93 : _GEN_7445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7447 = 10'h5e == _T_21 ? ram_94 : _GEN_7446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7448 = 10'h5f == _T_21 ? ram_95 : _GEN_7447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7449 = 10'h60 == _T_21 ? ram_96 : _GEN_7448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7450 = 10'h61 == _T_21 ? ram_97 : _GEN_7449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7451 = 10'h62 == _T_21 ? ram_98 : _GEN_7450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7452 = 10'h63 == _T_21 ? ram_99 : _GEN_7451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7453 = 10'h64 == _T_21 ? ram_100 : _GEN_7452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7454 = 10'h65 == _T_21 ? ram_101 : _GEN_7453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7455 = 10'h66 == _T_21 ? ram_102 : _GEN_7454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7456 = 10'h67 == _T_21 ? ram_103 : _GEN_7455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7457 = 10'h68 == _T_21 ? ram_104 : _GEN_7456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7458 = 10'h69 == _T_21 ? ram_105 : _GEN_7457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7459 = 10'h6a == _T_21 ? ram_106 : _GEN_7458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7460 = 10'h6b == _T_21 ? ram_107 : _GEN_7459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7461 = 10'h6c == _T_21 ? ram_108 : _GEN_7460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7462 = 10'h6d == _T_21 ? ram_109 : _GEN_7461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7463 = 10'h6e == _T_21 ? ram_110 : _GEN_7462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7464 = 10'h6f == _T_21 ? ram_111 : _GEN_7463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7465 = 10'h70 == _T_21 ? ram_112 : _GEN_7464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7466 = 10'h71 == _T_21 ? ram_113 : _GEN_7465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7467 = 10'h72 == _T_21 ? ram_114 : _GEN_7466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7468 = 10'h73 == _T_21 ? ram_115 : _GEN_7467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7469 = 10'h74 == _T_21 ? ram_116 : _GEN_7468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7470 = 10'h75 == _T_21 ? ram_117 : _GEN_7469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7471 = 10'h76 == _T_21 ? ram_118 : _GEN_7470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7472 = 10'h77 == _T_21 ? ram_119 : _GEN_7471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7473 = 10'h78 == _T_21 ? ram_120 : _GEN_7472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7474 = 10'h79 == _T_21 ? ram_121 : _GEN_7473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7475 = 10'h7a == _T_21 ? ram_122 : _GEN_7474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7476 = 10'h7b == _T_21 ? ram_123 : _GEN_7475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7477 = 10'h7c == _T_21 ? ram_124 : _GEN_7476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7478 = 10'h7d == _T_21 ? ram_125 : _GEN_7477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7479 = 10'h7e == _T_21 ? ram_126 : _GEN_7478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7480 = 10'h7f == _T_21 ? ram_127 : _GEN_7479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7481 = 10'h80 == _T_21 ? ram_128 : _GEN_7480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7482 = 10'h81 == _T_21 ? ram_129 : _GEN_7481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7483 = 10'h82 == _T_21 ? ram_130 : _GEN_7482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7484 = 10'h83 == _T_21 ? ram_131 : _GEN_7483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7485 = 10'h84 == _T_21 ? ram_132 : _GEN_7484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7486 = 10'h85 == _T_21 ? ram_133 : _GEN_7485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7487 = 10'h86 == _T_21 ? ram_134 : _GEN_7486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7488 = 10'h87 == _T_21 ? ram_135 : _GEN_7487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7489 = 10'h88 == _T_21 ? ram_136 : _GEN_7488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7490 = 10'h89 == _T_21 ? ram_137 : _GEN_7489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7491 = 10'h8a == _T_21 ? ram_138 : _GEN_7490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7492 = 10'h8b == _T_21 ? ram_139 : _GEN_7491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7493 = 10'h8c == _T_21 ? ram_140 : _GEN_7492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7494 = 10'h8d == _T_21 ? ram_141 : _GEN_7493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7495 = 10'h8e == _T_21 ? ram_142 : _GEN_7494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7496 = 10'h8f == _T_21 ? ram_143 : _GEN_7495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7497 = 10'h90 == _T_21 ? ram_144 : _GEN_7496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7498 = 10'h91 == _T_21 ? ram_145 : _GEN_7497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7499 = 10'h92 == _T_21 ? ram_146 : _GEN_7498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7500 = 10'h93 == _T_21 ? ram_147 : _GEN_7499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7501 = 10'h94 == _T_21 ? ram_148 : _GEN_7500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7502 = 10'h95 == _T_21 ? ram_149 : _GEN_7501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7503 = 10'h96 == _T_21 ? ram_150 : _GEN_7502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7504 = 10'h97 == _T_21 ? ram_151 : _GEN_7503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7505 = 10'h98 == _T_21 ? ram_152 : _GEN_7504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7506 = 10'h99 == _T_21 ? ram_153 : _GEN_7505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7507 = 10'h9a == _T_21 ? ram_154 : _GEN_7506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7508 = 10'h9b == _T_21 ? ram_155 : _GEN_7507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7509 = 10'h9c == _T_21 ? ram_156 : _GEN_7508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7510 = 10'h9d == _T_21 ? ram_157 : _GEN_7509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7511 = 10'h9e == _T_21 ? ram_158 : _GEN_7510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7512 = 10'h9f == _T_21 ? ram_159 : _GEN_7511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7513 = 10'ha0 == _T_21 ? ram_160 : _GEN_7512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7514 = 10'ha1 == _T_21 ? ram_161 : _GEN_7513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7515 = 10'ha2 == _T_21 ? ram_162 : _GEN_7514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7516 = 10'ha3 == _T_21 ? ram_163 : _GEN_7515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7517 = 10'ha4 == _T_21 ? ram_164 : _GEN_7516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7518 = 10'ha5 == _T_21 ? ram_165 : _GEN_7517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7519 = 10'ha6 == _T_21 ? ram_166 : _GEN_7518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7520 = 10'ha7 == _T_21 ? ram_167 : _GEN_7519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7521 = 10'ha8 == _T_21 ? ram_168 : _GEN_7520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7522 = 10'ha9 == _T_21 ? ram_169 : _GEN_7521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7523 = 10'haa == _T_21 ? ram_170 : _GEN_7522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7524 = 10'hab == _T_21 ? ram_171 : _GEN_7523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7525 = 10'hac == _T_21 ? ram_172 : _GEN_7524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7526 = 10'had == _T_21 ? ram_173 : _GEN_7525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7527 = 10'hae == _T_21 ? ram_174 : _GEN_7526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7528 = 10'haf == _T_21 ? ram_175 : _GEN_7527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7529 = 10'hb0 == _T_21 ? ram_176 : _GEN_7528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7530 = 10'hb1 == _T_21 ? ram_177 : _GEN_7529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7531 = 10'hb2 == _T_21 ? ram_178 : _GEN_7530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7532 = 10'hb3 == _T_21 ? ram_179 : _GEN_7531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7533 = 10'hb4 == _T_21 ? ram_180 : _GEN_7532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7534 = 10'hb5 == _T_21 ? ram_181 : _GEN_7533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7535 = 10'hb6 == _T_21 ? ram_182 : _GEN_7534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7536 = 10'hb7 == _T_21 ? ram_183 : _GEN_7535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7537 = 10'hb8 == _T_21 ? ram_184 : _GEN_7536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7538 = 10'hb9 == _T_21 ? ram_185 : _GEN_7537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7539 = 10'hba == _T_21 ? ram_186 : _GEN_7538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7540 = 10'hbb == _T_21 ? ram_187 : _GEN_7539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7541 = 10'hbc == _T_21 ? ram_188 : _GEN_7540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7542 = 10'hbd == _T_21 ? ram_189 : _GEN_7541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7543 = 10'hbe == _T_21 ? ram_190 : _GEN_7542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7544 = 10'hbf == _T_21 ? ram_191 : _GEN_7543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7545 = 10'hc0 == _T_21 ? ram_192 : _GEN_7544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7546 = 10'hc1 == _T_21 ? ram_193 : _GEN_7545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7547 = 10'hc2 == _T_21 ? ram_194 : _GEN_7546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7548 = 10'hc3 == _T_21 ? ram_195 : _GEN_7547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7549 = 10'hc4 == _T_21 ? ram_196 : _GEN_7548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7550 = 10'hc5 == _T_21 ? ram_197 : _GEN_7549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7551 = 10'hc6 == _T_21 ? ram_198 : _GEN_7550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7552 = 10'hc7 == _T_21 ? ram_199 : _GEN_7551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7553 = 10'hc8 == _T_21 ? ram_200 : _GEN_7552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7554 = 10'hc9 == _T_21 ? ram_201 : _GEN_7553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7555 = 10'hca == _T_21 ? ram_202 : _GEN_7554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7556 = 10'hcb == _T_21 ? ram_203 : _GEN_7555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7557 = 10'hcc == _T_21 ? ram_204 : _GEN_7556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7558 = 10'hcd == _T_21 ? ram_205 : _GEN_7557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7559 = 10'hce == _T_21 ? ram_206 : _GEN_7558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7560 = 10'hcf == _T_21 ? ram_207 : _GEN_7559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7561 = 10'hd0 == _T_21 ? ram_208 : _GEN_7560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7562 = 10'hd1 == _T_21 ? ram_209 : _GEN_7561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7563 = 10'hd2 == _T_21 ? ram_210 : _GEN_7562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7564 = 10'hd3 == _T_21 ? ram_211 : _GEN_7563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7565 = 10'hd4 == _T_21 ? ram_212 : _GEN_7564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7566 = 10'hd5 == _T_21 ? ram_213 : _GEN_7565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7567 = 10'hd6 == _T_21 ? ram_214 : _GEN_7566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7568 = 10'hd7 == _T_21 ? ram_215 : _GEN_7567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7569 = 10'hd8 == _T_21 ? ram_216 : _GEN_7568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7570 = 10'hd9 == _T_21 ? ram_217 : _GEN_7569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7571 = 10'hda == _T_21 ? ram_218 : _GEN_7570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7572 = 10'hdb == _T_21 ? ram_219 : _GEN_7571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7573 = 10'hdc == _T_21 ? ram_220 : _GEN_7572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7574 = 10'hdd == _T_21 ? ram_221 : _GEN_7573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7575 = 10'hde == _T_21 ? ram_222 : _GEN_7574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7576 = 10'hdf == _T_21 ? ram_223 : _GEN_7575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7577 = 10'he0 == _T_21 ? ram_224 : _GEN_7576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7578 = 10'he1 == _T_21 ? ram_225 : _GEN_7577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7579 = 10'he2 == _T_21 ? ram_226 : _GEN_7578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7580 = 10'he3 == _T_21 ? ram_227 : _GEN_7579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7581 = 10'he4 == _T_21 ? ram_228 : _GEN_7580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7582 = 10'he5 == _T_21 ? ram_229 : _GEN_7581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7583 = 10'he6 == _T_21 ? ram_230 : _GEN_7582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7584 = 10'he7 == _T_21 ? ram_231 : _GEN_7583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7585 = 10'he8 == _T_21 ? ram_232 : _GEN_7584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7586 = 10'he9 == _T_21 ? ram_233 : _GEN_7585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7587 = 10'hea == _T_21 ? ram_234 : _GEN_7586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7588 = 10'heb == _T_21 ? ram_235 : _GEN_7587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7589 = 10'hec == _T_21 ? ram_236 : _GEN_7588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7590 = 10'hed == _T_21 ? ram_237 : _GEN_7589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7591 = 10'hee == _T_21 ? ram_238 : _GEN_7590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7592 = 10'hef == _T_21 ? ram_239 : _GEN_7591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7593 = 10'hf0 == _T_21 ? ram_240 : _GEN_7592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7594 = 10'hf1 == _T_21 ? ram_241 : _GEN_7593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7595 = 10'hf2 == _T_21 ? ram_242 : _GEN_7594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7596 = 10'hf3 == _T_21 ? ram_243 : _GEN_7595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7597 = 10'hf4 == _T_21 ? ram_244 : _GEN_7596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7598 = 10'hf5 == _T_21 ? ram_245 : _GEN_7597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7599 = 10'hf6 == _T_21 ? ram_246 : _GEN_7598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7600 = 10'hf7 == _T_21 ? ram_247 : _GEN_7599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7601 = 10'hf8 == _T_21 ? ram_248 : _GEN_7600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7602 = 10'hf9 == _T_21 ? ram_249 : _GEN_7601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7603 = 10'hfa == _T_21 ? ram_250 : _GEN_7602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7604 = 10'hfb == _T_21 ? ram_251 : _GEN_7603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7605 = 10'hfc == _T_21 ? ram_252 : _GEN_7604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7606 = 10'hfd == _T_21 ? ram_253 : _GEN_7605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7607 = 10'hfe == _T_21 ? ram_254 : _GEN_7606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7608 = 10'hff == _T_21 ? ram_255 : _GEN_7607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7609 = 10'h100 == _T_21 ? ram_256 : _GEN_7608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7610 = 10'h101 == _T_21 ? ram_257 : _GEN_7609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7611 = 10'h102 == _T_21 ? ram_258 : _GEN_7610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7612 = 10'h103 == _T_21 ? ram_259 : _GEN_7611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7613 = 10'h104 == _T_21 ? ram_260 : _GEN_7612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7614 = 10'h105 == _T_21 ? ram_261 : _GEN_7613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7615 = 10'h106 == _T_21 ? ram_262 : _GEN_7614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7616 = 10'h107 == _T_21 ? ram_263 : _GEN_7615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7617 = 10'h108 == _T_21 ? ram_264 : _GEN_7616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7618 = 10'h109 == _T_21 ? ram_265 : _GEN_7617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7619 = 10'h10a == _T_21 ? ram_266 : _GEN_7618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7620 = 10'h10b == _T_21 ? ram_267 : _GEN_7619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7621 = 10'h10c == _T_21 ? ram_268 : _GEN_7620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7622 = 10'h10d == _T_21 ? ram_269 : _GEN_7621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7623 = 10'h10e == _T_21 ? ram_270 : _GEN_7622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7624 = 10'h10f == _T_21 ? ram_271 : _GEN_7623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7625 = 10'h110 == _T_21 ? ram_272 : _GEN_7624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7626 = 10'h111 == _T_21 ? ram_273 : _GEN_7625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7627 = 10'h112 == _T_21 ? ram_274 : _GEN_7626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7628 = 10'h113 == _T_21 ? ram_275 : _GEN_7627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7629 = 10'h114 == _T_21 ? ram_276 : _GEN_7628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7630 = 10'h115 == _T_21 ? ram_277 : _GEN_7629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7631 = 10'h116 == _T_21 ? ram_278 : _GEN_7630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7632 = 10'h117 == _T_21 ? ram_279 : _GEN_7631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7633 = 10'h118 == _T_21 ? ram_280 : _GEN_7632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7634 = 10'h119 == _T_21 ? ram_281 : _GEN_7633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7635 = 10'h11a == _T_21 ? ram_282 : _GEN_7634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7636 = 10'h11b == _T_21 ? ram_283 : _GEN_7635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7637 = 10'h11c == _T_21 ? ram_284 : _GEN_7636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7638 = 10'h11d == _T_21 ? ram_285 : _GEN_7637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7639 = 10'h11e == _T_21 ? ram_286 : _GEN_7638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7640 = 10'h11f == _T_21 ? ram_287 : _GEN_7639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7641 = 10'h120 == _T_21 ? ram_288 : _GEN_7640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7642 = 10'h121 == _T_21 ? ram_289 : _GEN_7641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7643 = 10'h122 == _T_21 ? ram_290 : _GEN_7642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7644 = 10'h123 == _T_21 ? ram_291 : _GEN_7643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7645 = 10'h124 == _T_21 ? ram_292 : _GEN_7644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7646 = 10'h125 == _T_21 ? ram_293 : _GEN_7645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7647 = 10'h126 == _T_21 ? ram_294 : _GEN_7646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7648 = 10'h127 == _T_21 ? ram_295 : _GEN_7647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7649 = 10'h128 == _T_21 ? ram_296 : _GEN_7648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7650 = 10'h129 == _T_21 ? ram_297 : _GEN_7649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7651 = 10'h12a == _T_21 ? ram_298 : _GEN_7650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7652 = 10'h12b == _T_21 ? ram_299 : _GEN_7651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7653 = 10'h12c == _T_21 ? ram_300 : _GEN_7652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7654 = 10'h12d == _T_21 ? ram_301 : _GEN_7653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7655 = 10'h12e == _T_21 ? ram_302 : _GEN_7654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7656 = 10'h12f == _T_21 ? ram_303 : _GEN_7655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7657 = 10'h130 == _T_21 ? ram_304 : _GEN_7656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7658 = 10'h131 == _T_21 ? ram_305 : _GEN_7657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7659 = 10'h132 == _T_21 ? ram_306 : _GEN_7658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7660 = 10'h133 == _T_21 ? ram_307 : _GEN_7659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7661 = 10'h134 == _T_21 ? ram_308 : _GEN_7660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7662 = 10'h135 == _T_21 ? ram_309 : _GEN_7661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7663 = 10'h136 == _T_21 ? ram_310 : _GEN_7662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7664 = 10'h137 == _T_21 ? ram_311 : _GEN_7663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7665 = 10'h138 == _T_21 ? ram_312 : _GEN_7664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7666 = 10'h139 == _T_21 ? ram_313 : _GEN_7665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7667 = 10'h13a == _T_21 ? ram_314 : _GEN_7666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7668 = 10'h13b == _T_21 ? ram_315 : _GEN_7667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7669 = 10'h13c == _T_21 ? ram_316 : _GEN_7668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7670 = 10'h13d == _T_21 ? ram_317 : _GEN_7669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7671 = 10'h13e == _T_21 ? ram_318 : _GEN_7670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7672 = 10'h13f == _T_21 ? ram_319 : _GEN_7671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7673 = 10'h140 == _T_21 ? ram_320 : _GEN_7672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7674 = 10'h141 == _T_21 ? ram_321 : _GEN_7673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7675 = 10'h142 == _T_21 ? ram_322 : _GEN_7674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7676 = 10'h143 == _T_21 ? ram_323 : _GEN_7675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7677 = 10'h144 == _T_21 ? ram_324 : _GEN_7676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7678 = 10'h145 == _T_21 ? ram_325 : _GEN_7677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7679 = 10'h146 == _T_21 ? ram_326 : _GEN_7678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7680 = 10'h147 == _T_21 ? ram_327 : _GEN_7679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7681 = 10'h148 == _T_21 ? ram_328 : _GEN_7680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7682 = 10'h149 == _T_21 ? ram_329 : _GEN_7681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7683 = 10'h14a == _T_21 ? ram_330 : _GEN_7682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7684 = 10'h14b == _T_21 ? ram_331 : _GEN_7683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7685 = 10'h14c == _T_21 ? ram_332 : _GEN_7684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7686 = 10'h14d == _T_21 ? ram_333 : _GEN_7685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7687 = 10'h14e == _T_21 ? ram_334 : _GEN_7686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7688 = 10'h14f == _T_21 ? ram_335 : _GEN_7687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7689 = 10'h150 == _T_21 ? ram_336 : _GEN_7688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7690 = 10'h151 == _T_21 ? ram_337 : _GEN_7689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7691 = 10'h152 == _T_21 ? ram_338 : _GEN_7690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7692 = 10'h153 == _T_21 ? ram_339 : _GEN_7691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7693 = 10'h154 == _T_21 ? ram_340 : _GEN_7692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7694 = 10'h155 == _T_21 ? ram_341 : _GEN_7693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7695 = 10'h156 == _T_21 ? ram_342 : _GEN_7694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7696 = 10'h157 == _T_21 ? ram_343 : _GEN_7695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7697 = 10'h158 == _T_21 ? ram_344 : _GEN_7696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7698 = 10'h159 == _T_21 ? ram_345 : _GEN_7697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7699 = 10'h15a == _T_21 ? ram_346 : _GEN_7698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7700 = 10'h15b == _T_21 ? ram_347 : _GEN_7699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7701 = 10'h15c == _T_21 ? ram_348 : _GEN_7700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7702 = 10'h15d == _T_21 ? ram_349 : _GEN_7701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7703 = 10'h15e == _T_21 ? ram_350 : _GEN_7702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7704 = 10'h15f == _T_21 ? ram_351 : _GEN_7703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7705 = 10'h160 == _T_21 ? ram_352 : _GEN_7704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7706 = 10'h161 == _T_21 ? ram_353 : _GEN_7705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7707 = 10'h162 == _T_21 ? ram_354 : _GEN_7706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7708 = 10'h163 == _T_21 ? ram_355 : _GEN_7707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7709 = 10'h164 == _T_21 ? ram_356 : _GEN_7708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7710 = 10'h165 == _T_21 ? ram_357 : _GEN_7709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7711 = 10'h166 == _T_21 ? ram_358 : _GEN_7710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7712 = 10'h167 == _T_21 ? ram_359 : _GEN_7711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7713 = 10'h168 == _T_21 ? ram_360 : _GEN_7712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7714 = 10'h169 == _T_21 ? ram_361 : _GEN_7713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7715 = 10'h16a == _T_21 ? ram_362 : _GEN_7714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7716 = 10'h16b == _T_21 ? ram_363 : _GEN_7715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7717 = 10'h16c == _T_21 ? ram_364 : _GEN_7716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7718 = 10'h16d == _T_21 ? ram_365 : _GEN_7717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7719 = 10'h16e == _T_21 ? ram_366 : _GEN_7718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7720 = 10'h16f == _T_21 ? ram_367 : _GEN_7719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7721 = 10'h170 == _T_21 ? ram_368 : _GEN_7720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7722 = 10'h171 == _T_21 ? ram_369 : _GEN_7721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7723 = 10'h172 == _T_21 ? ram_370 : _GEN_7722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7724 = 10'h173 == _T_21 ? ram_371 : _GEN_7723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7725 = 10'h174 == _T_21 ? ram_372 : _GEN_7724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7726 = 10'h175 == _T_21 ? ram_373 : _GEN_7725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7727 = 10'h176 == _T_21 ? ram_374 : _GEN_7726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7728 = 10'h177 == _T_21 ? ram_375 : _GEN_7727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7729 = 10'h178 == _T_21 ? ram_376 : _GEN_7728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7730 = 10'h179 == _T_21 ? ram_377 : _GEN_7729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7731 = 10'h17a == _T_21 ? ram_378 : _GEN_7730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7732 = 10'h17b == _T_21 ? ram_379 : _GEN_7731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7733 = 10'h17c == _T_21 ? ram_380 : _GEN_7732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7734 = 10'h17d == _T_21 ? ram_381 : _GEN_7733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7735 = 10'h17e == _T_21 ? ram_382 : _GEN_7734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7736 = 10'h17f == _T_21 ? ram_383 : _GEN_7735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7737 = 10'h180 == _T_21 ? ram_384 : _GEN_7736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7738 = 10'h181 == _T_21 ? ram_385 : _GEN_7737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7739 = 10'h182 == _T_21 ? ram_386 : _GEN_7738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7740 = 10'h183 == _T_21 ? ram_387 : _GEN_7739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7741 = 10'h184 == _T_21 ? ram_388 : _GEN_7740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7742 = 10'h185 == _T_21 ? ram_389 : _GEN_7741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7743 = 10'h186 == _T_21 ? ram_390 : _GEN_7742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7744 = 10'h187 == _T_21 ? ram_391 : _GEN_7743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7745 = 10'h188 == _T_21 ? ram_392 : _GEN_7744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7746 = 10'h189 == _T_21 ? ram_393 : _GEN_7745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7747 = 10'h18a == _T_21 ? ram_394 : _GEN_7746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7748 = 10'h18b == _T_21 ? ram_395 : _GEN_7747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7749 = 10'h18c == _T_21 ? ram_396 : _GEN_7748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7750 = 10'h18d == _T_21 ? ram_397 : _GEN_7749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7751 = 10'h18e == _T_21 ? ram_398 : _GEN_7750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7752 = 10'h18f == _T_21 ? ram_399 : _GEN_7751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7753 = 10'h190 == _T_21 ? ram_400 : _GEN_7752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7754 = 10'h191 == _T_21 ? ram_401 : _GEN_7753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7755 = 10'h192 == _T_21 ? ram_402 : _GEN_7754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7756 = 10'h193 == _T_21 ? ram_403 : _GEN_7755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7757 = 10'h194 == _T_21 ? ram_404 : _GEN_7756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7758 = 10'h195 == _T_21 ? ram_405 : _GEN_7757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7759 = 10'h196 == _T_21 ? ram_406 : _GEN_7758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7760 = 10'h197 == _T_21 ? ram_407 : _GEN_7759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7761 = 10'h198 == _T_21 ? ram_408 : _GEN_7760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7762 = 10'h199 == _T_21 ? ram_409 : _GEN_7761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7763 = 10'h19a == _T_21 ? ram_410 : _GEN_7762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7764 = 10'h19b == _T_21 ? ram_411 : _GEN_7763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7765 = 10'h19c == _T_21 ? ram_412 : _GEN_7764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7766 = 10'h19d == _T_21 ? ram_413 : _GEN_7765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7767 = 10'h19e == _T_21 ? ram_414 : _GEN_7766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7768 = 10'h19f == _T_21 ? ram_415 : _GEN_7767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7769 = 10'h1a0 == _T_21 ? ram_416 : _GEN_7768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7770 = 10'h1a1 == _T_21 ? ram_417 : _GEN_7769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7771 = 10'h1a2 == _T_21 ? ram_418 : _GEN_7770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7772 = 10'h1a3 == _T_21 ? ram_419 : _GEN_7771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7773 = 10'h1a4 == _T_21 ? ram_420 : _GEN_7772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7774 = 10'h1a5 == _T_21 ? ram_421 : _GEN_7773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7775 = 10'h1a6 == _T_21 ? ram_422 : _GEN_7774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7776 = 10'h1a7 == _T_21 ? ram_423 : _GEN_7775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7777 = 10'h1a8 == _T_21 ? ram_424 : _GEN_7776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7778 = 10'h1a9 == _T_21 ? ram_425 : _GEN_7777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7779 = 10'h1aa == _T_21 ? ram_426 : _GEN_7778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7780 = 10'h1ab == _T_21 ? ram_427 : _GEN_7779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7781 = 10'h1ac == _T_21 ? ram_428 : _GEN_7780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7782 = 10'h1ad == _T_21 ? ram_429 : _GEN_7781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7783 = 10'h1ae == _T_21 ? ram_430 : _GEN_7782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7784 = 10'h1af == _T_21 ? ram_431 : _GEN_7783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7785 = 10'h1b0 == _T_21 ? ram_432 : _GEN_7784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7786 = 10'h1b1 == _T_21 ? ram_433 : _GEN_7785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7787 = 10'h1b2 == _T_21 ? ram_434 : _GEN_7786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7788 = 10'h1b3 == _T_21 ? ram_435 : _GEN_7787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7789 = 10'h1b4 == _T_21 ? ram_436 : _GEN_7788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7790 = 10'h1b5 == _T_21 ? ram_437 : _GEN_7789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7791 = 10'h1b6 == _T_21 ? ram_438 : _GEN_7790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7792 = 10'h1b7 == _T_21 ? ram_439 : _GEN_7791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7793 = 10'h1b8 == _T_21 ? ram_440 : _GEN_7792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7794 = 10'h1b9 == _T_21 ? ram_441 : _GEN_7793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7795 = 10'h1ba == _T_21 ? ram_442 : _GEN_7794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7796 = 10'h1bb == _T_21 ? ram_443 : _GEN_7795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7797 = 10'h1bc == _T_21 ? ram_444 : _GEN_7796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7798 = 10'h1bd == _T_21 ? ram_445 : _GEN_7797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7799 = 10'h1be == _T_21 ? ram_446 : _GEN_7798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7800 = 10'h1bf == _T_21 ? ram_447 : _GEN_7799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7801 = 10'h1c0 == _T_21 ? ram_448 : _GEN_7800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7802 = 10'h1c1 == _T_21 ? ram_449 : _GEN_7801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7803 = 10'h1c2 == _T_21 ? ram_450 : _GEN_7802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7804 = 10'h1c3 == _T_21 ? ram_451 : _GEN_7803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7805 = 10'h1c4 == _T_21 ? ram_452 : _GEN_7804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7806 = 10'h1c5 == _T_21 ? ram_453 : _GEN_7805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7807 = 10'h1c6 == _T_21 ? ram_454 : _GEN_7806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7808 = 10'h1c7 == _T_21 ? ram_455 : _GEN_7807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7809 = 10'h1c8 == _T_21 ? ram_456 : _GEN_7808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7810 = 10'h1c9 == _T_21 ? ram_457 : _GEN_7809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7811 = 10'h1ca == _T_21 ? ram_458 : _GEN_7810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7812 = 10'h1cb == _T_21 ? ram_459 : _GEN_7811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7813 = 10'h1cc == _T_21 ? ram_460 : _GEN_7812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7814 = 10'h1cd == _T_21 ? ram_461 : _GEN_7813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7815 = 10'h1ce == _T_21 ? ram_462 : _GEN_7814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7816 = 10'h1cf == _T_21 ? ram_463 : _GEN_7815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7817 = 10'h1d0 == _T_21 ? ram_464 : _GEN_7816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7818 = 10'h1d1 == _T_21 ? ram_465 : _GEN_7817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7819 = 10'h1d2 == _T_21 ? ram_466 : _GEN_7818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7820 = 10'h1d3 == _T_21 ? ram_467 : _GEN_7819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7821 = 10'h1d4 == _T_21 ? ram_468 : _GEN_7820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7822 = 10'h1d5 == _T_21 ? ram_469 : _GEN_7821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7823 = 10'h1d6 == _T_21 ? ram_470 : _GEN_7822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7824 = 10'h1d7 == _T_21 ? ram_471 : _GEN_7823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7825 = 10'h1d8 == _T_21 ? ram_472 : _GEN_7824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7826 = 10'h1d9 == _T_21 ? ram_473 : _GEN_7825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7827 = 10'h1da == _T_21 ? ram_474 : _GEN_7826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7828 = 10'h1db == _T_21 ? ram_475 : _GEN_7827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7829 = 10'h1dc == _T_21 ? ram_476 : _GEN_7828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7830 = 10'h1dd == _T_21 ? ram_477 : _GEN_7829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7831 = 10'h1de == _T_21 ? ram_478 : _GEN_7830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7832 = 10'h1df == _T_21 ? ram_479 : _GEN_7831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7833 = 10'h1e0 == _T_21 ? ram_480 : _GEN_7832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7834 = 10'h1e1 == _T_21 ? ram_481 : _GEN_7833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7835 = 10'h1e2 == _T_21 ? ram_482 : _GEN_7834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7836 = 10'h1e3 == _T_21 ? ram_483 : _GEN_7835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7837 = 10'h1e4 == _T_21 ? ram_484 : _GEN_7836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7838 = 10'h1e5 == _T_21 ? ram_485 : _GEN_7837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7839 = 10'h1e6 == _T_21 ? ram_486 : _GEN_7838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7840 = 10'h1e7 == _T_21 ? ram_487 : _GEN_7839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7841 = 10'h1e8 == _T_21 ? ram_488 : _GEN_7840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7842 = 10'h1e9 == _T_21 ? ram_489 : _GEN_7841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7843 = 10'h1ea == _T_21 ? ram_490 : _GEN_7842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7844 = 10'h1eb == _T_21 ? ram_491 : _GEN_7843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7845 = 10'h1ec == _T_21 ? ram_492 : _GEN_7844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7846 = 10'h1ed == _T_21 ? ram_493 : _GEN_7845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7847 = 10'h1ee == _T_21 ? ram_494 : _GEN_7846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7848 = 10'h1ef == _T_21 ? ram_495 : _GEN_7847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7849 = 10'h1f0 == _T_21 ? ram_496 : _GEN_7848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7850 = 10'h1f1 == _T_21 ? ram_497 : _GEN_7849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7851 = 10'h1f2 == _T_21 ? ram_498 : _GEN_7850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7852 = 10'h1f3 == _T_21 ? ram_499 : _GEN_7851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7853 = 10'h1f4 == _T_21 ? ram_500 : _GEN_7852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7854 = 10'h1f5 == _T_21 ? ram_501 : _GEN_7853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7855 = 10'h1f6 == _T_21 ? ram_502 : _GEN_7854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7856 = 10'h1f7 == _T_21 ? ram_503 : _GEN_7855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7857 = 10'h1f8 == _T_21 ? ram_504 : _GEN_7856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7858 = 10'h1f9 == _T_21 ? ram_505 : _GEN_7857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7859 = 10'h1fa == _T_21 ? ram_506 : _GEN_7858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7860 = 10'h1fb == _T_21 ? ram_507 : _GEN_7859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7861 = 10'h1fc == _T_21 ? ram_508 : _GEN_7860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7862 = 10'h1fd == _T_21 ? ram_509 : _GEN_7861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7863 = 10'h1fe == _T_21 ? ram_510 : _GEN_7862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7864 = 10'h1ff == _T_21 ? ram_511 : _GEN_7863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7865 = 10'h200 == _T_21 ? ram_512 : _GEN_7864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7866 = 10'h201 == _T_21 ? ram_513 : _GEN_7865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7867 = 10'h202 == _T_21 ? ram_514 : _GEN_7866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7868 = 10'h203 == _T_21 ? ram_515 : _GEN_7867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7869 = 10'h204 == _T_21 ? ram_516 : _GEN_7868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7870 = 10'h205 == _T_21 ? ram_517 : _GEN_7869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7871 = 10'h206 == _T_21 ? ram_518 : _GEN_7870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7872 = 10'h207 == _T_21 ? ram_519 : _GEN_7871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7873 = 10'h208 == _T_21 ? ram_520 : _GEN_7872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7874 = 10'h209 == _T_21 ? ram_521 : _GEN_7873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7875 = 10'h20a == _T_21 ? ram_522 : _GEN_7874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7876 = 10'h20b == _T_21 ? ram_523 : _GEN_7875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_7877 = 10'h20c == _T_21 ? ram_524 : _GEN_7876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19075 = {{8190'd0}, _GEN_7877}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_207 = _GEN_19075 ^ _ram_T_206; // @[vga.scala 64:41]
  wire [287:0] _GEN_7878 = 10'h0 == _T_21 ? _ram_T_207[287:0] : _GEN_6828; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7879 = 10'h1 == _T_21 ? _ram_T_207[287:0] : _GEN_6829; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7880 = 10'h2 == _T_21 ? _ram_T_207[287:0] : _GEN_6830; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7881 = 10'h3 == _T_21 ? _ram_T_207[287:0] : _GEN_6831; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7882 = 10'h4 == _T_21 ? _ram_T_207[287:0] : _GEN_6832; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7883 = 10'h5 == _T_21 ? _ram_T_207[287:0] : _GEN_6833; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7884 = 10'h6 == _T_21 ? _ram_T_207[287:0] : _GEN_6834; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7885 = 10'h7 == _T_21 ? _ram_T_207[287:0] : _GEN_6835; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7886 = 10'h8 == _T_21 ? _ram_T_207[287:0] : _GEN_6836; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7887 = 10'h9 == _T_21 ? _ram_T_207[287:0] : _GEN_6837; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7888 = 10'ha == _T_21 ? _ram_T_207[287:0] : _GEN_6838; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7889 = 10'hb == _T_21 ? _ram_T_207[287:0] : _GEN_6839; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7890 = 10'hc == _T_21 ? _ram_T_207[287:0] : _GEN_6840; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7891 = 10'hd == _T_21 ? _ram_T_207[287:0] : _GEN_6841; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7892 = 10'he == _T_21 ? _ram_T_207[287:0] : _GEN_6842; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7893 = 10'hf == _T_21 ? _ram_T_207[287:0] : _GEN_6843; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7894 = 10'h10 == _T_21 ? _ram_T_207[287:0] : _GEN_6844; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7895 = 10'h11 == _T_21 ? _ram_T_207[287:0] : _GEN_6845; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7896 = 10'h12 == _T_21 ? _ram_T_207[287:0] : _GEN_6846; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7897 = 10'h13 == _T_21 ? _ram_T_207[287:0] : _GEN_6847; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7898 = 10'h14 == _T_21 ? _ram_T_207[287:0] : _GEN_6848; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7899 = 10'h15 == _T_21 ? _ram_T_207[287:0] : _GEN_6849; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7900 = 10'h16 == _T_21 ? _ram_T_207[287:0] : _GEN_6850; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7901 = 10'h17 == _T_21 ? _ram_T_207[287:0] : _GEN_6851; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7902 = 10'h18 == _T_21 ? _ram_T_207[287:0] : _GEN_6852; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7903 = 10'h19 == _T_21 ? _ram_T_207[287:0] : _GEN_6853; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7904 = 10'h1a == _T_21 ? _ram_T_207[287:0] : _GEN_6854; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7905 = 10'h1b == _T_21 ? _ram_T_207[287:0] : _GEN_6855; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7906 = 10'h1c == _T_21 ? _ram_T_207[287:0] : _GEN_6856; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7907 = 10'h1d == _T_21 ? _ram_T_207[287:0] : _GEN_6857; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7908 = 10'h1e == _T_21 ? _ram_T_207[287:0] : _GEN_6858; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7909 = 10'h1f == _T_21 ? _ram_T_207[287:0] : _GEN_6859; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7910 = 10'h20 == _T_21 ? _ram_T_207[287:0] : _GEN_6860; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7911 = 10'h21 == _T_21 ? _ram_T_207[287:0] : _GEN_6861; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7912 = 10'h22 == _T_21 ? _ram_T_207[287:0] : _GEN_6862; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7913 = 10'h23 == _T_21 ? _ram_T_207[287:0] : _GEN_6863; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7914 = 10'h24 == _T_21 ? _ram_T_207[287:0] : _GEN_6864; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7915 = 10'h25 == _T_21 ? _ram_T_207[287:0] : _GEN_6865; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7916 = 10'h26 == _T_21 ? _ram_T_207[287:0] : _GEN_6866; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7917 = 10'h27 == _T_21 ? _ram_T_207[287:0] : _GEN_6867; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7918 = 10'h28 == _T_21 ? _ram_T_207[287:0] : _GEN_6868; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7919 = 10'h29 == _T_21 ? _ram_T_207[287:0] : _GEN_6869; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7920 = 10'h2a == _T_21 ? _ram_T_207[287:0] : _GEN_6870; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7921 = 10'h2b == _T_21 ? _ram_T_207[287:0] : _GEN_6871; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7922 = 10'h2c == _T_21 ? _ram_T_207[287:0] : _GEN_6872; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7923 = 10'h2d == _T_21 ? _ram_T_207[287:0] : _GEN_6873; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7924 = 10'h2e == _T_21 ? _ram_T_207[287:0] : _GEN_6874; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7925 = 10'h2f == _T_21 ? _ram_T_207[287:0] : _GEN_6875; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7926 = 10'h30 == _T_21 ? _ram_T_207[287:0] : _GEN_6876; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7927 = 10'h31 == _T_21 ? _ram_T_207[287:0] : _GEN_6877; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7928 = 10'h32 == _T_21 ? _ram_T_207[287:0] : _GEN_6878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7929 = 10'h33 == _T_21 ? _ram_T_207[287:0] : _GEN_6879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7930 = 10'h34 == _T_21 ? _ram_T_207[287:0] : _GEN_6880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7931 = 10'h35 == _T_21 ? _ram_T_207[287:0] : _GEN_6881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7932 = 10'h36 == _T_21 ? _ram_T_207[287:0] : _GEN_6882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7933 = 10'h37 == _T_21 ? _ram_T_207[287:0] : _GEN_6883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7934 = 10'h38 == _T_21 ? _ram_T_207[287:0] : _GEN_6884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7935 = 10'h39 == _T_21 ? _ram_T_207[287:0] : _GEN_6885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7936 = 10'h3a == _T_21 ? _ram_T_207[287:0] : _GEN_6886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7937 = 10'h3b == _T_21 ? _ram_T_207[287:0] : _GEN_6887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7938 = 10'h3c == _T_21 ? _ram_T_207[287:0] : _GEN_6888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7939 = 10'h3d == _T_21 ? _ram_T_207[287:0] : _GEN_6889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7940 = 10'h3e == _T_21 ? _ram_T_207[287:0] : _GEN_6890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7941 = 10'h3f == _T_21 ? _ram_T_207[287:0] : _GEN_6891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7942 = 10'h40 == _T_21 ? _ram_T_207[287:0] : _GEN_6892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7943 = 10'h41 == _T_21 ? _ram_T_207[287:0] : _GEN_6893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7944 = 10'h42 == _T_21 ? _ram_T_207[287:0] : _GEN_6894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7945 = 10'h43 == _T_21 ? _ram_T_207[287:0] : _GEN_6895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7946 = 10'h44 == _T_21 ? _ram_T_207[287:0] : _GEN_6896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7947 = 10'h45 == _T_21 ? _ram_T_207[287:0] : _GEN_6897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7948 = 10'h46 == _T_21 ? _ram_T_207[287:0] : _GEN_6898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7949 = 10'h47 == _T_21 ? _ram_T_207[287:0] : _GEN_6899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7950 = 10'h48 == _T_21 ? _ram_T_207[287:0] : _GEN_6900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7951 = 10'h49 == _T_21 ? _ram_T_207[287:0] : _GEN_6901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7952 = 10'h4a == _T_21 ? _ram_T_207[287:0] : _GEN_6902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7953 = 10'h4b == _T_21 ? _ram_T_207[287:0] : _GEN_6903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7954 = 10'h4c == _T_21 ? _ram_T_207[287:0] : _GEN_6904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7955 = 10'h4d == _T_21 ? _ram_T_207[287:0] : _GEN_6905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7956 = 10'h4e == _T_21 ? _ram_T_207[287:0] : _GEN_6906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7957 = 10'h4f == _T_21 ? _ram_T_207[287:0] : _GEN_6907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7958 = 10'h50 == _T_21 ? _ram_T_207[287:0] : _GEN_6908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7959 = 10'h51 == _T_21 ? _ram_T_207[287:0] : _GEN_6909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7960 = 10'h52 == _T_21 ? _ram_T_207[287:0] : _GEN_6910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7961 = 10'h53 == _T_21 ? _ram_T_207[287:0] : _GEN_6911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7962 = 10'h54 == _T_21 ? _ram_T_207[287:0] : _GEN_6912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7963 = 10'h55 == _T_21 ? _ram_T_207[287:0] : _GEN_6913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7964 = 10'h56 == _T_21 ? _ram_T_207[287:0] : _GEN_6914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7965 = 10'h57 == _T_21 ? _ram_T_207[287:0] : _GEN_6915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7966 = 10'h58 == _T_21 ? _ram_T_207[287:0] : _GEN_6916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7967 = 10'h59 == _T_21 ? _ram_T_207[287:0] : _GEN_6917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7968 = 10'h5a == _T_21 ? _ram_T_207[287:0] : _GEN_6918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7969 = 10'h5b == _T_21 ? _ram_T_207[287:0] : _GEN_6919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7970 = 10'h5c == _T_21 ? _ram_T_207[287:0] : _GEN_6920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7971 = 10'h5d == _T_21 ? _ram_T_207[287:0] : _GEN_6921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7972 = 10'h5e == _T_21 ? _ram_T_207[287:0] : _GEN_6922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7973 = 10'h5f == _T_21 ? _ram_T_207[287:0] : _GEN_6923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7974 = 10'h60 == _T_21 ? _ram_T_207[287:0] : _GEN_6924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7975 = 10'h61 == _T_21 ? _ram_T_207[287:0] : _GEN_6925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7976 = 10'h62 == _T_21 ? _ram_T_207[287:0] : _GEN_6926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7977 = 10'h63 == _T_21 ? _ram_T_207[287:0] : _GEN_6927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7978 = 10'h64 == _T_21 ? _ram_T_207[287:0] : _GEN_6928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7979 = 10'h65 == _T_21 ? _ram_T_207[287:0] : _GEN_6929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7980 = 10'h66 == _T_21 ? _ram_T_207[287:0] : _GEN_6930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7981 = 10'h67 == _T_21 ? _ram_T_207[287:0] : _GEN_6931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7982 = 10'h68 == _T_21 ? _ram_T_207[287:0] : _GEN_6932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7983 = 10'h69 == _T_21 ? _ram_T_207[287:0] : _GEN_6933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7984 = 10'h6a == _T_21 ? _ram_T_207[287:0] : _GEN_6934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7985 = 10'h6b == _T_21 ? _ram_T_207[287:0] : _GEN_6935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7986 = 10'h6c == _T_21 ? _ram_T_207[287:0] : _GEN_6936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7987 = 10'h6d == _T_21 ? _ram_T_207[287:0] : _GEN_6937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7988 = 10'h6e == _T_21 ? _ram_T_207[287:0] : _GEN_6938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7989 = 10'h6f == _T_21 ? _ram_T_207[287:0] : _GEN_6939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7990 = 10'h70 == _T_21 ? _ram_T_207[287:0] : _GEN_6940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7991 = 10'h71 == _T_21 ? _ram_T_207[287:0] : _GEN_6941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7992 = 10'h72 == _T_21 ? _ram_T_207[287:0] : _GEN_6942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7993 = 10'h73 == _T_21 ? _ram_T_207[287:0] : _GEN_6943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7994 = 10'h74 == _T_21 ? _ram_T_207[287:0] : _GEN_6944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7995 = 10'h75 == _T_21 ? _ram_T_207[287:0] : _GEN_6945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7996 = 10'h76 == _T_21 ? _ram_T_207[287:0] : _GEN_6946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7997 = 10'h77 == _T_21 ? _ram_T_207[287:0] : _GEN_6947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7998 = 10'h78 == _T_21 ? _ram_T_207[287:0] : _GEN_6948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_7999 = 10'h79 == _T_21 ? _ram_T_207[287:0] : _GEN_6949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8000 = 10'h7a == _T_21 ? _ram_T_207[287:0] : _GEN_6950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8001 = 10'h7b == _T_21 ? _ram_T_207[287:0] : _GEN_6951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8002 = 10'h7c == _T_21 ? _ram_T_207[287:0] : _GEN_6952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8003 = 10'h7d == _T_21 ? _ram_T_207[287:0] : _GEN_6953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8004 = 10'h7e == _T_21 ? _ram_T_207[287:0] : _GEN_6954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8005 = 10'h7f == _T_21 ? _ram_T_207[287:0] : _GEN_6955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8006 = 10'h80 == _T_21 ? _ram_T_207[287:0] : _GEN_6956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8007 = 10'h81 == _T_21 ? _ram_T_207[287:0] : _GEN_6957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8008 = 10'h82 == _T_21 ? _ram_T_207[287:0] : _GEN_6958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8009 = 10'h83 == _T_21 ? _ram_T_207[287:0] : _GEN_6959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8010 = 10'h84 == _T_21 ? _ram_T_207[287:0] : _GEN_6960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8011 = 10'h85 == _T_21 ? _ram_T_207[287:0] : _GEN_6961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8012 = 10'h86 == _T_21 ? _ram_T_207[287:0] : _GEN_6962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8013 = 10'h87 == _T_21 ? _ram_T_207[287:0] : _GEN_6963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8014 = 10'h88 == _T_21 ? _ram_T_207[287:0] : _GEN_6964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8015 = 10'h89 == _T_21 ? _ram_T_207[287:0] : _GEN_6965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8016 = 10'h8a == _T_21 ? _ram_T_207[287:0] : _GEN_6966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8017 = 10'h8b == _T_21 ? _ram_T_207[287:0] : _GEN_6967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8018 = 10'h8c == _T_21 ? _ram_T_207[287:0] : _GEN_6968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8019 = 10'h8d == _T_21 ? _ram_T_207[287:0] : _GEN_6969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8020 = 10'h8e == _T_21 ? _ram_T_207[287:0] : _GEN_6970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8021 = 10'h8f == _T_21 ? _ram_T_207[287:0] : _GEN_6971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8022 = 10'h90 == _T_21 ? _ram_T_207[287:0] : _GEN_6972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8023 = 10'h91 == _T_21 ? _ram_T_207[287:0] : _GEN_6973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8024 = 10'h92 == _T_21 ? _ram_T_207[287:0] : _GEN_6974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8025 = 10'h93 == _T_21 ? _ram_T_207[287:0] : _GEN_6975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8026 = 10'h94 == _T_21 ? _ram_T_207[287:0] : _GEN_6976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8027 = 10'h95 == _T_21 ? _ram_T_207[287:0] : _GEN_6977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8028 = 10'h96 == _T_21 ? _ram_T_207[287:0] : _GEN_6978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8029 = 10'h97 == _T_21 ? _ram_T_207[287:0] : _GEN_6979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8030 = 10'h98 == _T_21 ? _ram_T_207[287:0] : _GEN_6980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8031 = 10'h99 == _T_21 ? _ram_T_207[287:0] : _GEN_6981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8032 = 10'h9a == _T_21 ? _ram_T_207[287:0] : _GEN_6982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8033 = 10'h9b == _T_21 ? _ram_T_207[287:0] : _GEN_6983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8034 = 10'h9c == _T_21 ? _ram_T_207[287:0] : _GEN_6984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8035 = 10'h9d == _T_21 ? _ram_T_207[287:0] : _GEN_6985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8036 = 10'h9e == _T_21 ? _ram_T_207[287:0] : _GEN_6986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8037 = 10'h9f == _T_21 ? _ram_T_207[287:0] : _GEN_6987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8038 = 10'ha0 == _T_21 ? _ram_T_207[287:0] : _GEN_6988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8039 = 10'ha1 == _T_21 ? _ram_T_207[287:0] : _GEN_6989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8040 = 10'ha2 == _T_21 ? _ram_T_207[287:0] : _GEN_6990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8041 = 10'ha3 == _T_21 ? _ram_T_207[287:0] : _GEN_6991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8042 = 10'ha4 == _T_21 ? _ram_T_207[287:0] : _GEN_6992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8043 = 10'ha5 == _T_21 ? _ram_T_207[287:0] : _GEN_6993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8044 = 10'ha6 == _T_21 ? _ram_T_207[287:0] : _GEN_6994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8045 = 10'ha7 == _T_21 ? _ram_T_207[287:0] : _GEN_6995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8046 = 10'ha8 == _T_21 ? _ram_T_207[287:0] : _GEN_6996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8047 = 10'ha9 == _T_21 ? _ram_T_207[287:0] : _GEN_6997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8048 = 10'haa == _T_21 ? _ram_T_207[287:0] : _GEN_6998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8049 = 10'hab == _T_21 ? _ram_T_207[287:0] : _GEN_6999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8050 = 10'hac == _T_21 ? _ram_T_207[287:0] : _GEN_7000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8051 = 10'had == _T_21 ? _ram_T_207[287:0] : _GEN_7001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8052 = 10'hae == _T_21 ? _ram_T_207[287:0] : _GEN_7002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8053 = 10'haf == _T_21 ? _ram_T_207[287:0] : _GEN_7003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8054 = 10'hb0 == _T_21 ? _ram_T_207[287:0] : _GEN_7004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8055 = 10'hb1 == _T_21 ? _ram_T_207[287:0] : _GEN_7005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8056 = 10'hb2 == _T_21 ? _ram_T_207[287:0] : _GEN_7006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8057 = 10'hb3 == _T_21 ? _ram_T_207[287:0] : _GEN_7007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8058 = 10'hb4 == _T_21 ? _ram_T_207[287:0] : _GEN_7008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8059 = 10'hb5 == _T_21 ? _ram_T_207[287:0] : _GEN_7009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8060 = 10'hb6 == _T_21 ? _ram_T_207[287:0] : _GEN_7010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8061 = 10'hb7 == _T_21 ? _ram_T_207[287:0] : _GEN_7011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8062 = 10'hb8 == _T_21 ? _ram_T_207[287:0] : _GEN_7012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8063 = 10'hb9 == _T_21 ? _ram_T_207[287:0] : _GEN_7013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8064 = 10'hba == _T_21 ? _ram_T_207[287:0] : _GEN_7014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8065 = 10'hbb == _T_21 ? _ram_T_207[287:0] : _GEN_7015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8066 = 10'hbc == _T_21 ? _ram_T_207[287:0] : _GEN_7016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8067 = 10'hbd == _T_21 ? _ram_T_207[287:0] : _GEN_7017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8068 = 10'hbe == _T_21 ? _ram_T_207[287:0] : _GEN_7018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8069 = 10'hbf == _T_21 ? _ram_T_207[287:0] : _GEN_7019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8070 = 10'hc0 == _T_21 ? _ram_T_207[287:0] : _GEN_7020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8071 = 10'hc1 == _T_21 ? _ram_T_207[287:0] : _GEN_7021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8072 = 10'hc2 == _T_21 ? _ram_T_207[287:0] : _GEN_7022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8073 = 10'hc3 == _T_21 ? _ram_T_207[287:0] : _GEN_7023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8074 = 10'hc4 == _T_21 ? _ram_T_207[287:0] : _GEN_7024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8075 = 10'hc5 == _T_21 ? _ram_T_207[287:0] : _GEN_7025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8076 = 10'hc6 == _T_21 ? _ram_T_207[287:0] : _GEN_7026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8077 = 10'hc7 == _T_21 ? _ram_T_207[287:0] : _GEN_7027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8078 = 10'hc8 == _T_21 ? _ram_T_207[287:0] : _GEN_7028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8079 = 10'hc9 == _T_21 ? _ram_T_207[287:0] : _GEN_7029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8080 = 10'hca == _T_21 ? _ram_T_207[287:0] : _GEN_7030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8081 = 10'hcb == _T_21 ? _ram_T_207[287:0] : _GEN_7031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8082 = 10'hcc == _T_21 ? _ram_T_207[287:0] : _GEN_7032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8083 = 10'hcd == _T_21 ? _ram_T_207[287:0] : _GEN_7033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8084 = 10'hce == _T_21 ? _ram_T_207[287:0] : _GEN_7034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8085 = 10'hcf == _T_21 ? _ram_T_207[287:0] : _GEN_7035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8086 = 10'hd0 == _T_21 ? _ram_T_207[287:0] : _GEN_7036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8087 = 10'hd1 == _T_21 ? _ram_T_207[287:0] : _GEN_7037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8088 = 10'hd2 == _T_21 ? _ram_T_207[287:0] : _GEN_7038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8089 = 10'hd3 == _T_21 ? _ram_T_207[287:0] : _GEN_7039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8090 = 10'hd4 == _T_21 ? _ram_T_207[287:0] : _GEN_7040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8091 = 10'hd5 == _T_21 ? _ram_T_207[287:0] : _GEN_7041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8092 = 10'hd6 == _T_21 ? _ram_T_207[287:0] : _GEN_7042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8093 = 10'hd7 == _T_21 ? _ram_T_207[287:0] : _GEN_7043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8094 = 10'hd8 == _T_21 ? _ram_T_207[287:0] : _GEN_7044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8095 = 10'hd9 == _T_21 ? _ram_T_207[287:0] : _GEN_7045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8096 = 10'hda == _T_21 ? _ram_T_207[287:0] : _GEN_7046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8097 = 10'hdb == _T_21 ? _ram_T_207[287:0] : _GEN_7047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8098 = 10'hdc == _T_21 ? _ram_T_207[287:0] : _GEN_7048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8099 = 10'hdd == _T_21 ? _ram_T_207[287:0] : _GEN_7049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8100 = 10'hde == _T_21 ? _ram_T_207[287:0] : _GEN_7050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8101 = 10'hdf == _T_21 ? _ram_T_207[287:0] : _GEN_7051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8102 = 10'he0 == _T_21 ? _ram_T_207[287:0] : _GEN_7052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8103 = 10'he1 == _T_21 ? _ram_T_207[287:0] : _GEN_7053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8104 = 10'he2 == _T_21 ? _ram_T_207[287:0] : _GEN_7054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8105 = 10'he3 == _T_21 ? _ram_T_207[287:0] : _GEN_7055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8106 = 10'he4 == _T_21 ? _ram_T_207[287:0] : _GEN_7056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8107 = 10'he5 == _T_21 ? _ram_T_207[287:0] : _GEN_7057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8108 = 10'he6 == _T_21 ? _ram_T_207[287:0] : _GEN_7058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8109 = 10'he7 == _T_21 ? _ram_T_207[287:0] : _GEN_7059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8110 = 10'he8 == _T_21 ? _ram_T_207[287:0] : _GEN_7060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8111 = 10'he9 == _T_21 ? _ram_T_207[287:0] : _GEN_7061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8112 = 10'hea == _T_21 ? _ram_T_207[287:0] : _GEN_7062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8113 = 10'heb == _T_21 ? _ram_T_207[287:0] : _GEN_7063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8114 = 10'hec == _T_21 ? _ram_T_207[287:0] : _GEN_7064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8115 = 10'hed == _T_21 ? _ram_T_207[287:0] : _GEN_7065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8116 = 10'hee == _T_21 ? _ram_T_207[287:0] : _GEN_7066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8117 = 10'hef == _T_21 ? _ram_T_207[287:0] : _GEN_7067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8118 = 10'hf0 == _T_21 ? _ram_T_207[287:0] : _GEN_7068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8119 = 10'hf1 == _T_21 ? _ram_T_207[287:0] : _GEN_7069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8120 = 10'hf2 == _T_21 ? _ram_T_207[287:0] : _GEN_7070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8121 = 10'hf3 == _T_21 ? _ram_T_207[287:0] : _GEN_7071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8122 = 10'hf4 == _T_21 ? _ram_T_207[287:0] : _GEN_7072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8123 = 10'hf5 == _T_21 ? _ram_T_207[287:0] : _GEN_7073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8124 = 10'hf6 == _T_21 ? _ram_T_207[287:0] : _GEN_7074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8125 = 10'hf7 == _T_21 ? _ram_T_207[287:0] : _GEN_7075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8126 = 10'hf8 == _T_21 ? _ram_T_207[287:0] : _GEN_7076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8127 = 10'hf9 == _T_21 ? _ram_T_207[287:0] : _GEN_7077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8128 = 10'hfa == _T_21 ? _ram_T_207[287:0] : _GEN_7078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8129 = 10'hfb == _T_21 ? _ram_T_207[287:0] : _GEN_7079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8130 = 10'hfc == _T_21 ? _ram_T_207[287:0] : _GEN_7080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8131 = 10'hfd == _T_21 ? _ram_T_207[287:0] : _GEN_7081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8132 = 10'hfe == _T_21 ? _ram_T_207[287:0] : _GEN_7082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8133 = 10'hff == _T_21 ? _ram_T_207[287:0] : _GEN_7083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8134 = 10'h100 == _T_21 ? _ram_T_207[287:0] : _GEN_7084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8135 = 10'h101 == _T_21 ? _ram_T_207[287:0] : _GEN_7085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8136 = 10'h102 == _T_21 ? _ram_T_207[287:0] : _GEN_7086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8137 = 10'h103 == _T_21 ? _ram_T_207[287:0] : _GEN_7087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8138 = 10'h104 == _T_21 ? _ram_T_207[287:0] : _GEN_7088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8139 = 10'h105 == _T_21 ? _ram_T_207[287:0] : _GEN_7089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8140 = 10'h106 == _T_21 ? _ram_T_207[287:0] : _GEN_7090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8141 = 10'h107 == _T_21 ? _ram_T_207[287:0] : _GEN_7091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8142 = 10'h108 == _T_21 ? _ram_T_207[287:0] : _GEN_7092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8143 = 10'h109 == _T_21 ? _ram_T_207[287:0] : _GEN_7093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8144 = 10'h10a == _T_21 ? _ram_T_207[287:0] : _GEN_7094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8145 = 10'h10b == _T_21 ? _ram_T_207[287:0] : _GEN_7095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8146 = 10'h10c == _T_21 ? _ram_T_207[287:0] : _GEN_7096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8147 = 10'h10d == _T_21 ? _ram_T_207[287:0] : _GEN_7097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8148 = 10'h10e == _T_21 ? _ram_T_207[287:0] : _GEN_7098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8149 = 10'h10f == _T_21 ? _ram_T_207[287:0] : _GEN_7099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8150 = 10'h110 == _T_21 ? _ram_T_207[287:0] : _GEN_7100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8151 = 10'h111 == _T_21 ? _ram_T_207[287:0] : _GEN_7101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8152 = 10'h112 == _T_21 ? _ram_T_207[287:0] : _GEN_7102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8153 = 10'h113 == _T_21 ? _ram_T_207[287:0] : _GEN_7103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8154 = 10'h114 == _T_21 ? _ram_T_207[287:0] : _GEN_7104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8155 = 10'h115 == _T_21 ? _ram_T_207[287:0] : _GEN_7105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8156 = 10'h116 == _T_21 ? _ram_T_207[287:0] : _GEN_7106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8157 = 10'h117 == _T_21 ? _ram_T_207[287:0] : _GEN_7107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8158 = 10'h118 == _T_21 ? _ram_T_207[287:0] : _GEN_7108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8159 = 10'h119 == _T_21 ? _ram_T_207[287:0] : _GEN_7109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8160 = 10'h11a == _T_21 ? _ram_T_207[287:0] : _GEN_7110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8161 = 10'h11b == _T_21 ? _ram_T_207[287:0] : _GEN_7111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8162 = 10'h11c == _T_21 ? _ram_T_207[287:0] : _GEN_7112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8163 = 10'h11d == _T_21 ? _ram_T_207[287:0] : _GEN_7113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8164 = 10'h11e == _T_21 ? _ram_T_207[287:0] : _GEN_7114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8165 = 10'h11f == _T_21 ? _ram_T_207[287:0] : _GEN_7115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8166 = 10'h120 == _T_21 ? _ram_T_207[287:0] : _GEN_7116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8167 = 10'h121 == _T_21 ? _ram_T_207[287:0] : _GEN_7117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8168 = 10'h122 == _T_21 ? _ram_T_207[287:0] : _GEN_7118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8169 = 10'h123 == _T_21 ? _ram_T_207[287:0] : _GEN_7119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8170 = 10'h124 == _T_21 ? _ram_T_207[287:0] : _GEN_7120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8171 = 10'h125 == _T_21 ? _ram_T_207[287:0] : _GEN_7121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8172 = 10'h126 == _T_21 ? _ram_T_207[287:0] : _GEN_7122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8173 = 10'h127 == _T_21 ? _ram_T_207[287:0] : _GEN_7123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8174 = 10'h128 == _T_21 ? _ram_T_207[287:0] : _GEN_7124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8175 = 10'h129 == _T_21 ? _ram_T_207[287:0] : _GEN_7125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8176 = 10'h12a == _T_21 ? _ram_T_207[287:0] : _GEN_7126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8177 = 10'h12b == _T_21 ? _ram_T_207[287:0] : _GEN_7127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8178 = 10'h12c == _T_21 ? _ram_T_207[287:0] : _GEN_7128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8179 = 10'h12d == _T_21 ? _ram_T_207[287:0] : _GEN_7129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8180 = 10'h12e == _T_21 ? _ram_T_207[287:0] : _GEN_7130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8181 = 10'h12f == _T_21 ? _ram_T_207[287:0] : _GEN_7131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8182 = 10'h130 == _T_21 ? _ram_T_207[287:0] : _GEN_7132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8183 = 10'h131 == _T_21 ? _ram_T_207[287:0] : _GEN_7133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8184 = 10'h132 == _T_21 ? _ram_T_207[287:0] : _GEN_7134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8185 = 10'h133 == _T_21 ? _ram_T_207[287:0] : _GEN_7135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8186 = 10'h134 == _T_21 ? _ram_T_207[287:0] : _GEN_7136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8187 = 10'h135 == _T_21 ? _ram_T_207[287:0] : _GEN_7137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8188 = 10'h136 == _T_21 ? _ram_T_207[287:0] : _GEN_7138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8189 = 10'h137 == _T_21 ? _ram_T_207[287:0] : _GEN_7139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8190 = 10'h138 == _T_21 ? _ram_T_207[287:0] : _GEN_7140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8191 = 10'h139 == _T_21 ? _ram_T_207[287:0] : _GEN_7141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8192 = 10'h13a == _T_21 ? _ram_T_207[287:0] : _GEN_7142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8193 = 10'h13b == _T_21 ? _ram_T_207[287:0] : _GEN_7143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8194 = 10'h13c == _T_21 ? _ram_T_207[287:0] : _GEN_7144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8195 = 10'h13d == _T_21 ? _ram_T_207[287:0] : _GEN_7145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8196 = 10'h13e == _T_21 ? _ram_T_207[287:0] : _GEN_7146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8197 = 10'h13f == _T_21 ? _ram_T_207[287:0] : _GEN_7147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8198 = 10'h140 == _T_21 ? _ram_T_207[287:0] : _GEN_7148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8199 = 10'h141 == _T_21 ? _ram_T_207[287:0] : _GEN_7149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8200 = 10'h142 == _T_21 ? _ram_T_207[287:0] : _GEN_7150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8201 = 10'h143 == _T_21 ? _ram_T_207[287:0] : _GEN_7151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8202 = 10'h144 == _T_21 ? _ram_T_207[287:0] : _GEN_7152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8203 = 10'h145 == _T_21 ? _ram_T_207[287:0] : _GEN_7153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8204 = 10'h146 == _T_21 ? _ram_T_207[287:0] : _GEN_7154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8205 = 10'h147 == _T_21 ? _ram_T_207[287:0] : _GEN_7155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8206 = 10'h148 == _T_21 ? _ram_T_207[287:0] : _GEN_7156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8207 = 10'h149 == _T_21 ? _ram_T_207[287:0] : _GEN_7157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8208 = 10'h14a == _T_21 ? _ram_T_207[287:0] : _GEN_7158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8209 = 10'h14b == _T_21 ? _ram_T_207[287:0] : _GEN_7159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8210 = 10'h14c == _T_21 ? _ram_T_207[287:0] : _GEN_7160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8211 = 10'h14d == _T_21 ? _ram_T_207[287:0] : _GEN_7161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8212 = 10'h14e == _T_21 ? _ram_T_207[287:0] : _GEN_7162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8213 = 10'h14f == _T_21 ? _ram_T_207[287:0] : _GEN_7163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8214 = 10'h150 == _T_21 ? _ram_T_207[287:0] : _GEN_7164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8215 = 10'h151 == _T_21 ? _ram_T_207[287:0] : _GEN_7165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8216 = 10'h152 == _T_21 ? _ram_T_207[287:0] : _GEN_7166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8217 = 10'h153 == _T_21 ? _ram_T_207[287:0] : _GEN_7167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8218 = 10'h154 == _T_21 ? _ram_T_207[287:0] : _GEN_7168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8219 = 10'h155 == _T_21 ? _ram_T_207[287:0] : _GEN_7169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8220 = 10'h156 == _T_21 ? _ram_T_207[287:0] : _GEN_7170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8221 = 10'h157 == _T_21 ? _ram_T_207[287:0] : _GEN_7171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8222 = 10'h158 == _T_21 ? _ram_T_207[287:0] : _GEN_7172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8223 = 10'h159 == _T_21 ? _ram_T_207[287:0] : _GEN_7173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8224 = 10'h15a == _T_21 ? _ram_T_207[287:0] : _GEN_7174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8225 = 10'h15b == _T_21 ? _ram_T_207[287:0] : _GEN_7175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8226 = 10'h15c == _T_21 ? _ram_T_207[287:0] : _GEN_7176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8227 = 10'h15d == _T_21 ? _ram_T_207[287:0] : _GEN_7177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8228 = 10'h15e == _T_21 ? _ram_T_207[287:0] : _GEN_7178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8229 = 10'h15f == _T_21 ? _ram_T_207[287:0] : _GEN_7179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8230 = 10'h160 == _T_21 ? _ram_T_207[287:0] : _GEN_7180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8231 = 10'h161 == _T_21 ? _ram_T_207[287:0] : _GEN_7181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8232 = 10'h162 == _T_21 ? _ram_T_207[287:0] : _GEN_7182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8233 = 10'h163 == _T_21 ? _ram_T_207[287:0] : _GEN_7183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8234 = 10'h164 == _T_21 ? _ram_T_207[287:0] : _GEN_7184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8235 = 10'h165 == _T_21 ? _ram_T_207[287:0] : _GEN_7185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8236 = 10'h166 == _T_21 ? _ram_T_207[287:0] : _GEN_7186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8237 = 10'h167 == _T_21 ? _ram_T_207[287:0] : _GEN_7187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8238 = 10'h168 == _T_21 ? _ram_T_207[287:0] : _GEN_7188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8239 = 10'h169 == _T_21 ? _ram_T_207[287:0] : _GEN_7189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8240 = 10'h16a == _T_21 ? _ram_T_207[287:0] : _GEN_7190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8241 = 10'h16b == _T_21 ? _ram_T_207[287:0] : _GEN_7191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8242 = 10'h16c == _T_21 ? _ram_T_207[287:0] : _GEN_7192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8243 = 10'h16d == _T_21 ? _ram_T_207[287:0] : _GEN_7193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8244 = 10'h16e == _T_21 ? _ram_T_207[287:0] : _GEN_7194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8245 = 10'h16f == _T_21 ? _ram_T_207[287:0] : _GEN_7195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8246 = 10'h170 == _T_21 ? _ram_T_207[287:0] : _GEN_7196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8247 = 10'h171 == _T_21 ? _ram_T_207[287:0] : _GEN_7197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8248 = 10'h172 == _T_21 ? _ram_T_207[287:0] : _GEN_7198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8249 = 10'h173 == _T_21 ? _ram_T_207[287:0] : _GEN_7199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8250 = 10'h174 == _T_21 ? _ram_T_207[287:0] : _GEN_7200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8251 = 10'h175 == _T_21 ? _ram_T_207[287:0] : _GEN_7201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8252 = 10'h176 == _T_21 ? _ram_T_207[287:0] : _GEN_7202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8253 = 10'h177 == _T_21 ? _ram_T_207[287:0] : _GEN_7203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8254 = 10'h178 == _T_21 ? _ram_T_207[287:0] : _GEN_7204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8255 = 10'h179 == _T_21 ? _ram_T_207[287:0] : _GEN_7205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8256 = 10'h17a == _T_21 ? _ram_T_207[287:0] : _GEN_7206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8257 = 10'h17b == _T_21 ? _ram_T_207[287:0] : _GEN_7207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8258 = 10'h17c == _T_21 ? _ram_T_207[287:0] : _GEN_7208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8259 = 10'h17d == _T_21 ? _ram_T_207[287:0] : _GEN_7209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8260 = 10'h17e == _T_21 ? _ram_T_207[287:0] : _GEN_7210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8261 = 10'h17f == _T_21 ? _ram_T_207[287:0] : _GEN_7211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8262 = 10'h180 == _T_21 ? _ram_T_207[287:0] : _GEN_7212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8263 = 10'h181 == _T_21 ? _ram_T_207[287:0] : _GEN_7213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8264 = 10'h182 == _T_21 ? _ram_T_207[287:0] : _GEN_7214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8265 = 10'h183 == _T_21 ? _ram_T_207[287:0] : _GEN_7215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8266 = 10'h184 == _T_21 ? _ram_T_207[287:0] : _GEN_7216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8267 = 10'h185 == _T_21 ? _ram_T_207[287:0] : _GEN_7217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8268 = 10'h186 == _T_21 ? _ram_T_207[287:0] : _GEN_7218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8269 = 10'h187 == _T_21 ? _ram_T_207[287:0] : _GEN_7219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8270 = 10'h188 == _T_21 ? _ram_T_207[287:0] : _GEN_7220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8271 = 10'h189 == _T_21 ? _ram_T_207[287:0] : _GEN_7221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8272 = 10'h18a == _T_21 ? _ram_T_207[287:0] : _GEN_7222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8273 = 10'h18b == _T_21 ? _ram_T_207[287:0] : _GEN_7223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8274 = 10'h18c == _T_21 ? _ram_T_207[287:0] : _GEN_7224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8275 = 10'h18d == _T_21 ? _ram_T_207[287:0] : _GEN_7225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8276 = 10'h18e == _T_21 ? _ram_T_207[287:0] : _GEN_7226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8277 = 10'h18f == _T_21 ? _ram_T_207[287:0] : _GEN_7227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8278 = 10'h190 == _T_21 ? _ram_T_207[287:0] : _GEN_7228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8279 = 10'h191 == _T_21 ? _ram_T_207[287:0] : _GEN_7229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8280 = 10'h192 == _T_21 ? _ram_T_207[287:0] : _GEN_7230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8281 = 10'h193 == _T_21 ? _ram_T_207[287:0] : _GEN_7231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8282 = 10'h194 == _T_21 ? _ram_T_207[287:0] : _GEN_7232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8283 = 10'h195 == _T_21 ? _ram_T_207[287:0] : _GEN_7233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8284 = 10'h196 == _T_21 ? _ram_T_207[287:0] : _GEN_7234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8285 = 10'h197 == _T_21 ? _ram_T_207[287:0] : _GEN_7235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8286 = 10'h198 == _T_21 ? _ram_T_207[287:0] : _GEN_7236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8287 = 10'h199 == _T_21 ? _ram_T_207[287:0] : _GEN_7237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8288 = 10'h19a == _T_21 ? _ram_T_207[287:0] : _GEN_7238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8289 = 10'h19b == _T_21 ? _ram_T_207[287:0] : _GEN_7239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8290 = 10'h19c == _T_21 ? _ram_T_207[287:0] : _GEN_7240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8291 = 10'h19d == _T_21 ? _ram_T_207[287:0] : _GEN_7241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8292 = 10'h19e == _T_21 ? _ram_T_207[287:0] : _GEN_7242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8293 = 10'h19f == _T_21 ? _ram_T_207[287:0] : _GEN_7243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8294 = 10'h1a0 == _T_21 ? _ram_T_207[287:0] : _GEN_7244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8295 = 10'h1a1 == _T_21 ? _ram_T_207[287:0] : _GEN_7245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8296 = 10'h1a2 == _T_21 ? _ram_T_207[287:0] : _GEN_7246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8297 = 10'h1a3 == _T_21 ? _ram_T_207[287:0] : _GEN_7247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8298 = 10'h1a4 == _T_21 ? _ram_T_207[287:0] : _GEN_7248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8299 = 10'h1a5 == _T_21 ? _ram_T_207[287:0] : _GEN_7249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8300 = 10'h1a6 == _T_21 ? _ram_T_207[287:0] : _GEN_7250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8301 = 10'h1a7 == _T_21 ? _ram_T_207[287:0] : _GEN_7251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8302 = 10'h1a8 == _T_21 ? _ram_T_207[287:0] : _GEN_7252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8303 = 10'h1a9 == _T_21 ? _ram_T_207[287:0] : _GEN_7253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8304 = 10'h1aa == _T_21 ? _ram_T_207[287:0] : _GEN_7254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8305 = 10'h1ab == _T_21 ? _ram_T_207[287:0] : _GEN_7255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8306 = 10'h1ac == _T_21 ? _ram_T_207[287:0] : _GEN_7256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8307 = 10'h1ad == _T_21 ? _ram_T_207[287:0] : _GEN_7257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8308 = 10'h1ae == _T_21 ? _ram_T_207[287:0] : _GEN_7258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8309 = 10'h1af == _T_21 ? _ram_T_207[287:0] : _GEN_7259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8310 = 10'h1b0 == _T_21 ? _ram_T_207[287:0] : _GEN_7260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8311 = 10'h1b1 == _T_21 ? _ram_T_207[287:0] : _GEN_7261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8312 = 10'h1b2 == _T_21 ? _ram_T_207[287:0] : _GEN_7262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8313 = 10'h1b3 == _T_21 ? _ram_T_207[287:0] : _GEN_7263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8314 = 10'h1b4 == _T_21 ? _ram_T_207[287:0] : _GEN_7264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8315 = 10'h1b5 == _T_21 ? _ram_T_207[287:0] : _GEN_7265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8316 = 10'h1b6 == _T_21 ? _ram_T_207[287:0] : _GEN_7266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8317 = 10'h1b7 == _T_21 ? _ram_T_207[287:0] : _GEN_7267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8318 = 10'h1b8 == _T_21 ? _ram_T_207[287:0] : _GEN_7268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8319 = 10'h1b9 == _T_21 ? _ram_T_207[287:0] : _GEN_7269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8320 = 10'h1ba == _T_21 ? _ram_T_207[287:0] : _GEN_7270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8321 = 10'h1bb == _T_21 ? _ram_T_207[287:0] : _GEN_7271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8322 = 10'h1bc == _T_21 ? _ram_T_207[287:0] : _GEN_7272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8323 = 10'h1bd == _T_21 ? _ram_T_207[287:0] : _GEN_7273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8324 = 10'h1be == _T_21 ? _ram_T_207[287:0] : _GEN_7274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8325 = 10'h1bf == _T_21 ? _ram_T_207[287:0] : _GEN_7275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8326 = 10'h1c0 == _T_21 ? _ram_T_207[287:0] : _GEN_7276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8327 = 10'h1c1 == _T_21 ? _ram_T_207[287:0] : _GEN_7277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8328 = 10'h1c2 == _T_21 ? _ram_T_207[287:0] : _GEN_7278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8329 = 10'h1c3 == _T_21 ? _ram_T_207[287:0] : _GEN_7279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8330 = 10'h1c4 == _T_21 ? _ram_T_207[287:0] : _GEN_7280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8331 = 10'h1c5 == _T_21 ? _ram_T_207[287:0] : _GEN_7281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8332 = 10'h1c6 == _T_21 ? _ram_T_207[287:0] : _GEN_7282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8333 = 10'h1c7 == _T_21 ? _ram_T_207[287:0] : _GEN_7283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8334 = 10'h1c8 == _T_21 ? _ram_T_207[287:0] : _GEN_7284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8335 = 10'h1c9 == _T_21 ? _ram_T_207[287:0] : _GEN_7285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8336 = 10'h1ca == _T_21 ? _ram_T_207[287:0] : _GEN_7286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8337 = 10'h1cb == _T_21 ? _ram_T_207[287:0] : _GEN_7287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8338 = 10'h1cc == _T_21 ? _ram_T_207[287:0] : _GEN_7288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8339 = 10'h1cd == _T_21 ? _ram_T_207[287:0] : _GEN_7289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8340 = 10'h1ce == _T_21 ? _ram_T_207[287:0] : _GEN_7290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8341 = 10'h1cf == _T_21 ? _ram_T_207[287:0] : _GEN_7291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8342 = 10'h1d0 == _T_21 ? _ram_T_207[287:0] : _GEN_7292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8343 = 10'h1d1 == _T_21 ? _ram_T_207[287:0] : _GEN_7293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8344 = 10'h1d2 == _T_21 ? _ram_T_207[287:0] : _GEN_7294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8345 = 10'h1d3 == _T_21 ? _ram_T_207[287:0] : _GEN_7295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8346 = 10'h1d4 == _T_21 ? _ram_T_207[287:0] : _GEN_7296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8347 = 10'h1d5 == _T_21 ? _ram_T_207[287:0] : _GEN_7297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8348 = 10'h1d6 == _T_21 ? _ram_T_207[287:0] : _GEN_7298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8349 = 10'h1d7 == _T_21 ? _ram_T_207[287:0] : _GEN_7299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8350 = 10'h1d8 == _T_21 ? _ram_T_207[287:0] : _GEN_7300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8351 = 10'h1d9 == _T_21 ? _ram_T_207[287:0] : _GEN_7301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8352 = 10'h1da == _T_21 ? _ram_T_207[287:0] : _GEN_7302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8353 = 10'h1db == _T_21 ? _ram_T_207[287:0] : _GEN_7303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8354 = 10'h1dc == _T_21 ? _ram_T_207[287:0] : _GEN_7304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8355 = 10'h1dd == _T_21 ? _ram_T_207[287:0] : _GEN_7305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8356 = 10'h1de == _T_21 ? _ram_T_207[287:0] : _GEN_7306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8357 = 10'h1df == _T_21 ? _ram_T_207[287:0] : _GEN_7307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8358 = 10'h1e0 == _T_21 ? _ram_T_207[287:0] : _GEN_7308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8359 = 10'h1e1 == _T_21 ? _ram_T_207[287:0] : _GEN_7309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8360 = 10'h1e2 == _T_21 ? _ram_T_207[287:0] : _GEN_7310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8361 = 10'h1e3 == _T_21 ? _ram_T_207[287:0] : _GEN_7311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8362 = 10'h1e4 == _T_21 ? _ram_T_207[287:0] : _GEN_7312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8363 = 10'h1e5 == _T_21 ? _ram_T_207[287:0] : _GEN_7313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8364 = 10'h1e6 == _T_21 ? _ram_T_207[287:0] : _GEN_7314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8365 = 10'h1e7 == _T_21 ? _ram_T_207[287:0] : _GEN_7315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8366 = 10'h1e8 == _T_21 ? _ram_T_207[287:0] : _GEN_7316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8367 = 10'h1e9 == _T_21 ? _ram_T_207[287:0] : _GEN_7317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8368 = 10'h1ea == _T_21 ? _ram_T_207[287:0] : _GEN_7318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8369 = 10'h1eb == _T_21 ? _ram_T_207[287:0] : _GEN_7319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8370 = 10'h1ec == _T_21 ? _ram_T_207[287:0] : _GEN_7320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8371 = 10'h1ed == _T_21 ? _ram_T_207[287:0] : _GEN_7321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8372 = 10'h1ee == _T_21 ? _ram_T_207[287:0] : _GEN_7322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8373 = 10'h1ef == _T_21 ? _ram_T_207[287:0] : _GEN_7323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8374 = 10'h1f0 == _T_21 ? _ram_T_207[287:0] : _GEN_7324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8375 = 10'h1f1 == _T_21 ? _ram_T_207[287:0] : _GEN_7325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8376 = 10'h1f2 == _T_21 ? _ram_T_207[287:0] : _GEN_7326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8377 = 10'h1f3 == _T_21 ? _ram_T_207[287:0] : _GEN_7327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8378 = 10'h1f4 == _T_21 ? _ram_T_207[287:0] : _GEN_7328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8379 = 10'h1f5 == _T_21 ? _ram_T_207[287:0] : _GEN_7329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8380 = 10'h1f6 == _T_21 ? _ram_T_207[287:0] : _GEN_7330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8381 = 10'h1f7 == _T_21 ? _ram_T_207[287:0] : _GEN_7331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8382 = 10'h1f8 == _T_21 ? _ram_T_207[287:0] : _GEN_7332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8383 = 10'h1f9 == _T_21 ? _ram_T_207[287:0] : _GEN_7333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8384 = 10'h1fa == _T_21 ? _ram_T_207[287:0] : _GEN_7334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8385 = 10'h1fb == _T_21 ? _ram_T_207[287:0] : _GEN_7335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8386 = 10'h1fc == _T_21 ? _ram_T_207[287:0] : _GEN_7336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8387 = 10'h1fd == _T_21 ? _ram_T_207[287:0] : _GEN_7337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8388 = 10'h1fe == _T_21 ? _ram_T_207[287:0] : _GEN_7338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8389 = 10'h1ff == _T_21 ? _ram_T_207[287:0] : _GEN_7339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8390 = 10'h200 == _T_21 ? _ram_T_207[287:0] : _GEN_7340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8391 = 10'h201 == _T_21 ? _ram_T_207[287:0] : _GEN_7341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8392 = 10'h202 == _T_21 ? _ram_T_207[287:0] : _GEN_7342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8393 = 10'h203 == _T_21 ? _ram_T_207[287:0] : _GEN_7343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8394 = 10'h204 == _T_21 ? _ram_T_207[287:0] : _GEN_7344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8395 = 10'h205 == _T_21 ? _ram_T_207[287:0] : _GEN_7345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8396 = 10'h206 == _T_21 ? _ram_T_207[287:0] : _GEN_7346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8397 = 10'h207 == _T_21 ? _ram_T_207[287:0] : _GEN_7347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8398 = 10'h208 == _T_21 ? _ram_T_207[287:0] : _GEN_7348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8399 = 10'h209 == _T_21 ? _ram_T_207[287:0] : _GEN_7349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8400 = 10'h20a == _T_21 ? _ram_T_207[287:0] : _GEN_7350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8401 = 10'h20b == _T_21 ? _ram_T_207[287:0] : _GEN_7351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8402 = 10'h20c == _T_21 ? _ram_T_207[287:0] : _GEN_7352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_23 = h + 10'h8; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_8 = vga_mem_ram_MPORT_72_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_8 = vga_mem_ram_MPORT_73_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_8 = vga_mem_ram_MPORT_74_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_8 = vga_mem_ram_MPORT_75_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_8 = vga_mem_ram_MPORT_76_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_8 = vga_mem_ram_MPORT_77_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_8 = vga_mem_ram_MPORT_78_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_8 = vga_mem_ram_MPORT_79_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_8 = vga_mem_ram_MPORT_80_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_228 = {278'h0,ram_hi_hi_hi_lo_8,ram_hi_hi_lo_8,ram_hi_lo_hi_8,ram_hi_lo_lo_8,ram_lo_hi_hi_hi_8,
    ram_lo_hi_hi_lo_8,ram_lo_hi_lo_8,ram_lo_lo_hi_8,ram_lo_lo_lo_8}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19076 = {{8191'd0}, _ram_T_228}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_232 = _GEN_19076 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_8404 = 10'h1 == _T_23 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8405 = 10'h2 == _T_23 ? ram_2 : _GEN_8404; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8406 = 10'h3 == _T_23 ? ram_3 : _GEN_8405; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8407 = 10'h4 == _T_23 ? ram_4 : _GEN_8406; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8408 = 10'h5 == _T_23 ? ram_5 : _GEN_8407; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8409 = 10'h6 == _T_23 ? ram_6 : _GEN_8408; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8410 = 10'h7 == _T_23 ? ram_7 : _GEN_8409; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8411 = 10'h8 == _T_23 ? ram_8 : _GEN_8410; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8412 = 10'h9 == _T_23 ? ram_9 : _GEN_8411; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8413 = 10'ha == _T_23 ? ram_10 : _GEN_8412; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8414 = 10'hb == _T_23 ? ram_11 : _GEN_8413; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8415 = 10'hc == _T_23 ? ram_12 : _GEN_8414; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8416 = 10'hd == _T_23 ? ram_13 : _GEN_8415; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8417 = 10'he == _T_23 ? ram_14 : _GEN_8416; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8418 = 10'hf == _T_23 ? ram_15 : _GEN_8417; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8419 = 10'h10 == _T_23 ? ram_16 : _GEN_8418; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8420 = 10'h11 == _T_23 ? ram_17 : _GEN_8419; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8421 = 10'h12 == _T_23 ? ram_18 : _GEN_8420; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8422 = 10'h13 == _T_23 ? ram_19 : _GEN_8421; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8423 = 10'h14 == _T_23 ? ram_20 : _GEN_8422; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8424 = 10'h15 == _T_23 ? ram_21 : _GEN_8423; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8425 = 10'h16 == _T_23 ? ram_22 : _GEN_8424; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8426 = 10'h17 == _T_23 ? ram_23 : _GEN_8425; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8427 = 10'h18 == _T_23 ? ram_24 : _GEN_8426; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8428 = 10'h19 == _T_23 ? ram_25 : _GEN_8427; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8429 = 10'h1a == _T_23 ? ram_26 : _GEN_8428; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8430 = 10'h1b == _T_23 ? ram_27 : _GEN_8429; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8431 = 10'h1c == _T_23 ? ram_28 : _GEN_8430; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8432 = 10'h1d == _T_23 ? ram_29 : _GEN_8431; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8433 = 10'h1e == _T_23 ? ram_30 : _GEN_8432; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8434 = 10'h1f == _T_23 ? ram_31 : _GEN_8433; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8435 = 10'h20 == _T_23 ? ram_32 : _GEN_8434; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8436 = 10'h21 == _T_23 ? ram_33 : _GEN_8435; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8437 = 10'h22 == _T_23 ? ram_34 : _GEN_8436; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8438 = 10'h23 == _T_23 ? ram_35 : _GEN_8437; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8439 = 10'h24 == _T_23 ? ram_36 : _GEN_8438; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8440 = 10'h25 == _T_23 ? ram_37 : _GEN_8439; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8441 = 10'h26 == _T_23 ? ram_38 : _GEN_8440; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8442 = 10'h27 == _T_23 ? ram_39 : _GEN_8441; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8443 = 10'h28 == _T_23 ? ram_40 : _GEN_8442; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8444 = 10'h29 == _T_23 ? ram_41 : _GEN_8443; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8445 = 10'h2a == _T_23 ? ram_42 : _GEN_8444; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8446 = 10'h2b == _T_23 ? ram_43 : _GEN_8445; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8447 = 10'h2c == _T_23 ? ram_44 : _GEN_8446; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8448 = 10'h2d == _T_23 ? ram_45 : _GEN_8447; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8449 = 10'h2e == _T_23 ? ram_46 : _GEN_8448; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8450 = 10'h2f == _T_23 ? ram_47 : _GEN_8449; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8451 = 10'h30 == _T_23 ? ram_48 : _GEN_8450; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8452 = 10'h31 == _T_23 ? ram_49 : _GEN_8451; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8453 = 10'h32 == _T_23 ? ram_50 : _GEN_8452; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8454 = 10'h33 == _T_23 ? ram_51 : _GEN_8453; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8455 = 10'h34 == _T_23 ? ram_52 : _GEN_8454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8456 = 10'h35 == _T_23 ? ram_53 : _GEN_8455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8457 = 10'h36 == _T_23 ? ram_54 : _GEN_8456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8458 = 10'h37 == _T_23 ? ram_55 : _GEN_8457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8459 = 10'h38 == _T_23 ? ram_56 : _GEN_8458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8460 = 10'h39 == _T_23 ? ram_57 : _GEN_8459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8461 = 10'h3a == _T_23 ? ram_58 : _GEN_8460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8462 = 10'h3b == _T_23 ? ram_59 : _GEN_8461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8463 = 10'h3c == _T_23 ? ram_60 : _GEN_8462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8464 = 10'h3d == _T_23 ? ram_61 : _GEN_8463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8465 = 10'h3e == _T_23 ? ram_62 : _GEN_8464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8466 = 10'h3f == _T_23 ? ram_63 : _GEN_8465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8467 = 10'h40 == _T_23 ? ram_64 : _GEN_8466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8468 = 10'h41 == _T_23 ? ram_65 : _GEN_8467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8469 = 10'h42 == _T_23 ? ram_66 : _GEN_8468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8470 = 10'h43 == _T_23 ? ram_67 : _GEN_8469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8471 = 10'h44 == _T_23 ? ram_68 : _GEN_8470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8472 = 10'h45 == _T_23 ? ram_69 : _GEN_8471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8473 = 10'h46 == _T_23 ? ram_70 : _GEN_8472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8474 = 10'h47 == _T_23 ? ram_71 : _GEN_8473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8475 = 10'h48 == _T_23 ? ram_72 : _GEN_8474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8476 = 10'h49 == _T_23 ? ram_73 : _GEN_8475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8477 = 10'h4a == _T_23 ? ram_74 : _GEN_8476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8478 = 10'h4b == _T_23 ? ram_75 : _GEN_8477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8479 = 10'h4c == _T_23 ? ram_76 : _GEN_8478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8480 = 10'h4d == _T_23 ? ram_77 : _GEN_8479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8481 = 10'h4e == _T_23 ? ram_78 : _GEN_8480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8482 = 10'h4f == _T_23 ? ram_79 : _GEN_8481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8483 = 10'h50 == _T_23 ? ram_80 : _GEN_8482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8484 = 10'h51 == _T_23 ? ram_81 : _GEN_8483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8485 = 10'h52 == _T_23 ? ram_82 : _GEN_8484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8486 = 10'h53 == _T_23 ? ram_83 : _GEN_8485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8487 = 10'h54 == _T_23 ? ram_84 : _GEN_8486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8488 = 10'h55 == _T_23 ? ram_85 : _GEN_8487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8489 = 10'h56 == _T_23 ? ram_86 : _GEN_8488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8490 = 10'h57 == _T_23 ? ram_87 : _GEN_8489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8491 = 10'h58 == _T_23 ? ram_88 : _GEN_8490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8492 = 10'h59 == _T_23 ? ram_89 : _GEN_8491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8493 = 10'h5a == _T_23 ? ram_90 : _GEN_8492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8494 = 10'h5b == _T_23 ? ram_91 : _GEN_8493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8495 = 10'h5c == _T_23 ? ram_92 : _GEN_8494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8496 = 10'h5d == _T_23 ? ram_93 : _GEN_8495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8497 = 10'h5e == _T_23 ? ram_94 : _GEN_8496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8498 = 10'h5f == _T_23 ? ram_95 : _GEN_8497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8499 = 10'h60 == _T_23 ? ram_96 : _GEN_8498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8500 = 10'h61 == _T_23 ? ram_97 : _GEN_8499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8501 = 10'h62 == _T_23 ? ram_98 : _GEN_8500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8502 = 10'h63 == _T_23 ? ram_99 : _GEN_8501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8503 = 10'h64 == _T_23 ? ram_100 : _GEN_8502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8504 = 10'h65 == _T_23 ? ram_101 : _GEN_8503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8505 = 10'h66 == _T_23 ? ram_102 : _GEN_8504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8506 = 10'h67 == _T_23 ? ram_103 : _GEN_8505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8507 = 10'h68 == _T_23 ? ram_104 : _GEN_8506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8508 = 10'h69 == _T_23 ? ram_105 : _GEN_8507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8509 = 10'h6a == _T_23 ? ram_106 : _GEN_8508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8510 = 10'h6b == _T_23 ? ram_107 : _GEN_8509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8511 = 10'h6c == _T_23 ? ram_108 : _GEN_8510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8512 = 10'h6d == _T_23 ? ram_109 : _GEN_8511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8513 = 10'h6e == _T_23 ? ram_110 : _GEN_8512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8514 = 10'h6f == _T_23 ? ram_111 : _GEN_8513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8515 = 10'h70 == _T_23 ? ram_112 : _GEN_8514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8516 = 10'h71 == _T_23 ? ram_113 : _GEN_8515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8517 = 10'h72 == _T_23 ? ram_114 : _GEN_8516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8518 = 10'h73 == _T_23 ? ram_115 : _GEN_8517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8519 = 10'h74 == _T_23 ? ram_116 : _GEN_8518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8520 = 10'h75 == _T_23 ? ram_117 : _GEN_8519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8521 = 10'h76 == _T_23 ? ram_118 : _GEN_8520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8522 = 10'h77 == _T_23 ? ram_119 : _GEN_8521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8523 = 10'h78 == _T_23 ? ram_120 : _GEN_8522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8524 = 10'h79 == _T_23 ? ram_121 : _GEN_8523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8525 = 10'h7a == _T_23 ? ram_122 : _GEN_8524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8526 = 10'h7b == _T_23 ? ram_123 : _GEN_8525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8527 = 10'h7c == _T_23 ? ram_124 : _GEN_8526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8528 = 10'h7d == _T_23 ? ram_125 : _GEN_8527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8529 = 10'h7e == _T_23 ? ram_126 : _GEN_8528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8530 = 10'h7f == _T_23 ? ram_127 : _GEN_8529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8531 = 10'h80 == _T_23 ? ram_128 : _GEN_8530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8532 = 10'h81 == _T_23 ? ram_129 : _GEN_8531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8533 = 10'h82 == _T_23 ? ram_130 : _GEN_8532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8534 = 10'h83 == _T_23 ? ram_131 : _GEN_8533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8535 = 10'h84 == _T_23 ? ram_132 : _GEN_8534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8536 = 10'h85 == _T_23 ? ram_133 : _GEN_8535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8537 = 10'h86 == _T_23 ? ram_134 : _GEN_8536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8538 = 10'h87 == _T_23 ? ram_135 : _GEN_8537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8539 = 10'h88 == _T_23 ? ram_136 : _GEN_8538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8540 = 10'h89 == _T_23 ? ram_137 : _GEN_8539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8541 = 10'h8a == _T_23 ? ram_138 : _GEN_8540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8542 = 10'h8b == _T_23 ? ram_139 : _GEN_8541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8543 = 10'h8c == _T_23 ? ram_140 : _GEN_8542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8544 = 10'h8d == _T_23 ? ram_141 : _GEN_8543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8545 = 10'h8e == _T_23 ? ram_142 : _GEN_8544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8546 = 10'h8f == _T_23 ? ram_143 : _GEN_8545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8547 = 10'h90 == _T_23 ? ram_144 : _GEN_8546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8548 = 10'h91 == _T_23 ? ram_145 : _GEN_8547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8549 = 10'h92 == _T_23 ? ram_146 : _GEN_8548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8550 = 10'h93 == _T_23 ? ram_147 : _GEN_8549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8551 = 10'h94 == _T_23 ? ram_148 : _GEN_8550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8552 = 10'h95 == _T_23 ? ram_149 : _GEN_8551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8553 = 10'h96 == _T_23 ? ram_150 : _GEN_8552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8554 = 10'h97 == _T_23 ? ram_151 : _GEN_8553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8555 = 10'h98 == _T_23 ? ram_152 : _GEN_8554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8556 = 10'h99 == _T_23 ? ram_153 : _GEN_8555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8557 = 10'h9a == _T_23 ? ram_154 : _GEN_8556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8558 = 10'h9b == _T_23 ? ram_155 : _GEN_8557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8559 = 10'h9c == _T_23 ? ram_156 : _GEN_8558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8560 = 10'h9d == _T_23 ? ram_157 : _GEN_8559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8561 = 10'h9e == _T_23 ? ram_158 : _GEN_8560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8562 = 10'h9f == _T_23 ? ram_159 : _GEN_8561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8563 = 10'ha0 == _T_23 ? ram_160 : _GEN_8562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8564 = 10'ha1 == _T_23 ? ram_161 : _GEN_8563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8565 = 10'ha2 == _T_23 ? ram_162 : _GEN_8564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8566 = 10'ha3 == _T_23 ? ram_163 : _GEN_8565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8567 = 10'ha4 == _T_23 ? ram_164 : _GEN_8566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8568 = 10'ha5 == _T_23 ? ram_165 : _GEN_8567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8569 = 10'ha6 == _T_23 ? ram_166 : _GEN_8568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8570 = 10'ha7 == _T_23 ? ram_167 : _GEN_8569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8571 = 10'ha8 == _T_23 ? ram_168 : _GEN_8570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8572 = 10'ha9 == _T_23 ? ram_169 : _GEN_8571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8573 = 10'haa == _T_23 ? ram_170 : _GEN_8572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8574 = 10'hab == _T_23 ? ram_171 : _GEN_8573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8575 = 10'hac == _T_23 ? ram_172 : _GEN_8574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8576 = 10'had == _T_23 ? ram_173 : _GEN_8575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8577 = 10'hae == _T_23 ? ram_174 : _GEN_8576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8578 = 10'haf == _T_23 ? ram_175 : _GEN_8577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8579 = 10'hb0 == _T_23 ? ram_176 : _GEN_8578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8580 = 10'hb1 == _T_23 ? ram_177 : _GEN_8579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8581 = 10'hb2 == _T_23 ? ram_178 : _GEN_8580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8582 = 10'hb3 == _T_23 ? ram_179 : _GEN_8581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8583 = 10'hb4 == _T_23 ? ram_180 : _GEN_8582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8584 = 10'hb5 == _T_23 ? ram_181 : _GEN_8583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8585 = 10'hb6 == _T_23 ? ram_182 : _GEN_8584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8586 = 10'hb7 == _T_23 ? ram_183 : _GEN_8585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8587 = 10'hb8 == _T_23 ? ram_184 : _GEN_8586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8588 = 10'hb9 == _T_23 ? ram_185 : _GEN_8587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8589 = 10'hba == _T_23 ? ram_186 : _GEN_8588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8590 = 10'hbb == _T_23 ? ram_187 : _GEN_8589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8591 = 10'hbc == _T_23 ? ram_188 : _GEN_8590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8592 = 10'hbd == _T_23 ? ram_189 : _GEN_8591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8593 = 10'hbe == _T_23 ? ram_190 : _GEN_8592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8594 = 10'hbf == _T_23 ? ram_191 : _GEN_8593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8595 = 10'hc0 == _T_23 ? ram_192 : _GEN_8594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8596 = 10'hc1 == _T_23 ? ram_193 : _GEN_8595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8597 = 10'hc2 == _T_23 ? ram_194 : _GEN_8596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8598 = 10'hc3 == _T_23 ? ram_195 : _GEN_8597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8599 = 10'hc4 == _T_23 ? ram_196 : _GEN_8598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8600 = 10'hc5 == _T_23 ? ram_197 : _GEN_8599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8601 = 10'hc6 == _T_23 ? ram_198 : _GEN_8600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8602 = 10'hc7 == _T_23 ? ram_199 : _GEN_8601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8603 = 10'hc8 == _T_23 ? ram_200 : _GEN_8602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8604 = 10'hc9 == _T_23 ? ram_201 : _GEN_8603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8605 = 10'hca == _T_23 ? ram_202 : _GEN_8604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8606 = 10'hcb == _T_23 ? ram_203 : _GEN_8605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8607 = 10'hcc == _T_23 ? ram_204 : _GEN_8606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8608 = 10'hcd == _T_23 ? ram_205 : _GEN_8607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8609 = 10'hce == _T_23 ? ram_206 : _GEN_8608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8610 = 10'hcf == _T_23 ? ram_207 : _GEN_8609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8611 = 10'hd0 == _T_23 ? ram_208 : _GEN_8610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8612 = 10'hd1 == _T_23 ? ram_209 : _GEN_8611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8613 = 10'hd2 == _T_23 ? ram_210 : _GEN_8612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8614 = 10'hd3 == _T_23 ? ram_211 : _GEN_8613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8615 = 10'hd4 == _T_23 ? ram_212 : _GEN_8614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8616 = 10'hd5 == _T_23 ? ram_213 : _GEN_8615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8617 = 10'hd6 == _T_23 ? ram_214 : _GEN_8616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8618 = 10'hd7 == _T_23 ? ram_215 : _GEN_8617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8619 = 10'hd8 == _T_23 ? ram_216 : _GEN_8618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8620 = 10'hd9 == _T_23 ? ram_217 : _GEN_8619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8621 = 10'hda == _T_23 ? ram_218 : _GEN_8620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8622 = 10'hdb == _T_23 ? ram_219 : _GEN_8621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8623 = 10'hdc == _T_23 ? ram_220 : _GEN_8622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8624 = 10'hdd == _T_23 ? ram_221 : _GEN_8623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8625 = 10'hde == _T_23 ? ram_222 : _GEN_8624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8626 = 10'hdf == _T_23 ? ram_223 : _GEN_8625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8627 = 10'he0 == _T_23 ? ram_224 : _GEN_8626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8628 = 10'he1 == _T_23 ? ram_225 : _GEN_8627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8629 = 10'he2 == _T_23 ? ram_226 : _GEN_8628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8630 = 10'he3 == _T_23 ? ram_227 : _GEN_8629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8631 = 10'he4 == _T_23 ? ram_228 : _GEN_8630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8632 = 10'he5 == _T_23 ? ram_229 : _GEN_8631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8633 = 10'he6 == _T_23 ? ram_230 : _GEN_8632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8634 = 10'he7 == _T_23 ? ram_231 : _GEN_8633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8635 = 10'he8 == _T_23 ? ram_232 : _GEN_8634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8636 = 10'he9 == _T_23 ? ram_233 : _GEN_8635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8637 = 10'hea == _T_23 ? ram_234 : _GEN_8636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8638 = 10'heb == _T_23 ? ram_235 : _GEN_8637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8639 = 10'hec == _T_23 ? ram_236 : _GEN_8638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8640 = 10'hed == _T_23 ? ram_237 : _GEN_8639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8641 = 10'hee == _T_23 ? ram_238 : _GEN_8640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8642 = 10'hef == _T_23 ? ram_239 : _GEN_8641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8643 = 10'hf0 == _T_23 ? ram_240 : _GEN_8642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8644 = 10'hf1 == _T_23 ? ram_241 : _GEN_8643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8645 = 10'hf2 == _T_23 ? ram_242 : _GEN_8644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8646 = 10'hf3 == _T_23 ? ram_243 : _GEN_8645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8647 = 10'hf4 == _T_23 ? ram_244 : _GEN_8646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8648 = 10'hf5 == _T_23 ? ram_245 : _GEN_8647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8649 = 10'hf6 == _T_23 ? ram_246 : _GEN_8648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8650 = 10'hf7 == _T_23 ? ram_247 : _GEN_8649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8651 = 10'hf8 == _T_23 ? ram_248 : _GEN_8650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8652 = 10'hf9 == _T_23 ? ram_249 : _GEN_8651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8653 = 10'hfa == _T_23 ? ram_250 : _GEN_8652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8654 = 10'hfb == _T_23 ? ram_251 : _GEN_8653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8655 = 10'hfc == _T_23 ? ram_252 : _GEN_8654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8656 = 10'hfd == _T_23 ? ram_253 : _GEN_8655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8657 = 10'hfe == _T_23 ? ram_254 : _GEN_8656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8658 = 10'hff == _T_23 ? ram_255 : _GEN_8657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8659 = 10'h100 == _T_23 ? ram_256 : _GEN_8658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8660 = 10'h101 == _T_23 ? ram_257 : _GEN_8659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8661 = 10'h102 == _T_23 ? ram_258 : _GEN_8660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8662 = 10'h103 == _T_23 ? ram_259 : _GEN_8661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8663 = 10'h104 == _T_23 ? ram_260 : _GEN_8662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8664 = 10'h105 == _T_23 ? ram_261 : _GEN_8663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8665 = 10'h106 == _T_23 ? ram_262 : _GEN_8664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8666 = 10'h107 == _T_23 ? ram_263 : _GEN_8665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8667 = 10'h108 == _T_23 ? ram_264 : _GEN_8666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8668 = 10'h109 == _T_23 ? ram_265 : _GEN_8667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8669 = 10'h10a == _T_23 ? ram_266 : _GEN_8668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8670 = 10'h10b == _T_23 ? ram_267 : _GEN_8669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8671 = 10'h10c == _T_23 ? ram_268 : _GEN_8670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8672 = 10'h10d == _T_23 ? ram_269 : _GEN_8671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8673 = 10'h10e == _T_23 ? ram_270 : _GEN_8672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8674 = 10'h10f == _T_23 ? ram_271 : _GEN_8673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8675 = 10'h110 == _T_23 ? ram_272 : _GEN_8674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8676 = 10'h111 == _T_23 ? ram_273 : _GEN_8675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8677 = 10'h112 == _T_23 ? ram_274 : _GEN_8676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8678 = 10'h113 == _T_23 ? ram_275 : _GEN_8677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8679 = 10'h114 == _T_23 ? ram_276 : _GEN_8678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8680 = 10'h115 == _T_23 ? ram_277 : _GEN_8679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8681 = 10'h116 == _T_23 ? ram_278 : _GEN_8680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8682 = 10'h117 == _T_23 ? ram_279 : _GEN_8681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8683 = 10'h118 == _T_23 ? ram_280 : _GEN_8682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8684 = 10'h119 == _T_23 ? ram_281 : _GEN_8683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8685 = 10'h11a == _T_23 ? ram_282 : _GEN_8684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8686 = 10'h11b == _T_23 ? ram_283 : _GEN_8685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8687 = 10'h11c == _T_23 ? ram_284 : _GEN_8686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8688 = 10'h11d == _T_23 ? ram_285 : _GEN_8687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8689 = 10'h11e == _T_23 ? ram_286 : _GEN_8688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8690 = 10'h11f == _T_23 ? ram_287 : _GEN_8689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8691 = 10'h120 == _T_23 ? ram_288 : _GEN_8690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8692 = 10'h121 == _T_23 ? ram_289 : _GEN_8691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8693 = 10'h122 == _T_23 ? ram_290 : _GEN_8692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8694 = 10'h123 == _T_23 ? ram_291 : _GEN_8693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8695 = 10'h124 == _T_23 ? ram_292 : _GEN_8694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8696 = 10'h125 == _T_23 ? ram_293 : _GEN_8695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8697 = 10'h126 == _T_23 ? ram_294 : _GEN_8696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8698 = 10'h127 == _T_23 ? ram_295 : _GEN_8697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8699 = 10'h128 == _T_23 ? ram_296 : _GEN_8698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8700 = 10'h129 == _T_23 ? ram_297 : _GEN_8699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8701 = 10'h12a == _T_23 ? ram_298 : _GEN_8700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8702 = 10'h12b == _T_23 ? ram_299 : _GEN_8701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8703 = 10'h12c == _T_23 ? ram_300 : _GEN_8702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8704 = 10'h12d == _T_23 ? ram_301 : _GEN_8703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8705 = 10'h12e == _T_23 ? ram_302 : _GEN_8704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8706 = 10'h12f == _T_23 ? ram_303 : _GEN_8705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8707 = 10'h130 == _T_23 ? ram_304 : _GEN_8706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8708 = 10'h131 == _T_23 ? ram_305 : _GEN_8707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8709 = 10'h132 == _T_23 ? ram_306 : _GEN_8708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8710 = 10'h133 == _T_23 ? ram_307 : _GEN_8709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8711 = 10'h134 == _T_23 ? ram_308 : _GEN_8710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8712 = 10'h135 == _T_23 ? ram_309 : _GEN_8711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8713 = 10'h136 == _T_23 ? ram_310 : _GEN_8712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8714 = 10'h137 == _T_23 ? ram_311 : _GEN_8713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8715 = 10'h138 == _T_23 ? ram_312 : _GEN_8714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8716 = 10'h139 == _T_23 ? ram_313 : _GEN_8715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8717 = 10'h13a == _T_23 ? ram_314 : _GEN_8716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8718 = 10'h13b == _T_23 ? ram_315 : _GEN_8717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8719 = 10'h13c == _T_23 ? ram_316 : _GEN_8718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8720 = 10'h13d == _T_23 ? ram_317 : _GEN_8719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8721 = 10'h13e == _T_23 ? ram_318 : _GEN_8720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8722 = 10'h13f == _T_23 ? ram_319 : _GEN_8721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8723 = 10'h140 == _T_23 ? ram_320 : _GEN_8722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8724 = 10'h141 == _T_23 ? ram_321 : _GEN_8723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8725 = 10'h142 == _T_23 ? ram_322 : _GEN_8724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8726 = 10'h143 == _T_23 ? ram_323 : _GEN_8725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8727 = 10'h144 == _T_23 ? ram_324 : _GEN_8726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8728 = 10'h145 == _T_23 ? ram_325 : _GEN_8727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8729 = 10'h146 == _T_23 ? ram_326 : _GEN_8728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8730 = 10'h147 == _T_23 ? ram_327 : _GEN_8729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8731 = 10'h148 == _T_23 ? ram_328 : _GEN_8730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8732 = 10'h149 == _T_23 ? ram_329 : _GEN_8731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8733 = 10'h14a == _T_23 ? ram_330 : _GEN_8732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8734 = 10'h14b == _T_23 ? ram_331 : _GEN_8733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8735 = 10'h14c == _T_23 ? ram_332 : _GEN_8734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8736 = 10'h14d == _T_23 ? ram_333 : _GEN_8735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8737 = 10'h14e == _T_23 ? ram_334 : _GEN_8736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8738 = 10'h14f == _T_23 ? ram_335 : _GEN_8737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8739 = 10'h150 == _T_23 ? ram_336 : _GEN_8738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8740 = 10'h151 == _T_23 ? ram_337 : _GEN_8739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8741 = 10'h152 == _T_23 ? ram_338 : _GEN_8740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8742 = 10'h153 == _T_23 ? ram_339 : _GEN_8741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8743 = 10'h154 == _T_23 ? ram_340 : _GEN_8742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8744 = 10'h155 == _T_23 ? ram_341 : _GEN_8743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8745 = 10'h156 == _T_23 ? ram_342 : _GEN_8744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8746 = 10'h157 == _T_23 ? ram_343 : _GEN_8745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8747 = 10'h158 == _T_23 ? ram_344 : _GEN_8746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8748 = 10'h159 == _T_23 ? ram_345 : _GEN_8747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8749 = 10'h15a == _T_23 ? ram_346 : _GEN_8748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8750 = 10'h15b == _T_23 ? ram_347 : _GEN_8749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8751 = 10'h15c == _T_23 ? ram_348 : _GEN_8750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8752 = 10'h15d == _T_23 ? ram_349 : _GEN_8751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8753 = 10'h15e == _T_23 ? ram_350 : _GEN_8752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8754 = 10'h15f == _T_23 ? ram_351 : _GEN_8753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8755 = 10'h160 == _T_23 ? ram_352 : _GEN_8754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8756 = 10'h161 == _T_23 ? ram_353 : _GEN_8755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8757 = 10'h162 == _T_23 ? ram_354 : _GEN_8756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8758 = 10'h163 == _T_23 ? ram_355 : _GEN_8757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8759 = 10'h164 == _T_23 ? ram_356 : _GEN_8758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8760 = 10'h165 == _T_23 ? ram_357 : _GEN_8759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8761 = 10'h166 == _T_23 ? ram_358 : _GEN_8760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8762 = 10'h167 == _T_23 ? ram_359 : _GEN_8761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8763 = 10'h168 == _T_23 ? ram_360 : _GEN_8762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8764 = 10'h169 == _T_23 ? ram_361 : _GEN_8763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8765 = 10'h16a == _T_23 ? ram_362 : _GEN_8764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8766 = 10'h16b == _T_23 ? ram_363 : _GEN_8765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8767 = 10'h16c == _T_23 ? ram_364 : _GEN_8766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8768 = 10'h16d == _T_23 ? ram_365 : _GEN_8767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8769 = 10'h16e == _T_23 ? ram_366 : _GEN_8768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8770 = 10'h16f == _T_23 ? ram_367 : _GEN_8769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8771 = 10'h170 == _T_23 ? ram_368 : _GEN_8770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8772 = 10'h171 == _T_23 ? ram_369 : _GEN_8771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8773 = 10'h172 == _T_23 ? ram_370 : _GEN_8772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8774 = 10'h173 == _T_23 ? ram_371 : _GEN_8773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8775 = 10'h174 == _T_23 ? ram_372 : _GEN_8774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8776 = 10'h175 == _T_23 ? ram_373 : _GEN_8775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8777 = 10'h176 == _T_23 ? ram_374 : _GEN_8776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8778 = 10'h177 == _T_23 ? ram_375 : _GEN_8777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8779 = 10'h178 == _T_23 ? ram_376 : _GEN_8778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8780 = 10'h179 == _T_23 ? ram_377 : _GEN_8779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8781 = 10'h17a == _T_23 ? ram_378 : _GEN_8780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8782 = 10'h17b == _T_23 ? ram_379 : _GEN_8781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8783 = 10'h17c == _T_23 ? ram_380 : _GEN_8782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8784 = 10'h17d == _T_23 ? ram_381 : _GEN_8783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8785 = 10'h17e == _T_23 ? ram_382 : _GEN_8784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8786 = 10'h17f == _T_23 ? ram_383 : _GEN_8785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8787 = 10'h180 == _T_23 ? ram_384 : _GEN_8786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8788 = 10'h181 == _T_23 ? ram_385 : _GEN_8787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8789 = 10'h182 == _T_23 ? ram_386 : _GEN_8788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8790 = 10'h183 == _T_23 ? ram_387 : _GEN_8789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8791 = 10'h184 == _T_23 ? ram_388 : _GEN_8790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8792 = 10'h185 == _T_23 ? ram_389 : _GEN_8791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8793 = 10'h186 == _T_23 ? ram_390 : _GEN_8792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8794 = 10'h187 == _T_23 ? ram_391 : _GEN_8793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8795 = 10'h188 == _T_23 ? ram_392 : _GEN_8794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8796 = 10'h189 == _T_23 ? ram_393 : _GEN_8795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8797 = 10'h18a == _T_23 ? ram_394 : _GEN_8796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8798 = 10'h18b == _T_23 ? ram_395 : _GEN_8797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8799 = 10'h18c == _T_23 ? ram_396 : _GEN_8798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8800 = 10'h18d == _T_23 ? ram_397 : _GEN_8799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8801 = 10'h18e == _T_23 ? ram_398 : _GEN_8800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8802 = 10'h18f == _T_23 ? ram_399 : _GEN_8801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8803 = 10'h190 == _T_23 ? ram_400 : _GEN_8802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8804 = 10'h191 == _T_23 ? ram_401 : _GEN_8803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8805 = 10'h192 == _T_23 ? ram_402 : _GEN_8804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8806 = 10'h193 == _T_23 ? ram_403 : _GEN_8805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8807 = 10'h194 == _T_23 ? ram_404 : _GEN_8806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8808 = 10'h195 == _T_23 ? ram_405 : _GEN_8807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8809 = 10'h196 == _T_23 ? ram_406 : _GEN_8808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8810 = 10'h197 == _T_23 ? ram_407 : _GEN_8809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8811 = 10'h198 == _T_23 ? ram_408 : _GEN_8810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8812 = 10'h199 == _T_23 ? ram_409 : _GEN_8811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8813 = 10'h19a == _T_23 ? ram_410 : _GEN_8812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8814 = 10'h19b == _T_23 ? ram_411 : _GEN_8813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8815 = 10'h19c == _T_23 ? ram_412 : _GEN_8814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8816 = 10'h19d == _T_23 ? ram_413 : _GEN_8815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8817 = 10'h19e == _T_23 ? ram_414 : _GEN_8816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8818 = 10'h19f == _T_23 ? ram_415 : _GEN_8817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8819 = 10'h1a0 == _T_23 ? ram_416 : _GEN_8818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8820 = 10'h1a1 == _T_23 ? ram_417 : _GEN_8819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8821 = 10'h1a2 == _T_23 ? ram_418 : _GEN_8820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8822 = 10'h1a3 == _T_23 ? ram_419 : _GEN_8821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8823 = 10'h1a4 == _T_23 ? ram_420 : _GEN_8822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8824 = 10'h1a5 == _T_23 ? ram_421 : _GEN_8823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8825 = 10'h1a6 == _T_23 ? ram_422 : _GEN_8824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8826 = 10'h1a7 == _T_23 ? ram_423 : _GEN_8825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8827 = 10'h1a8 == _T_23 ? ram_424 : _GEN_8826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8828 = 10'h1a9 == _T_23 ? ram_425 : _GEN_8827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8829 = 10'h1aa == _T_23 ? ram_426 : _GEN_8828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8830 = 10'h1ab == _T_23 ? ram_427 : _GEN_8829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8831 = 10'h1ac == _T_23 ? ram_428 : _GEN_8830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8832 = 10'h1ad == _T_23 ? ram_429 : _GEN_8831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8833 = 10'h1ae == _T_23 ? ram_430 : _GEN_8832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8834 = 10'h1af == _T_23 ? ram_431 : _GEN_8833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8835 = 10'h1b0 == _T_23 ? ram_432 : _GEN_8834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8836 = 10'h1b1 == _T_23 ? ram_433 : _GEN_8835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8837 = 10'h1b2 == _T_23 ? ram_434 : _GEN_8836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8838 = 10'h1b3 == _T_23 ? ram_435 : _GEN_8837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8839 = 10'h1b4 == _T_23 ? ram_436 : _GEN_8838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8840 = 10'h1b5 == _T_23 ? ram_437 : _GEN_8839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8841 = 10'h1b6 == _T_23 ? ram_438 : _GEN_8840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8842 = 10'h1b7 == _T_23 ? ram_439 : _GEN_8841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8843 = 10'h1b8 == _T_23 ? ram_440 : _GEN_8842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8844 = 10'h1b9 == _T_23 ? ram_441 : _GEN_8843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8845 = 10'h1ba == _T_23 ? ram_442 : _GEN_8844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8846 = 10'h1bb == _T_23 ? ram_443 : _GEN_8845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8847 = 10'h1bc == _T_23 ? ram_444 : _GEN_8846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8848 = 10'h1bd == _T_23 ? ram_445 : _GEN_8847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8849 = 10'h1be == _T_23 ? ram_446 : _GEN_8848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8850 = 10'h1bf == _T_23 ? ram_447 : _GEN_8849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8851 = 10'h1c0 == _T_23 ? ram_448 : _GEN_8850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8852 = 10'h1c1 == _T_23 ? ram_449 : _GEN_8851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8853 = 10'h1c2 == _T_23 ? ram_450 : _GEN_8852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8854 = 10'h1c3 == _T_23 ? ram_451 : _GEN_8853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8855 = 10'h1c4 == _T_23 ? ram_452 : _GEN_8854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8856 = 10'h1c5 == _T_23 ? ram_453 : _GEN_8855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8857 = 10'h1c6 == _T_23 ? ram_454 : _GEN_8856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8858 = 10'h1c7 == _T_23 ? ram_455 : _GEN_8857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8859 = 10'h1c8 == _T_23 ? ram_456 : _GEN_8858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8860 = 10'h1c9 == _T_23 ? ram_457 : _GEN_8859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8861 = 10'h1ca == _T_23 ? ram_458 : _GEN_8860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8862 = 10'h1cb == _T_23 ? ram_459 : _GEN_8861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8863 = 10'h1cc == _T_23 ? ram_460 : _GEN_8862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8864 = 10'h1cd == _T_23 ? ram_461 : _GEN_8863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8865 = 10'h1ce == _T_23 ? ram_462 : _GEN_8864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8866 = 10'h1cf == _T_23 ? ram_463 : _GEN_8865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8867 = 10'h1d0 == _T_23 ? ram_464 : _GEN_8866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8868 = 10'h1d1 == _T_23 ? ram_465 : _GEN_8867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8869 = 10'h1d2 == _T_23 ? ram_466 : _GEN_8868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8870 = 10'h1d3 == _T_23 ? ram_467 : _GEN_8869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8871 = 10'h1d4 == _T_23 ? ram_468 : _GEN_8870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8872 = 10'h1d5 == _T_23 ? ram_469 : _GEN_8871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8873 = 10'h1d6 == _T_23 ? ram_470 : _GEN_8872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8874 = 10'h1d7 == _T_23 ? ram_471 : _GEN_8873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8875 = 10'h1d8 == _T_23 ? ram_472 : _GEN_8874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8876 = 10'h1d9 == _T_23 ? ram_473 : _GEN_8875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8877 = 10'h1da == _T_23 ? ram_474 : _GEN_8876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8878 = 10'h1db == _T_23 ? ram_475 : _GEN_8877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8879 = 10'h1dc == _T_23 ? ram_476 : _GEN_8878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8880 = 10'h1dd == _T_23 ? ram_477 : _GEN_8879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8881 = 10'h1de == _T_23 ? ram_478 : _GEN_8880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8882 = 10'h1df == _T_23 ? ram_479 : _GEN_8881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8883 = 10'h1e0 == _T_23 ? ram_480 : _GEN_8882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8884 = 10'h1e1 == _T_23 ? ram_481 : _GEN_8883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8885 = 10'h1e2 == _T_23 ? ram_482 : _GEN_8884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8886 = 10'h1e3 == _T_23 ? ram_483 : _GEN_8885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8887 = 10'h1e4 == _T_23 ? ram_484 : _GEN_8886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8888 = 10'h1e5 == _T_23 ? ram_485 : _GEN_8887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8889 = 10'h1e6 == _T_23 ? ram_486 : _GEN_8888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8890 = 10'h1e7 == _T_23 ? ram_487 : _GEN_8889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8891 = 10'h1e8 == _T_23 ? ram_488 : _GEN_8890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8892 = 10'h1e9 == _T_23 ? ram_489 : _GEN_8891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8893 = 10'h1ea == _T_23 ? ram_490 : _GEN_8892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8894 = 10'h1eb == _T_23 ? ram_491 : _GEN_8893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8895 = 10'h1ec == _T_23 ? ram_492 : _GEN_8894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8896 = 10'h1ed == _T_23 ? ram_493 : _GEN_8895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8897 = 10'h1ee == _T_23 ? ram_494 : _GEN_8896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8898 = 10'h1ef == _T_23 ? ram_495 : _GEN_8897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8899 = 10'h1f0 == _T_23 ? ram_496 : _GEN_8898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8900 = 10'h1f1 == _T_23 ? ram_497 : _GEN_8899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8901 = 10'h1f2 == _T_23 ? ram_498 : _GEN_8900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8902 = 10'h1f3 == _T_23 ? ram_499 : _GEN_8901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8903 = 10'h1f4 == _T_23 ? ram_500 : _GEN_8902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8904 = 10'h1f5 == _T_23 ? ram_501 : _GEN_8903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8905 = 10'h1f6 == _T_23 ? ram_502 : _GEN_8904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8906 = 10'h1f7 == _T_23 ? ram_503 : _GEN_8905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8907 = 10'h1f8 == _T_23 ? ram_504 : _GEN_8906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8908 = 10'h1f9 == _T_23 ? ram_505 : _GEN_8907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8909 = 10'h1fa == _T_23 ? ram_506 : _GEN_8908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8910 = 10'h1fb == _T_23 ? ram_507 : _GEN_8909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8911 = 10'h1fc == _T_23 ? ram_508 : _GEN_8910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8912 = 10'h1fd == _T_23 ? ram_509 : _GEN_8911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8913 = 10'h1fe == _T_23 ? ram_510 : _GEN_8912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8914 = 10'h1ff == _T_23 ? ram_511 : _GEN_8913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8915 = 10'h200 == _T_23 ? ram_512 : _GEN_8914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8916 = 10'h201 == _T_23 ? ram_513 : _GEN_8915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8917 = 10'h202 == _T_23 ? ram_514 : _GEN_8916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8918 = 10'h203 == _T_23 ? ram_515 : _GEN_8917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8919 = 10'h204 == _T_23 ? ram_516 : _GEN_8918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8920 = 10'h205 == _T_23 ? ram_517 : _GEN_8919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8921 = 10'h206 == _T_23 ? ram_518 : _GEN_8920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8922 = 10'h207 == _T_23 ? ram_519 : _GEN_8921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8923 = 10'h208 == _T_23 ? ram_520 : _GEN_8922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8924 = 10'h209 == _T_23 ? ram_521 : _GEN_8923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8925 = 10'h20a == _T_23 ? ram_522 : _GEN_8924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8926 = 10'h20b == _T_23 ? ram_523 : _GEN_8925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_8927 = 10'h20c == _T_23 ? ram_524 : _GEN_8926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19077 = {{8190'd0}, _GEN_8927}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_233 = _GEN_19077 ^ _ram_T_232; // @[vga.scala 64:41]
  wire [287:0] _GEN_8928 = 10'h0 == _T_23 ? _ram_T_233[287:0] : _GEN_7878; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8929 = 10'h1 == _T_23 ? _ram_T_233[287:0] : _GEN_7879; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8930 = 10'h2 == _T_23 ? _ram_T_233[287:0] : _GEN_7880; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8931 = 10'h3 == _T_23 ? _ram_T_233[287:0] : _GEN_7881; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8932 = 10'h4 == _T_23 ? _ram_T_233[287:0] : _GEN_7882; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8933 = 10'h5 == _T_23 ? _ram_T_233[287:0] : _GEN_7883; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8934 = 10'h6 == _T_23 ? _ram_T_233[287:0] : _GEN_7884; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8935 = 10'h7 == _T_23 ? _ram_T_233[287:0] : _GEN_7885; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8936 = 10'h8 == _T_23 ? _ram_T_233[287:0] : _GEN_7886; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8937 = 10'h9 == _T_23 ? _ram_T_233[287:0] : _GEN_7887; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8938 = 10'ha == _T_23 ? _ram_T_233[287:0] : _GEN_7888; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8939 = 10'hb == _T_23 ? _ram_T_233[287:0] : _GEN_7889; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8940 = 10'hc == _T_23 ? _ram_T_233[287:0] : _GEN_7890; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8941 = 10'hd == _T_23 ? _ram_T_233[287:0] : _GEN_7891; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8942 = 10'he == _T_23 ? _ram_T_233[287:0] : _GEN_7892; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8943 = 10'hf == _T_23 ? _ram_T_233[287:0] : _GEN_7893; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8944 = 10'h10 == _T_23 ? _ram_T_233[287:0] : _GEN_7894; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8945 = 10'h11 == _T_23 ? _ram_T_233[287:0] : _GEN_7895; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8946 = 10'h12 == _T_23 ? _ram_T_233[287:0] : _GEN_7896; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8947 = 10'h13 == _T_23 ? _ram_T_233[287:0] : _GEN_7897; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8948 = 10'h14 == _T_23 ? _ram_T_233[287:0] : _GEN_7898; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8949 = 10'h15 == _T_23 ? _ram_T_233[287:0] : _GEN_7899; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8950 = 10'h16 == _T_23 ? _ram_T_233[287:0] : _GEN_7900; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8951 = 10'h17 == _T_23 ? _ram_T_233[287:0] : _GEN_7901; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8952 = 10'h18 == _T_23 ? _ram_T_233[287:0] : _GEN_7902; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8953 = 10'h19 == _T_23 ? _ram_T_233[287:0] : _GEN_7903; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8954 = 10'h1a == _T_23 ? _ram_T_233[287:0] : _GEN_7904; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8955 = 10'h1b == _T_23 ? _ram_T_233[287:0] : _GEN_7905; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8956 = 10'h1c == _T_23 ? _ram_T_233[287:0] : _GEN_7906; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8957 = 10'h1d == _T_23 ? _ram_T_233[287:0] : _GEN_7907; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8958 = 10'h1e == _T_23 ? _ram_T_233[287:0] : _GEN_7908; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8959 = 10'h1f == _T_23 ? _ram_T_233[287:0] : _GEN_7909; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8960 = 10'h20 == _T_23 ? _ram_T_233[287:0] : _GEN_7910; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8961 = 10'h21 == _T_23 ? _ram_T_233[287:0] : _GEN_7911; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8962 = 10'h22 == _T_23 ? _ram_T_233[287:0] : _GEN_7912; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8963 = 10'h23 == _T_23 ? _ram_T_233[287:0] : _GEN_7913; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8964 = 10'h24 == _T_23 ? _ram_T_233[287:0] : _GEN_7914; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8965 = 10'h25 == _T_23 ? _ram_T_233[287:0] : _GEN_7915; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8966 = 10'h26 == _T_23 ? _ram_T_233[287:0] : _GEN_7916; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8967 = 10'h27 == _T_23 ? _ram_T_233[287:0] : _GEN_7917; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8968 = 10'h28 == _T_23 ? _ram_T_233[287:0] : _GEN_7918; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8969 = 10'h29 == _T_23 ? _ram_T_233[287:0] : _GEN_7919; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8970 = 10'h2a == _T_23 ? _ram_T_233[287:0] : _GEN_7920; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8971 = 10'h2b == _T_23 ? _ram_T_233[287:0] : _GEN_7921; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8972 = 10'h2c == _T_23 ? _ram_T_233[287:0] : _GEN_7922; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8973 = 10'h2d == _T_23 ? _ram_T_233[287:0] : _GEN_7923; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8974 = 10'h2e == _T_23 ? _ram_T_233[287:0] : _GEN_7924; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8975 = 10'h2f == _T_23 ? _ram_T_233[287:0] : _GEN_7925; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8976 = 10'h30 == _T_23 ? _ram_T_233[287:0] : _GEN_7926; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8977 = 10'h31 == _T_23 ? _ram_T_233[287:0] : _GEN_7927; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8978 = 10'h32 == _T_23 ? _ram_T_233[287:0] : _GEN_7928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8979 = 10'h33 == _T_23 ? _ram_T_233[287:0] : _GEN_7929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8980 = 10'h34 == _T_23 ? _ram_T_233[287:0] : _GEN_7930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8981 = 10'h35 == _T_23 ? _ram_T_233[287:0] : _GEN_7931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8982 = 10'h36 == _T_23 ? _ram_T_233[287:0] : _GEN_7932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8983 = 10'h37 == _T_23 ? _ram_T_233[287:0] : _GEN_7933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8984 = 10'h38 == _T_23 ? _ram_T_233[287:0] : _GEN_7934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8985 = 10'h39 == _T_23 ? _ram_T_233[287:0] : _GEN_7935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8986 = 10'h3a == _T_23 ? _ram_T_233[287:0] : _GEN_7936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8987 = 10'h3b == _T_23 ? _ram_T_233[287:0] : _GEN_7937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8988 = 10'h3c == _T_23 ? _ram_T_233[287:0] : _GEN_7938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8989 = 10'h3d == _T_23 ? _ram_T_233[287:0] : _GEN_7939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8990 = 10'h3e == _T_23 ? _ram_T_233[287:0] : _GEN_7940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8991 = 10'h3f == _T_23 ? _ram_T_233[287:0] : _GEN_7941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8992 = 10'h40 == _T_23 ? _ram_T_233[287:0] : _GEN_7942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8993 = 10'h41 == _T_23 ? _ram_T_233[287:0] : _GEN_7943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8994 = 10'h42 == _T_23 ? _ram_T_233[287:0] : _GEN_7944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8995 = 10'h43 == _T_23 ? _ram_T_233[287:0] : _GEN_7945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8996 = 10'h44 == _T_23 ? _ram_T_233[287:0] : _GEN_7946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8997 = 10'h45 == _T_23 ? _ram_T_233[287:0] : _GEN_7947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8998 = 10'h46 == _T_23 ? _ram_T_233[287:0] : _GEN_7948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_8999 = 10'h47 == _T_23 ? _ram_T_233[287:0] : _GEN_7949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9000 = 10'h48 == _T_23 ? _ram_T_233[287:0] : _GEN_7950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9001 = 10'h49 == _T_23 ? _ram_T_233[287:0] : _GEN_7951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9002 = 10'h4a == _T_23 ? _ram_T_233[287:0] : _GEN_7952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9003 = 10'h4b == _T_23 ? _ram_T_233[287:0] : _GEN_7953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9004 = 10'h4c == _T_23 ? _ram_T_233[287:0] : _GEN_7954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9005 = 10'h4d == _T_23 ? _ram_T_233[287:0] : _GEN_7955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9006 = 10'h4e == _T_23 ? _ram_T_233[287:0] : _GEN_7956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9007 = 10'h4f == _T_23 ? _ram_T_233[287:0] : _GEN_7957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9008 = 10'h50 == _T_23 ? _ram_T_233[287:0] : _GEN_7958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9009 = 10'h51 == _T_23 ? _ram_T_233[287:0] : _GEN_7959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9010 = 10'h52 == _T_23 ? _ram_T_233[287:0] : _GEN_7960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9011 = 10'h53 == _T_23 ? _ram_T_233[287:0] : _GEN_7961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9012 = 10'h54 == _T_23 ? _ram_T_233[287:0] : _GEN_7962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9013 = 10'h55 == _T_23 ? _ram_T_233[287:0] : _GEN_7963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9014 = 10'h56 == _T_23 ? _ram_T_233[287:0] : _GEN_7964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9015 = 10'h57 == _T_23 ? _ram_T_233[287:0] : _GEN_7965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9016 = 10'h58 == _T_23 ? _ram_T_233[287:0] : _GEN_7966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9017 = 10'h59 == _T_23 ? _ram_T_233[287:0] : _GEN_7967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9018 = 10'h5a == _T_23 ? _ram_T_233[287:0] : _GEN_7968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9019 = 10'h5b == _T_23 ? _ram_T_233[287:0] : _GEN_7969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9020 = 10'h5c == _T_23 ? _ram_T_233[287:0] : _GEN_7970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9021 = 10'h5d == _T_23 ? _ram_T_233[287:0] : _GEN_7971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9022 = 10'h5e == _T_23 ? _ram_T_233[287:0] : _GEN_7972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9023 = 10'h5f == _T_23 ? _ram_T_233[287:0] : _GEN_7973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9024 = 10'h60 == _T_23 ? _ram_T_233[287:0] : _GEN_7974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9025 = 10'h61 == _T_23 ? _ram_T_233[287:0] : _GEN_7975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9026 = 10'h62 == _T_23 ? _ram_T_233[287:0] : _GEN_7976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9027 = 10'h63 == _T_23 ? _ram_T_233[287:0] : _GEN_7977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9028 = 10'h64 == _T_23 ? _ram_T_233[287:0] : _GEN_7978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9029 = 10'h65 == _T_23 ? _ram_T_233[287:0] : _GEN_7979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9030 = 10'h66 == _T_23 ? _ram_T_233[287:0] : _GEN_7980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9031 = 10'h67 == _T_23 ? _ram_T_233[287:0] : _GEN_7981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9032 = 10'h68 == _T_23 ? _ram_T_233[287:0] : _GEN_7982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9033 = 10'h69 == _T_23 ? _ram_T_233[287:0] : _GEN_7983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9034 = 10'h6a == _T_23 ? _ram_T_233[287:0] : _GEN_7984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9035 = 10'h6b == _T_23 ? _ram_T_233[287:0] : _GEN_7985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9036 = 10'h6c == _T_23 ? _ram_T_233[287:0] : _GEN_7986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9037 = 10'h6d == _T_23 ? _ram_T_233[287:0] : _GEN_7987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9038 = 10'h6e == _T_23 ? _ram_T_233[287:0] : _GEN_7988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9039 = 10'h6f == _T_23 ? _ram_T_233[287:0] : _GEN_7989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9040 = 10'h70 == _T_23 ? _ram_T_233[287:0] : _GEN_7990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9041 = 10'h71 == _T_23 ? _ram_T_233[287:0] : _GEN_7991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9042 = 10'h72 == _T_23 ? _ram_T_233[287:0] : _GEN_7992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9043 = 10'h73 == _T_23 ? _ram_T_233[287:0] : _GEN_7993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9044 = 10'h74 == _T_23 ? _ram_T_233[287:0] : _GEN_7994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9045 = 10'h75 == _T_23 ? _ram_T_233[287:0] : _GEN_7995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9046 = 10'h76 == _T_23 ? _ram_T_233[287:0] : _GEN_7996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9047 = 10'h77 == _T_23 ? _ram_T_233[287:0] : _GEN_7997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9048 = 10'h78 == _T_23 ? _ram_T_233[287:0] : _GEN_7998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9049 = 10'h79 == _T_23 ? _ram_T_233[287:0] : _GEN_7999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9050 = 10'h7a == _T_23 ? _ram_T_233[287:0] : _GEN_8000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9051 = 10'h7b == _T_23 ? _ram_T_233[287:0] : _GEN_8001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9052 = 10'h7c == _T_23 ? _ram_T_233[287:0] : _GEN_8002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9053 = 10'h7d == _T_23 ? _ram_T_233[287:0] : _GEN_8003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9054 = 10'h7e == _T_23 ? _ram_T_233[287:0] : _GEN_8004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9055 = 10'h7f == _T_23 ? _ram_T_233[287:0] : _GEN_8005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9056 = 10'h80 == _T_23 ? _ram_T_233[287:0] : _GEN_8006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9057 = 10'h81 == _T_23 ? _ram_T_233[287:0] : _GEN_8007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9058 = 10'h82 == _T_23 ? _ram_T_233[287:0] : _GEN_8008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9059 = 10'h83 == _T_23 ? _ram_T_233[287:0] : _GEN_8009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9060 = 10'h84 == _T_23 ? _ram_T_233[287:0] : _GEN_8010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9061 = 10'h85 == _T_23 ? _ram_T_233[287:0] : _GEN_8011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9062 = 10'h86 == _T_23 ? _ram_T_233[287:0] : _GEN_8012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9063 = 10'h87 == _T_23 ? _ram_T_233[287:0] : _GEN_8013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9064 = 10'h88 == _T_23 ? _ram_T_233[287:0] : _GEN_8014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9065 = 10'h89 == _T_23 ? _ram_T_233[287:0] : _GEN_8015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9066 = 10'h8a == _T_23 ? _ram_T_233[287:0] : _GEN_8016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9067 = 10'h8b == _T_23 ? _ram_T_233[287:0] : _GEN_8017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9068 = 10'h8c == _T_23 ? _ram_T_233[287:0] : _GEN_8018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9069 = 10'h8d == _T_23 ? _ram_T_233[287:0] : _GEN_8019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9070 = 10'h8e == _T_23 ? _ram_T_233[287:0] : _GEN_8020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9071 = 10'h8f == _T_23 ? _ram_T_233[287:0] : _GEN_8021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9072 = 10'h90 == _T_23 ? _ram_T_233[287:0] : _GEN_8022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9073 = 10'h91 == _T_23 ? _ram_T_233[287:0] : _GEN_8023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9074 = 10'h92 == _T_23 ? _ram_T_233[287:0] : _GEN_8024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9075 = 10'h93 == _T_23 ? _ram_T_233[287:0] : _GEN_8025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9076 = 10'h94 == _T_23 ? _ram_T_233[287:0] : _GEN_8026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9077 = 10'h95 == _T_23 ? _ram_T_233[287:0] : _GEN_8027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9078 = 10'h96 == _T_23 ? _ram_T_233[287:0] : _GEN_8028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9079 = 10'h97 == _T_23 ? _ram_T_233[287:0] : _GEN_8029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9080 = 10'h98 == _T_23 ? _ram_T_233[287:0] : _GEN_8030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9081 = 10'h99 == _T_23 ? _ram_T_233[287:0] : _GEN_8031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9082 = 10'h9a == _T_23 ? _ram_T_233[287:0] : _GEN_8032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9083 = 10'h9b == _T_23 ? _ram_T_233[287:0] : _GEN_8033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9084 = 10'h9c == _T_23 ? _ram_T_233[287:0] : _GEN_8034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9085 = 10'h9d == _T_23 ? _ram_T_233[287:0] : _GEN_8035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9086 = 10'h9e == _T_23 ? _ram_T_233[287:0] : _GEN_8036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9087 = 10'h9f == _T_23 ? _ram_T_233[287:0] : _GEN_8037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9088 = 10'ha0 == _T_23 ? _ram_T_233[287:0] : _GEN_8038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9089 = 10'ha1 == _T_23 ? _ram_T_233[287:0] : _GEN_8039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9090 = 10'ha2 == _T_23 ? _ram_T_233[287:0] : _GEN_8040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9091 = 10'ha3 == _T_23 ? _ram_T_233[287:0] : _GEN_8041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9092 = 10'ha4 == _T_23 ? _ram_T_233[287:0] : _GEN_8042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9093 = 10'ha5 == _T_23 ? _ram_T_233[287:0] : _GEN_8043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9094 = 10'ha6 == _T_23 ? _ram_T_233[287:0] : _GEN_8044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9095 = 10'ha7 == _T_23 ? _ram_T_233[287:0] : _GEN_8045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9096 = 10'ha8 == _T_23 ? _ram_T_233[287:0] : _GEN_8046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9097 = 10'ha9 == _T_23 ? _ram_T_233[287:0] : _GEN_8047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9098 = 10'haa == _T_23 ? _ram_T_233[287:0] : _GEN_8048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9099 = 10'hab == _T_23 ? _ram_T_233[287:0] : _GEN_8049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9100 = 10'hac == _T_23 ? _ram_T_233[287:0] : _GEN_8050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9101 = 10'had == _T_23 ? _ram_T_233[287:0] : _GEN_8051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9102 = 10'hae == _T_23 ? _ram_T_233[287:0] : _GEN_8052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9103 = 10'haf == _T_23 ? _ram_T_233[287:0] : _GEN_8053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9104 = 10'hb0 == _T_23 ? _ram_T_233[287:0] : _GEN_8054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9105 = 10'hb1 == _T_23 ? _ram_T_233[287:0] : _GEN_8055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9106 = 10'hb2 == _T_23 ? _ram_T_233[287:0] : _GEN_8056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9107 = 10'hb3 == _T_23 ? _ram_T_233[287:0] : _GEN_8057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9108 = 10'hb4 == _T_23 ? _ram_T_233[287:0] : _GEN_8058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9109 = 10'hb5 == _T_23 ? _ram_T_233[287:0] : _GEN_8059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9110 = 10'hb6 == _T_23 ? _ram_T_233[287:0] : _GEN_8060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9111 = 10'hb7 == _T_23 ? _ram_T_233[287:0] : _GEN_8061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9112 = 10'hb8 == _T_23 ? _ram_T_233[287:0] : _GEN_8062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9113 = 10'hb9 == _T_23 ? _ram_T_233[287:0] : _GEN_8063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9114 = 10'hba == _T_23 ? _ram_T_233[287:0] : _GEN_8064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9115 = 10'hbb == _T_23 ? _ram_T_233[287:0] : _GEN_8065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9116 = 10'hbc == _T_23 ? _ram_T_233[287:0] : _GEN_8066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9117 = 10'hbd == _T_23 ? _ram_T_233[287:0] : _GEN_8067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9118 = 10'hbe == _T_23 ? _ram_T_233[287:0] : _GEN_8068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9119 = 10'hbf == _T_23 ? _ram_T_233[287:0] : _GEN_8069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9120 = 10'hc0 == _T_23 ? _ram_T_233[287:0] : _GEN_8070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9121 = 10'hc1 == _T_23 ? _ram_T_233[287:0] : _GEN_8071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9122 = 10'hc2 == _T_23 ? _ram_T_233[287:0] : _GEN_8072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9123 = 10'hc3 == _T_23 ? _ram_T_233[287:0] : _GEN_8073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9124 = 10'hc4 == _T_23 ? _ram_T_233[287:0] : _GEN_8074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9125 = 10'hc5 == _T_23 ? _ram_T_233[287:0] : _GEN_8075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9126 = 10'hc6 == _T_23 ? _ram_T_233[287:0] : _GEN_8076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9127 = 10'hc7 == _T_23 ? _ram_T_233[287:0] : _GEN_8077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9128 = 10'hc8 == _T_23 ? _ram_T_233[287:0] : _GEN_8078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9129 = 10'hc9 == _T_23 ? _ram_T_233[287:0] : _GEN_8079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9130 = 10'hca == _T_23 ? _ram_T_233[287:0] : _GEN_8080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9131 = 10'hcb == _T_23 ? _ram_T_233[287:0] : _GEN_8081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9132 = 10'hcc == _T_23 ? _ram_T_233[287:0] : _GEN_8082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9133 = 10'hcd == _T_23 ? _ram_T_233[287:0] : _GEN_8083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9134 = 10'hce == _T_23 ? _ram_T_233[287:0] : _GEN_8084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9135 = 10'hcf == _T_23 ? _ram_T_233[287:0] : _GEN_8085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9136 = 10'hd0 == _T_23 ? _ram_T_233[287:0] : _GEN_8086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9137 = 10'hd1 == _T_23 ? _ram_T_233[287:0] : _GEN_8087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9138 = 10'hd2 == _T_23 ? _ram_T_233[287:0] : _GEN_8088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9139 = 10'hd3 == _T_23 ? _ram_T_233[287:0] : _GEN_8089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9140 = 10'hd4 == _T_23 ? _ram_T_233[287:0] : _GEN_8090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9141 = 10'hd5 == _T_23 ? _ram_T_233[287:0] : _GEN_8091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9142 = 10'hd6 == _T_23 ? _ram_T_233[287:0] : _GEN_8092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9143 = 10'hd7 == _T_23 ? _ram_T_233[287:0] : _GEN_8093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9144 = 10'hd8 == _T_23 ? _ram_T_233[287:0] : _GEN_8094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9145 = 10'hd9 == _T_23 ? _ram_T_233[287:0] : _GEN_8095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9146 = 10'hda == _T_23 ? _ram_T_233[287:0] : _GEN_8096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9147 = 10'hdb == _T_23 ? _ram_T_233[287:0] : _GEN_8097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9148 = 10'hdc == _T_23 ? _ram_T_233[287:0] : _GEN_8098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9149 = 10'hdd == _T_23 ? _ram_T_233[287:0] : _GEN_8099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9150 = 10'hde == _T_23 ? _ram_T_233[287:0] : _GEN_8100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9151 = 10'hdf == _T_23 ? _ram_T_233[287:0] : _GEN_8101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9152 = 10'he0 == _T_23 ? _ram_T_233[287:0] : _GEN_8102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9153 = 10'he1 == _T_23 ? _ram_T_233[287:0] : _GEN_8103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9154 = 10'he2 == _T_23 ? _ram_T_233[287:0] : _GEN_8104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9155 = 10'he3 == _T_23 ? _ram_T_233[287:0] : _GEN_8105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9156 = 10'he4 == _T_23 ? _ram_T_233[287:0] : _GEN_8106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9157 = 10'he5 == _T_23 ? _ram_T_233[287:0] : _GEN_8107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9158 = 10'he6 == _T_23 ? _ram_T_233[287:0] : _GEN_8108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9159 = 10'he7 == _T_23 ? _ram_T_233[287:0] : _GEN_8109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9160 = 10'he8 == _T_23 ? _ram_T_233[287:0] : _GEN_8110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9161 = 10'he9 == _T_23 ? _ram_T_233[287:0] : _GEN_8111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9162 = 10'hea == _T_23 ? _ram_T_233[287:0] : _GEN_8112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9163 = 10'heb == _T_23 ? _ram_T_233[287:0] : _GEN_8113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9164 = 10'hec == _T_23 ? _ram_T_233[287:0] : _GEN_8114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9165 = 10'hed == _T_23 ? _ram_T_233[287:0] : _GEN_8115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9166 = 10'hee == _T_23 ? _ram_T_233[287:0] : _GEN_8116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9167 = 10'hef == _T_23 ? _ram_T_233[287:0] : _GEN_8117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9168 = 10'hf0 == _T_23 ? _ram_T_233[287:0] : _GEN_8118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9169 = 10'hf1 == _T_23 ? _ram_T_233[287:0] : _GEN_8119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9170 = 10'hf2 == _T_23 ? _ram_T_233[287:0] : _GEN_8120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9171 = 10'hf3 == _T_23 ? _ram_T_233[287:0] : _GEN_8121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9172 = 10'hf4 == _T_23 ? _ram_T_233[287:0] : _GEN_8122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9173 = 10'hf5 == _T_23 ? _ram_T_233[287:0] : _GEN_8123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9174 = 10'hf6 == _T_23 ? _ram_T_233[287:0] : _GEN_8124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9175 = 10'hf7 == _T_23 ? _ram_T_233[287:0] : _GEN_8125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9176 = 10'hf8 == _T_23 ? _ram_T_233[287:0] : _GEN_8126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9177 = 10'hf9 == _T_23 ? _ram_T_233[287:0] : _GEN_8127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9178 = 10'hfa == _T_23 ? _ram_T_233[287:0] : _GEN_8128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9179 = 10'hfb == _T_23 ? _ram_T_233[287:0] : _GEN_8129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9180 = 10'hfc == _T_23 ? _ram_T_233[287:0] : _GEN_8130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9181 = 10'hfd == _T_23 ? _ram_T_233[287:0] : _GEN_8131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9182 = 10'hfe == _T_23 ? _ram_T_233[287:0] : _GEN_8132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9183 = 10'hff == _T_23 ? _ram_T_233[287:0] : _GEN_8133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9184 = 10'h100 == _T_23 ? _ram_T_233[287:0] : _GEN_8134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9185 = 10'h101 == _T_23 ? _ram_T_233[287:0] : _GEN_8135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9186 = 10'h102 == _T_23 ? _ram_T_233[287:0] : _GEN_8136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9187 = 10'h103 == _T_23 ? _ram_T_233[287:0] : _GEN_8137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9188 = 10'h104 == _T_23 ? _ram_T_233[287:0] : _GEN_8138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9189 = 10'h105 == _T_23 ? _ram_T_233[287:0] : _GEN_8139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9190 = 10'h106 == _T_23 ? _ram_T_233[287:0] : _GEN_8140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9191 = 10'h107 == _T_23 ? _ram_T_233[287:0] : _GEN_8141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9192 = 10'h108 == _T_23 ? _ram_T_233[287:0] : _GEN_8142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9193 = 10'h109 == _T_23 ? _ram_T_233[287:0] : _GEN_8143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9194 = 10'h10a == _T_23 ? _ram_T_233[287:0] : _GEN_8144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9195 = 10'h10b == _T_23 ? _ram_T_233[287:0] : _GEN_8145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9196 = 10'h10c == _T_23 ? _ram_T_233[287:0] : _GEN_8146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9197 = 10'h10d == _T_23 ? _ram_T_233[287:0] : _GEN_8147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9198 = 10'h10e == _T_23 ? _ram_T_233[287:0] : _GEN_8148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9199 = 10'h10f == _T_23 ? _ram_T_233[287:0] : _GEN_8149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9200 = 10'h110 == _T_23 ? _ram_T_233[287:0] : _GEN_8150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9201 = 10'h111 == _T_23 ? _ram_T_233[287:0] : _GEN_8151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9202 = 10'h112 == _T_23 ? _ram_T_233[287:0] : _GEN_8152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9203 = 10'h113 == _T_23 ? _ram_T_233[287:0] : _GEN_8153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9204 = 10'h114 == _T_23 ? _ram_T_233[287:0] : _GEN_8154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9205 = 10'h115 == _T_23 ? _ram_T_233[287:0] : _GEN_8155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9206 = 10'h116 == _T_23 ? _ram_T_233[287:0] : _GEN_8156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9207 = 10'h117 == _T_23 ? _ram_T_233[287:0] : _GEN_8157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9208 = 10'h118 == _T_23 ? _ram_T_233[287:0] : _GEN_8158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9209 = 10'h119 == _T_23 ? _ram_T_233[287:0] : _GEN_8159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9210 = 10'h11a == _T_23 ? _ram_T_233[287:0] : _GEN_8160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9211 = 10'h11b == _T_23 ? _ram_T_233[287:0] : _GEN_8161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9212 = 10'h11c == _T_23 ? _ram_T_233[287:0] : _GEN_8162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9213 = 10'h11d == _T_23 ? _ram_T_233[287:0] : _GEN_8163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9214 = 10'h11e == _T_23 ? _ram_T_233[287:0] : _GEN_8164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9215 = 10'h11f == _T_23 ? _ram_T_233[287:0] : _GEN_8165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9216 = 10'h120 == _T_23 ? _ram_T_233[287:0] : _GEN_8166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9217 = 10'h121 == _T_23 ? _ram_T_233[287:0] : _GEN_8167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9218 = 10'h122 == _T_23 ? _ram_T_233[287:0] : _GEN_8168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9219 = 10'h123 == _T_23 ? _ram_T_233[287:0] : _GEN_8169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9220 = 10'h124 == _T_23 ? _ram_T_233[287:0] : _GEN_8170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9221 = 10'h125 == _T_23 ? _ram_T_233[287:0] : _GEN_8171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9222 = 10'h126 == _T_23 ? _ram_T_233[287:0] : _GEN_8172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9223 = 10'h127 == _T_23 ? _ram_T_233[287:0] : _GEN_8173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9224 = 10'h128 == _T_23 ? _ram_T_233[287:0] : _GEN_8174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9225 = 10'h129 == _T_23 ? _ram_T_233[287:0] : _GEN_8175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9226 = 10'h12a == _T_23 ? _ram_T_233[287:0] : _GEN_8176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9227 = 10'h12b == _T_23 ? _ram_T_233[287:0] : _GEN_8177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9228 = 10'h12c == _T_23 ? _ram_T_233[287:0] : _GEN_8178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9229 = 10'h12d == _T_23 ? _ram_T_233[287:0] : _GEN_8179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9230 = 10'h12e == _T_23 ? _ram_T_233[287:0] : _GEN_8180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9231 = 10'h12f == _T_23 ? _ram_T_233[287:0] : _GEN_8181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9232 = 10'h130 == _T_23 ? _ram_T_233[287:0] : _GEN_8182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9233 = 10'h131 == _T_23 ? _ram_T_233[287:0] : _GEN_8183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9234 = 10'h132 == _T_23 ? _ram_T_233[287:0] : _GEN_8184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9235 = 10'h133 == _T_23 ? _ram_T_233[287:0] : _GEN_8185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9236 = 10'h134 == _T_23 ? _ram_T_233[287:0] : _GEN_8186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9237 = 10'h135 == _T_23 ? _ram_T_233[287:0] : _GEN_8187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9238 = 10'h136 == _T_23 ? _ram_T_233[287:0] : _GEN_8188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9239 = 10'h137 == _T_23 ? _ram_T_233[287:0] : _GEN_8189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9240 = 10'h138 == _T_23 ? _ram_T_233[287:0] : _GEN_8190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9241 = 10'h139 == _T_23 ? _ram_T_233[287:0] : _GEN_8191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9242 = 10'h13a == _T_23 ? _ram_T_233[287:0] : _GEN_8192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9243 = 10'h13b == _T_23 ? _ram_T_233[287:0] : _GEN_8193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9244 = 10'h13c == _T_23 ? _ram_T_233[287:0] : _GEN_8194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9245 = 10'h13d == _T_23 ? _ram_T_233[287:0] : _GEN_8195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9246 = 10'h13e == _T_23 ? _ram_T_233[287:0] : _GEN_8196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9247 = 10'h13f == _T_23 ? _ram_T_233[287:0] : _GEN_8197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9248 = 10'h140 == _T_23 ? _ram_T_233[287:0] : _GEN_8198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9249 = 10'h141 == _T_23 ? _ram_T_233[287:0] : _GEN_8199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9250 = 10'h142 == _T_23 ? _ram_T_233[287:0] : _GEN_8200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9251 = 10'h143 == _T_23 ? _ram_T_233[287:0] : _GEN_8201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9252 = 10'h144 == _T_23 ? _ram_T_233[287:0] : _GEN_8202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9253 = 10'h145 == _T_23 ? _ram_T_233[287:0] : _GEN_8203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9254 = 10'h146 == _T_23 ? _ram_T_233[287:0] : _GEN_8204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9255 = 10'h147 == _T_23 ? _ram_T_233[287:0] : _GEN_8205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9256 = 10'h148 == _T_23 ? _ram_T_233[287:0] : _GEN_8206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9257 = 10'h149 == _T_23 ? _ram_T_233[287:0] : _GEN_8207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9258 = 10'h14a == _T_23 ? _ram_T_233[287:0] : _GEN_8208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9259 = 10'h14b == _T_23 ? _ram_T_233[287:0] : _GEN_8209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9260 = 10'h14c == _T_23 ? _ram_T_233[287:0] : _GEN_8210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9261 = 10'h14d == _T_23 ? _ram_T_233[287:0] : _GEN_8211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9262 = 10'h14e == _T_23 ? _ram_T_233[287:0] : _GEN_8212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9263 = 10'h14f == _T_23 ? _ram_T_233[287:0] : _GEN_8213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9264 = 10'h150 == _T_23 ? _ram_T_233[287:0] : _GEN_8214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9265 = 10'h151 == _T_23 ? _ram_T_233[287:0] : _GEN_8215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9266 = 10'h152 == _T_23 ? _ram_T_233[287:0] : _GEN_8216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9267 = 10'h153 == _T_23 ? _ram_T_233[287:0] : _GEN_8217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9268 = 10'h154 == _T_23 ? _ram_T_233[287:0] : _GEN_8218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9269 = 10'h155 == _T_23 ? _ram_T_233[287:0] : _GEN_8219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9270 = 10'h156 == _T_23 ? _ram_T_233[287:0] : _GEN_8220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9271 = 10'h157 == _T_23 ? _ram_T_233[287:0] : _GEN_8221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9272 = 10'h158 == _T_23 ? _ram_T_233[287:0] : _GEN_8222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9273 = 10'h159 == _T_23 ? _ram_T_233[287:0] : _GEN_8223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9274 = 10'h15a == _T_23 ? _ram_T_233[287:0] : _GEN_8224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9275 = 10'h15b == _T_23 ? _ram_T_233[287:0] : _GEN_8225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9276 = 10'h15c == _T_23 ? _ram_T_233[287:0] : _GEN_8226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9277 = 10'h15d == _T_23 ? _ram_T_233[287:0] : _GEN_8227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9278 = 10'h15e == _T_23 ? _ram_T_233[287:0] : _GEN_8228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9279 = 10'h15f == _T_23 ? _ram_T_233[287:0] : _GEN_8229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9280 = 10'h160 == _T_23 ? _ram_T_233[287:0] : _GEN_8230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9281 = 10'h161 == _T_23 ? _ram_T_233[287:0] : _GEN_8231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9282 = 10'h162 == _T_23 ? _ram_T_233[287:0] : _GEN_8232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9283 = 10'h163 == _T_23 ? _ram_T_233[287:0] : _GEN_8233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9284 = 10'h164 == _T_23 ? _ram_T_233[287:0] : _GEN_8234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9285 = 10'h165 == _T_23 ? _ram_T_233[287:0] : _GEN_8235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9286 = 10'h166 == _T_23 ? _ram_T_233[287:0] : _GEN_8236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9287 = 10'h167 == _T_23 ? _ram_T_233[287:0] : _GEN_8237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9288 = 10'h168 == _T_23 ? _ram_T_233[287:0] : _GEN_8238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9289 = 10'h169 == _T_23 ? _ram_T_233[287:0] : _GEN_8239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9290 = 10'h16a == _T_23 ? _ram_T_233[287:0] : _GEN_8240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9291 = 10'h16b == _T_23 ? _ram_T_233[287:0] : _GEN_8241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9292 = 10'h16c == _T_23 ? _ram_T_233[287:0] : _GEN_8242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9293 = 10'h16d == _T_23 ? _ram_T_233[287:0] : _GEN_8243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9294 = 10'h16e == _T_23 ? _ram_T_233[287:0] : _GEN_8244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9295 = 10'h16f == _T_23 ? _ram_T_233[287:0] : _GEN_8245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9296 = 10'h170 == _T_23 ? _ram_T_233[287:0] : _GEN_8246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9297 = 10'h171 == _T_23 ? _ram_T_233[287:0] : _GEN_8247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9298 = 10'h172 == _T_23 ? _ram_T_233[287:0] : _GEN_8248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9299 = 10'h173 == _T_23 ? _ram_T_233[287:0] : _GEN_8249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9300 = 10'h174 == _T_23 ? _ram_T_233[287:0] : _GEN_8250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9301 = 10'h175 == _T_23 ? _ram_T_233[287:0] : _GEN_8251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9302 = 10'h176 == _T_23 ? _ram_T_233[287:0] : _GEN_8252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9303 = 10'h177 == _T_23 ? _ram_T_233[287:0] : _GEN_8253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9304 = 10'h178 == _T_23 ? _ram_T_233[287:0] : _GEN_8254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9305 = 10'h179 == _T_23 ? _ram_T_233[287:0] : _GEN_8255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9306 = 10'h17a == _T_23 ? _ram_T_233[287:0] : _GEN_8256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9307 = 10'h17b == _T_23 ? _ram_T_233[287:0] : _GEN_8257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9308 = 10'h17c == _T_23 ? _ram_T_233[287:0] : _GEN_8258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9309 = 10'h17d == _T_23 ? _ram_T_233[287:0] : _GEN_8259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9310 = 10'h17e == _T_23 ? _ram_T_233[287:0] : _GEN_8260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9311 = 10'h17f == _T_23 ? _ram_T_233[287:0] : _GEN_8261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9312 = 10'h180 == _T_23 ? _ram_T_233[287:0] : _GEN_8262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9313 = 10'h181 == _T_23 ? _ram_T_233[287:0] : _GEN_8263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9314 = 10'h182 == _T_23 ? _ram_T_233[287:0] : _GEN_8264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9315 = 10'h183 == _T_23 ? _ram_T_233[287:0] : _GEN_8265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9316 = 10'h184 == _T_23 ? _ram_T_233[287:0] : _GEN_8266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9317 = 10'h185 == _T_23 ? _ram_T_233[287:0] : _GEN_8267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9318 = 10'h186 == _T_23 ? _ram_T_233[287:0] : _GEN_8268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9319 = 10'h187 == _T_23 ? _ram_T_233[287:0] : _GEN_8269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9320 = 10'h188 == _T_23 ? _ram_T_233[287:0] : _GEN_8270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9321 = 10'h189 == _T_23 ? _ram_T_233[287:0] : _GEN_8271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9322 = 10'h18a == _T_23 ? _ram_T_233[287:0] : _GEN_8272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9323 = 10'h18b == _T_23 ? _ram_T_233[287:0] : _GEN_8273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9324 = 10'h18c == _T_23 ? _ram_T_233[287:0] : _GEN_8274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9325 = 10'h18d == _T_23 ? _ram_T_233[287:0] : _GEN_8275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9326 = 10'h18e == _T_23 ? _ram_T_233[287:0] : _GEN_8276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9327 = 10'h18f == _T_23 ? _ram_T_233[287:0] : _GEN_8277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9328 = 10'h190 == _T_23 ? _ram_T_233[287:0] : _GEN_8278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9329 = 10'h191 == _T_23 ? _ram_T_233[287:0] : _GEN_8279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9330 = 10'h192 == _T_23 ? _ram_T_233[287:0] : _GEN_8280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9331 = 10'h193 == _T_23 ? _ram_T_233[287:0] : _GEN_8281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9332 = 10'h194 == _T_23 ? _ram_T_233[287:0] : _GEN_8282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9333 = 10'h195 == _T_23 ? _ram_T_233[287:0] : _GEN_8283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9334 = 10'h196 == _T_23 ? _ram_T_233[287:0] : _GEN_8284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9335 = 10'h197 == _T_23 ? _ram_T_233[287:0] : _GEN_8285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9336 = 10'h198 == _T_23 ? _ram_T_233[287:0] : _GEN_8286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9337 = 10'h199 == _T_23 ? _ram_T_233[287:0] : _GEN_8287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9338 = 10'h19a == _T_23 ? _ram_T_233[287:0] : _GEN_8288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9339 = 10'h19b == _T_23 ? _ram_T_233[287:0] : _GEN_8289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9340 = 10'h19c == _T_23 ? _ram_T_233[287:0] : _GEN_8290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9341 = 10'h19d == _T_23 ? _ram_T_233[287:0] : _GEN_8291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9342 = 10'h19e == _T_23 ? _ram_T_233[287:0] : _GEN_8292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9343 = 10'h19f == _T_23 ? _ram_T_233[287:0] : _GEN_8293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9344 = 10'h1a0 == _T_23 ? _ram_T_233[287:0] : _GEN_8294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9345 = 10'h1a1 == _T_23 ? _ram_T_233[287:0] : _GEN_8295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9346 = 10'h1a2 == _T_23 ? _ram_T_233[287:0] : _GEN_8296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9347 = 10'h1a3 == _T_23 ? _ram_T_233[287:0] : _GEN_8297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9348 = 10'h1a4 == _T_23 ? _ram_T_233[287:0] : _GEN_8298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9349 = 10'h1a5 == _T_23 ? _ram_T_233[287:0] : _GEN_8299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9350 = 10'h1a6 == _T_23 ? _ram_T_233[287:0] : _GEN_8300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9351 = 10'h1a7 == _T_23 ? _ram_T_233[287:0] : _GEN_8301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9352 = 10'h1a8 == _T_23 ? _ram_T_233[287:0] : _GEN_8302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9353 = 10'h1a9 == _T_23 ? _ram_T_233[287:0] : _GEN_8303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9354 = 10'h1aa == _T_23 ? _ram_T_233[287:0] : _GEN_8304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9355 = 10'h1ab == _T_23 ? _ram_T_233[287:0] : _GEN_8305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9356 = 10'h1ac == _T_23 ? _ram_T_233[287:0] : _GEN_8306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9357 = 10'h1ad == _T_23 ? _ram_T_233[287:0] : _GEN_8307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9358 = 10'h1ae == _T_23 ? _ram_T_233[287:0] : _GEN_8308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9359 = 10'h1af == _T_23 ? _ram_T_233[287:0] : _GEN_8309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9360 = 10'h1b0 == _T_23 ? _ram_T_233[287:0] : _GEN_8310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9361 = 10'h1b1 == _T_23 ? _ram_T_233[287:0] : _GEN_8311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9362 = 10'h1b2 == _T_23 ? _ram_T_233[287:0] : _GEN_8312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9363 = 10'h1b3 == _T_23 ? _ram_T_233[287:0] : _GEN_8313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9364 = 10'h1b4 == _T_23 ? _ram_T_233[287:0] : _GEN_8314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9365 = 10'h1b5 == _T_23 ? _ram_T_233[287:0] : _GEN_8315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9366 = 10'h1b6 == _T_23 ? _ram_T_233[287:0] : _GEN_8316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9367 = 10'h1b7 == _T_23 ? _ram_T_233[287:0] : _GEN_8317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9368 = 10'h1b8 == _T_23 ? _ram_T_233[287:0] : _GEN_8318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9369 = 10'h1b9 == _T_23 ? _ram_T_233[287:0] : _GEN_8319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9370 = 10'h1ba == _T_23 ? _ram_T_233[287:0] : _GEN_8320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9371 = 10'h1bb == _T_23 ? _ram_T_233[287:0] : _GEN_8321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9372 = 10'h1bc == _T_23 ? _ram_T_233[287:0] : _GEN_8322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9373 = 10'h1bd == _T_23 ? _ram_T_233[287:0] : _GEN_8323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9374 = 10'h1be == _T_23 ? _ram_T_233[287:0] : _GEN_8324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9375 = 10'h1bf == _T_23 ? _ram_T_233[287:0] : _GEN_8325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9376 = 10'h1c0 == _T_23 ? _ram_T_233[287:0] : _GEN_8326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9377 = 10'h1c1 == _T_23 ? _ram_T_233[287:0] : _GEN_8327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9378 = 10'h1c2 == _T_23 ? _ram_T_233[287:0] : _GEN_8328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9379 = 10'h1c3 == _T_23 ? _ram_T_233[287:0] : _GEN_8329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9380 = 10'h1c4 == _T_23 ? _ram_T_233[287:0] : _GEN_8330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9381 = 10'h1c5 == _T_23 ? _ram_T_233[287:0] : _GEN_8331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9382 = 10'h1c6 == _T_23 ? _ram_T_233[287:0] : _GEN_8332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9383 = 10'h1c7 == _T_23 ? _ram_T_233[287:0] : _GEN_8333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9384 = 10'h1c8 == _T_23 ? _ram_T_233[287:0] : _GEN_8334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9385 = 10'h1c9 == _T_23 ? _ram_T_233[287:0] : _GEN_8335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9386 = 10'h1ca == _T_23 ? _ram_T_233[287:0] : _GEN_8336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9387 = 10'h1cb == _T_23 ? _ram_T_233[287:0] : _GEN_8337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9388 = 10'h1cc == _T_23 ? _ram_T_233[287:0] : _GEN_8338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9389 = 10'h1cd == _T_23 ? _ram_T_233[287:0] : _GEN_8339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9390 = 10'h1ce == _T_23 ? _ram_T_233[287:0] : _GEN_8340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9391 = 10'h1cf == _T_23 ? _ram_T_233[287:0] : _GEN_8341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9392 = 10'h1d0 == _T_23 ? _ram_T_233[287:0] : _GEN_8342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9393 = 10'h1d1 == _T_23 ? _ram_T_233[287:0] : _GEN_8343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9394 = 10'h1d2 == _T_23 ? _ram_T_233[287:0] : _GEN_8344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9395 = 10'h1d3 == _T_23 ? _ram_T_233[287:0] : _GEN_8345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9396 = 10'h1d4 == _T_23 ? _ram_T_233[287:0] : _GEN_8346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9397 = 10'h1d5 == _T_23 ? _ram_T_233[287:0] : _GEN_8347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9398 = 10'h1d6 == _T_23 ? _ram_T_233[287:0] : _GEN_8348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9399 = 10'h1d7 == _T_23 ? _ram_T_233[287:0] : _GEN_8349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9400 = 10'h1d8 == _T_23 ? _ram_T_233[287:0] : _GEN_8350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9401 = 10'h1d9 == _T_23 ? _ram_T_233[287:0] : _GEN_8351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9402 = 10'h1da == _T_23 ? _ram_T_233[287:0] : _GEN_8352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9403 = 10'h1db == _T_23 ? _ram_T_233[287:0] : _GEN_8353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9404 = 10'h1dc == _T_23 ? _ram_T_233[287:0] : _GEN_8354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9405 = 10'h1dd == _T_23 ? _ram_T_233[287:0] : _GEN_8355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9406 = 10'h1de == _T_23 ? _ram_T_233[287:0] : _GEN_8356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9407 = 10'h1df == _T_23 ? _ram_T_233[287:0] : _GEN_8357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9408 = 10'h1e0 == _T_23 ? _ram_T_233[287:0] : _GEN_8358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9409 = 10'h1e1 == _T_23 ? _ram_T_233[287:0] : _GEN_8359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9410 = 10'h1e2 == _T_23 ? _ram_T_233[287:0] : _GEN_8360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9411 = 10'h1e3 == _T_23 ? _ram_T_233[287:0] : _GEN_8361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9412 = 10'h1e4 == _T_23 ? _ram_T_233[287:0] : _GEN_8362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9413 = 10'h1e5 == _T_23 ? _ram_T_233[287:0] : _GEN_8363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9414 = 10'h1e6 == _T_23 ? _ram_T_233[287:0] : _GEN_8364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9415 = 10'h1e7 == _T_23 ? _ram_T_233[287:0] : _GEN_8365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9416 = 10'h1e8 == _T_23 ? _ram_T_233[287:0] : _GEN_8366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9417 = 10'h1e9 == _T_23 ? _ram_T_233[287:0] : _GEN_8367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9418 = 10'h1ea == _T_23 ? _ram_T_233[287:0] : _GEN_8368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9419 = 10'h1eb == _T_23 ? _ram_T_233[287:0] : _GEN_8369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9420 = 10'h1ec == _T_23 ? _ram_T_233[287:0] : _GEN_8370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9421 = 10'h1ed == _T_23 ? _ram_T_233[287:0] : _GEN_8371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9422 = 10'h1ee == _T_23 ? _ram_T_233[287:0] : _GEN_8372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9423 = 10'h1ef == _T_23 ? _ram_T_233[287:0] : _GEN_8373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9424 = 10'h1f0 == _T_23 ? _ram_T_233[287:0] : _GEN_8374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9425 = 10'h1f1 == _T_23 ? _ram_T_233[287:0] : _GEN_8375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9426 = 10'h1f2 == _T_23 ? _ram_T_233[287:0] : _GEN_8376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9427 = 10'h1f3 == _T_23 ? _ram_T_233[287:0] : _GEN_8377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9428 = 10'h1f4 == _T_23 ? _ram_T_233[287:0] : _GEN_8378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9429 = 10'h1f5 == _T_23 ? _ram_T_233[287:0] : _GEN_8379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9430 = 10'h1f6 == _T_23 ? _ram_T_233[287:0] : _GEN_8380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9431 = 10'h1f7 == _T_23 ? _ram_T_233[287:0] : _GEN_8381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9432 = 10'h1f8 == _T_23 ? _ram_T_233[287:0] : _GEN_8382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9433 = 10'h1f9 == _T_23 ? _ram_T_233[287:0] : _GEN_8383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9434 = 10'h1fa == _T_23 ? _ram_T_233[287:0] : _GEN_8384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9435 = 10'h1fb == _T_23 ? _ram_T_233[287:0] : _GEN_8385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9436 = 10'h1fc == _T_23 ? _ram_T_233[287:0] : _GEN_8386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9437 = 10'h1fd == _T_23 ? _ram_T_233[287:0] : _GEN_8387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9438 = 10'h1fe == _T_23 ? _ram_T_233[287:0] : _GEN_8388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9439 = 10'h1ff == _T_23 ? _ram_T_233[287:0] : _GEN_8389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9440 = 10'h200 == _T_23 ? _ram_T_233[287:0] : _GEN_8390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9441 = 10'h201 == _T_23 ? _ram_T_233[287:0] : _GEN_8391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9442 = 10'h202 == _T_23 ? _ram_T_233[287:0] : _GEN_8392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9443 = 10'h203 == _T_23 ? _ram_T_233[287:0] : _GEN_8393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9444 = 10'h204 == _T_23 ? _ram_T_233[287:0] : _GEN_8394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9445 = 10'h205 == _T_23 ? _ram_T_233[287:0] : _GEN_8395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9446 = 10'h206 == _T_23 ? _ram_T_233[287:0] : _GEN_8396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9447 = 10'h207 == _T_23 ? _ram_T_233[287:0] : _GEN_8397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9448 = 10'h208 == _T_23 ? _ram_T_233[287:0] : _GEN_8398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9449 = 10'h209 == _T_23 ? _ram_T_233[287:0] : _GEN_8399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9450 = 10'h20a == _T_23 ? _ram_T_233[287:0] : _GEN_8400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9451 = 10'h20b == _T_23 ? _ram_T_233[287:0] : _GEN_8401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9452 = 10'h20c == _T_23 ? _ram_T_233[287:0] : _GEN_8402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_25 = h + 10'h9; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_9 = vga_mem_ram_MPORT_81_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_9 = vga_mem_ram_MPORT_82_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_9 = vga_mem_ram_MPORT_83_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_9 = vga_mem_ram_MPORT_84_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_9 = vga_mem_ram_MPORT_85_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_9 = vga_mem_ram_MPORT_86_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_9 = vga_mem_ram_MPORT_87_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_9 = vga_mem_ram_MPORT_88_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_9 = vga_mem_ram_MPORT_89_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_254 = {278'h0,ram_hi_hi_hi_lo_9,ram_hi_hi_lo_9,ram_hi_lo_hi_9,ram_hi_lo_lo_9,ram_lo_hi_hi_hi_9,
    ram_lo_hi_hi_lo_9,ram_lo_hi_lo_9,ram_lo_lo_hi_9,ram_lo_lo_lo_9}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19078 = {{8191'd0}, _ram_T_254}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_258 = _GEN_19078 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_9454 = 10'h1 == _T_25 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9455 = 10'h2 == _T_25 ? ram_2 : _GEN_9454; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9456 = 10'h3 == _T_25 ? ram_3 : _GEN_9455; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9457 = 10'h4 == _T_25 ? ram_4 : _GEN_9456; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9458 = 10'h5 == _T_25 ? ram_5 : _GEN_9457; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9459 = 10'h6 == _T_25 ? ram_6 : _GEN_9458; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9460 = 10'h7 == _T_25 ? ram_7 : _GEN_9459; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9461 = 10'h8 == _T_25 ? ram_8 : _GEN_9460; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9462 = 10'h9 == _T_25 ? ram_9 : _GEN_9461; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9463 = 10'ha == _T_25 ? ram_10 : _GEN_9462; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9464 = 10'hb == _T_25 ? ram_11 : _GEN_9463; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9465 = 10'hc == _T_25 ? ram_12 : _GEN_9464; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9466 = 10'hd == _T_25 ? ram_13 : _GEN_9465; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9467 = 10'he == _T_25 ? ram_14 : _GEN_9466; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9468 = 10'hf == _T_25 ? ram_15 : _GEN_9467; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9469 = 10'h10 == _T_25 ? ram_16 : _GEN_9468; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9470 = 10'h11 == _T_25 ? ram_17 : _GEN_9469; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9471 = 10'h12 == _T_25 ? ram_18 : _GEN_9470; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9472 = 10'h13 == _T_25 ? ram_19 : _GEN_9471; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9473 = 10'h14 == _T_25 ? ram_20 : _GEN_9472; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9474 = 10'h15 == _T_25 ? ram_21 : _GEN_9473; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9475 = 10'h16 == _T_25 ? ram_22 : _GEN_9474; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9476 = 10'h17 == _T_25 ? ram_23 : _GEN_9475; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9477 = 10'h18 == _T_25 ? ram_24 : _GEN_9476; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9478 = 10'h19 == _T_25 ? ram_25 : _GEN_9477; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9479 = 10'h1a == _T_25 ? ram_26 : _GEN_9478; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9480 = 10'h1b == _T_25 ? ram_27 : _GEN_9479; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9481 = 10'h1c == _T_25 ? ram_28 : _GEN_9480; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9482 = 10'h1d == _T_25 ? ram_29 : _GEN_9481; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9483 = 10'h1e == _T_25 ? ram_30 : _GEN_9482; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9484 = 10'h1f == _T_25 ? ram_31 : _GEN_9483; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9485 = 10'h20 == _T_25 ? ram_32 : _GEN_9484; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9486 = 10'h21 == _T_25 ? ram_33 : _GEN_9485; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9487 = 10'h22 == _T_25 ? ram_34 : _GEN_9486; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9488 = 10'h23 == _T_25 ? ram_35 : _GEN_9487; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9489 = 10'h24 == _T_25 ? ram_36 : _GEN_9488; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9490 = 10'h25 == _T_25 ? ram_37 : _GEN_9489; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9491 = 10'h26 == _T_25 ? ram_38 : _GEN_9490; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9492 = 10'h27 == _T_25 ? ram_39 : _GEN_9491; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9493 = 10'h28 == _T_25 ? ram_40 : _GEN_9492; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9494 = 10'h29 == _T_25 ? ram_41 : _GEN_9493; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9495 = 10'h2a == _T_25 ? ram_42 : _GEN_9494; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9496 = 10'h2b == _T_25 ? ram_43 : _GEN_9495; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9497 = 10'h2c == _T_25 ? ram_44 : _GEN_9496; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9498 = 10'h2d == _T_25 ? ram_45 : _GEN_9497; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9499 = 10'h2e == _T_25 ? ram_46 : _GEN_9498; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9500 = 10'h2f == _T_25 ? ram_47 : _GEN_9499; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9501 = 10'h30 == _T_25 ? ram_48 : _GEN_9500; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9502 = 10'h31 == _T_25 ? ram_49 : _GEN_9501; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9503 = 10'h32 == _T_25 ? ram_50 : _GEN_9502; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9504 = 10'h33 == _T_25 ? ram_51 : _GEN_9503; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9505 = 10'h34 == _T_25 ? ram_52 : _GEN_9504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9506 = 10'h35 == _T_25 ? ram_53 : _GEN_9505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9507 = 10'h36 == _T_25 ? ram_54 : _GEN_9506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9508 = 10'h37 == _T_25 ? ram_55 : _GEN_9507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9509 = 10'h38 == _T_25 ? ram_56 : _GEN_9508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9510 = 10'h39 == _T_25 ? ram_57 : _GEN_9509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9511 = 10'h3a == _T_25 ? ram_58 : _GEN_9510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9512 = 10'h3b == _T_25 ? ram_59 : _GEN_9511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9513 = 10'h3c == _T_25 ? ram_60 : _GEN_9512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9514 = 10'h3d == _T_25 ? ram_61 : _GEN_9513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9515 = 10'h3e == _T_25 ? ram_62 : _GEN_9514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9516 = 10'h3f == _T_25 ? ram_63 : _GEN_9515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9517 = 10'h40 == _T_25 ? ram_64 : _GEN_9516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9518 = 10'h41 == _T_25 ? ram_65 : _GEN_9517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9519 = 10'h42 == _T_25 ? ram_66 : _GEN_9518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9520 = 10'h43 == _T_25 ? ram_67 : _GEN_9519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9521 = 10'h44 == _T_25 ? ram_68 : _GEN_9520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9522 = 10'h45 == _T_25 ? ram_69 : _GEN_9521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9523 = 10'h46 == _T_25 ? ram_70 : _GEN_9522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9524 = 10'h47 == _T_25 ? ram_71 : _GEN_9523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9525 = 10'h48 == _T_25 ? ram_72 : _GEN_9524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9526 = 10'h49 == _T_25 ? ram_73 : _GEN_9525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9527 = 10'h4a == _T_25 ? ram_74 : _GEN_9526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9528 = 10'h4b == _T_25 ? ram_75 : _GEN_9527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9529 = 10'h4c == _T_25 ? ram_76 : _GEN_9528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9530 = 10'h4d == _T_25 ? ram_77 : _GEN_9529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9531 = 10'h4e == _T_25 ? ram_78 : _GEN_9530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9532 = 10'h4f == _T_25 ? ram_79 : _GEN_9531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9533 = 10'h50 == _T_25 ? ram_80 : _GEN_9532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9534 = 10'h51 == _T_25 ? ram_81 : _GEN_9533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9535 = 10'h52 == _T_25 ? ram_82 : _GEN_9534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9536 = 10'h53 == _T_25 ? ram_83 : _GEN_9535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9537 = 10'h54 == _T_25 ? ram_84 : _GEN_9536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9538 = 10'h55 == _T_25 ? ram_85 : _GEN_9537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9539 = 10'h56 == _T_25 ? ram_86 : _GEN_9538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9540 = 10'h57 == _T_25 ? ram_87 : _GEN_9539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9541 = 10'h58 == _T_25 ? ram_88 : _GEN_9540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9542 = 10'h59 == _T_25 ? ram_89 : _GEN_9541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9543 = 10'h5a == _T_25 ? ram_90 : _GEN_9542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9544 = 10'h5b == _T_25 ? ram_91 : _GEN_9543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9545 = 10'h5c == _T_25 ? ram_92 : _GEN_9544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9546 = 10'h5d == _T_25 ? ram_93 : _GEN_9545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9547 = 10'h5e == _T_25 ? ram_94 : _GEN_9546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9548 = 10'h5f == _T_25 ? ram_95 : _GEN_9547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9549 = 10'h60 == _T_25 ? ram_96 : _GEN_9548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9550 = 10'h61 == _T_25 ? ram_97 : _GEN_9549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9551 = 10'h62 == _T_25 ? ram_98 : _GEN_9550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9552 = 10'h63 == _T_25 ? ram_99 : _GEN_9551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9553 = 10'h64 == _T_25 ? ram_100 : _GEN_9552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9554 = 10'h65 == _T_25 ? ram_101 : _GEN_9553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9555 = 10'h66 == _T_25 ? ram_102 : _GEN_9554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9556 = 10'h67 == _T_25 ? ram_103 : _GEN_9555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9557 = 10'h68 == _T_25 ? ram_104 : _GEN_9556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9558 = 10'h69 == _T_25 ? ram_105 : _GEN_9557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9559 = 10'h6a == _T_25 ? ram_106 : _GEN_9558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9560 = 10'h6b == _T_25 ? ram_107 : _GEN_9559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9561 = 10'h6c == _T_25 ? ram_108 : _GEN_9560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9562 = 10'h6d == _T_25 ? ram_109 : _GEN_9561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9563 = 10'h6e == _T_25 ? ram_110 : _GEN_9562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9564 = 10'h6f == _T_25 ? ram_111 : _GEN_9563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9565 = 10'h70 == _T_25 ? ram_112 : _GEN_9564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9566 = 10'h71 == _T_25 ? ram_113 : _GEN_9565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9567 = 10'h72 == _T_25 ? ram_114 : _GEN_9566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9568 = 10'h73 == _T_25 ? ram_115 : _GEN_9567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9569 = 10'h74 == _T_25 ? ram_116 : _GEN_9568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9570 = 10'h75 == _T_25 ? ram_117 : _GEN_9569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9571 = 10'h76 == _T_25 ? ram_118 : _GEN_9570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9572 = 10'h77 == _T_25 ? ram_119 : _GEN_9571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9573 = 10'h78 == _T_25 ? ram_120 : _GEN_9572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9574 = 10'h79 == _T_25 ? ram_121 : _GEN_9573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9575 = 10'h7a == _T_25 ? ram_122 : _GEN_9574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9576 = 10'h7b == _T_25 ? ram_123 : _GEN_9575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9577 = 10'h7c == _T_25 ? ram_124 : _GEN_9576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9578 = 10'h7d == _T_25 ? ram_125 : _GEN_9577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9579 = 10'h7e == _T_25 ? ram_126 : _GEN_9578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9580 = 10'h7f == _T_25 ? ram_127 : _GEN_9579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9581 = 10'h80 == _T_25 ? ram_128 : _GEN_9580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9582 = 10'h81 == _T_25 ? ram_129 : _GEN_9581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9583 = 10'h82 == _T_25 ? ram_130 : _GEN_9582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9584 = 10'h83 == _T_25 ? ram_131 : _GEN_9583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9585 = 10'h84 == _T_25 ? ram_132 : _GEN_9584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9586 = 10'h85 == _T_25 ? ram_133 : _GEN_9585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9587 = 10'h86 == _T_25 ? ram_134 : _GEN_9586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9588 = 10'h87 == _T_25 ? ram_135 : _GEN_9587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9589 = 10'h88 == _T_25 ? ram_136 : _GEN_9588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9590 = 10'h89 == _T_25 ? ram_137 : _GEN_9589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9591 = 10'h8a == _T_25 ? ram_138 : _GEN_9590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9592 = 10'h8b == _T_25 ? ram_139 : _GEN_9591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9593 = 10'h8c == _T_25 ? ram_140 : _GEN_9592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9594 = 10'h8d == _T_25 ? ram_141 : _GEN_9593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9595 = 10'h8e == _T_25 ? ram_142 : _GEN_9594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9596 = 10'h8f == _T_25 ? ram_143 : _GEN_9595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9597 = 10'h90 == _T_25 ? ram_144 : _GEN_9596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9598 = 10'h91 == _T_25 ? ram_145 : _GEN_9597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9599 = 10'h92 == _T_25 ? ram_146 : _GEN_9598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9600 = 10'h93 == _T_25 ? ram_147 : _GEN_9599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9601 = 10'h94 == _T_25 ? ram_148 : _GEN_9600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9602 = 10'h95 == _T_25 ? ram_149 : _GEN_9601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9603 = 10'h96 == _T_25 ? ram_150 : _GEN_9602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9604 = 10'h97 == _T_25 ? ram_151 : _GEN_9603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9605 = 10'h98 == _T_25 ? ram_152 : _GEN_9604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9606 = 10'h99 == _T_25 ? ram_153 : _GEN_9605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9607 = 10'h9a == _T_25 ? ram_154 : _GEN_9606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9608 = 10'h9b == _T_25 ? ram_155 : _GEN_9607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9609 = 10'h9c == _T_25 ? ram_156 : _GEN_9608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9610 = 10'h9d == _T_25 ? ram_157 : _GEN_9609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9611 = 10'h9e == _T_25 ? ram_158 : _GEN_9610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9612 = 10'h9f == _T_25 ? ram_159 : _GEN_9611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9613 = 10'ha0 == _T_25 ? ram_160 : _GEN_9612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9614 = 10'ha1 == _T_25 ? ram_161 : _GEN_9613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9615 = 10'ha2 == _T_25 ? ram_162 : _GEN_9614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9616 = 10'ha3 == _T_25 ? ram_163 : _GEN_9615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9617 = 10'ha4 == _T_25 ? ram_164 : _GEN_9616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9618 = 10'ha5 == _T_25 ? ram_165 : _GEN_9617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9619 = 10'ha6 == _T_25 ? ram_166 : _GEN_9618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9620 = 10'ha7 == _T_25 ? ram_167 : _GEN_9619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9621 = 10'ha8 == _T_25 ? ram_168 : _GEN_9620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9622 = 10'ha9 == _T_25 ? ram_169 : _GEN_9621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9623 = 10'haa == _T_25 ? ram_170 : _GEN_9622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9624 = 10'hab == _T_25 ? ram_171 : _GEN_9623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9625 = 10'hac == _T_25 ? ram_172 : _GEN_9624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9626 = 10'had == _T_25 ? ram_173 : _GEN_9625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9627 = 10'hae == _T_25 ? ram_174 : _GEN_9626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9628 = 10'haf == _T_25 ? ram_175 : _GEN_9627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9629 = 10'hb0 == _T_25 ? ram_176 : _GEN_9628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9630 = 10'hb1 == _T_25 ? ram_177 : _GEN_9629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9631 = 10'hb2 == _T_25 ? ram_178 : _GEN_9630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9632 = 10'hb3 == _T_25 ? ram_179 : _GEN_9631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9633 = 10'hb4 == _T_25 ? ram_180 : _GEN_9632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9634 = 10'hb5 == _T_25 ? ram_181 : _GEN_9633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9635 = 10'hb6 == _T_25 ? ram_182 : _GEN_9634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9636 = 10'hb7 == _T_25 ? ram_183 : _GEN_9635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9637 = 10'hb8 == _T_25 ? ram_184 : _GEN_9636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9638 = 10'hb9 == _T_25 ? ram_185 : _GEN_9637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9639 = 10'hba == _T_25 ? ram_186 : _GEN_9638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9640 = 10'hbb == _T_25 ? ram_187 : _GEN_9639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9641 = 10'hbc == _T_25 ? ram_188 : _GEN_9640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9642 = 10'hbd == _T_25 ? ram_189 : _GEN_9641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9643 = 10'hbe == _T_25 ? ram_190 : _GEN_9642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9644 = 10'hbf == _T_25 ? ram_191 : _GEN_9643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9645 = 10'hc0 == _T_25 ? ram_192 : _GEN_9644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9646 = 10'hc1 == _T_25 ? ram_193 : _GEN_9645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9647 = 10'hc2 == _T_25 ? ram_194 : _GEN_9646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9648 = 10'hc3 == _T_25 ? ram_195 : _GEN_9647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9649 = 10'hc4 == _T_25 ? ram_196 : _GEN_9648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9650 = 10'hc5 == _T_25 ? ram_197 : _GEN_9649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9651 = 10'hc6 == _T_25 ? ram_198 : _GEN_9650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9652 = 10'hc7 == _T_25 ? ram_199 : _GEN_9651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9653 = 10'hc8 == _T_25 ? ram_200 : _GEN_9652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9654 = 10'hc9 == _T_25 ? ram_201 : _GEN_9653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9655 = 10'hca == _T_25 ? ram_202 : _GEN_9654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9656 = 10'hcb == _T_25 ? ram_203 : _GEN_9655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9657 = 10'hcc == _T_25 ? ram_204 : _GEN_9656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9658 = 10'hcd == _T_25 ? ram_205 : _GEN_9657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9659 = 10'hce == _T_25 ? ram_206 : _GEN_9658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9660 = 10'hcf == _T_25 ? ram_207 : _GEN_9659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9661 = 10'hd0 == _T_25 ? ram_208 : _GEN_9660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9662 = 10'hd1 == _T_25 ? ram_209 : _GEN_9661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9663 = 10'hd2 == _T_25 ? ram_210 : _GEN_9662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9664 = 10'hd3 == _T_25 ? ram_211 : _GEN_9663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9665 = 10'hd4 == _T_25 ? ram_212 : _GEN_9664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9666 = 10'hd5 == _T_25 ? ram_213 : _GEN_9665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9667 = 10'hd6 == _T_25 ? ram_214 : _GEN_9666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9668 = 10'hd7 == _T_25 ? ram_215 : _GEN_9667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9669 = 10'hd8 == _T_25 ? ram_216 : _GEN_9668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9670 = 10'hd9 == _T_25 ? ram_217 : _GEN_9669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9671 = 10'hda == _T_25 ? ram_218 : _GEN_9670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9672 = 10'hdb == _T_25 ? ram_219 : _GEN_9671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9673 = 10'hdc == _T_25 ? ram_220 : _GEN_9672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9674 = 10'hdd == _T_25 ? ram_221 : _GEN_9673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9675 = 10'hde == _T_25 ? ram_222 : _GEN_9674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9676 = 10'hdf == _T_25 ? ram_223 : _GEN_9675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9677 = 10'he0 == _T_25 ? ram_224 : _GEN_9676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9678 = 10'he1 == _T_25 ? ram_225 : _GEN_9677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9679 = 10'he2 == _T_25 ? ram_226 : _GEN_9678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9680 = 10'he3 == _T_25 ? ram_227 : _GEN_9679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9681 = 10'he4 == _T_25 ? ram_228 : _GEN_9680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9682 = 10'he5 == _T_25 ? ram_229 : _GEN_9681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9683 = 10'he6 == _T_25 ? ram_230 : _GEN_9682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9684 = 10'he7 == _T_25 ? ram_231 : _GEN_9683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9685 = 10'he8 == _T_25 ? ram_232 : _GEN_9684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9686 = 10'he9 == _T_25 ? ram_233 : _GEN_9685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9687 = 10'hea == _T_25 ? ram_234 : _GEN_9686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9688 = 10'heb == _T_25 ? ram_235 : _GEN_9687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9689 = 10'hec == _T_25 ? ram_236 : _GEN_9688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9690 = 10'hed == _T_25 ? ram_237 : _GEN_9689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9691 = 10'hee == _T_25 ? ram_238 : _GEN_9690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9692 = 10'hef == _T_25 ? ram_239 : _GEN_9691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9693 = 10'hf0 == _T_25 ? ram_240 : _GEN_9692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9694 = 10'hf1 == _T_25 ? ram_241 : _GEN_9693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9695 = 10'hf2 == _T_25 ? ram_242 : _GEN_9694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9696 = 10'hf3 == _T_25 ? ram_243 : _GEN_9695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9697 = 10'hf4 == _T_25 ? ram_244 : _GEN_9696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9698 = 10'hf5 == _T_25 ? ram_245 : _GEN_9697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9699 = 10'hf6 == _T_25 ? ram_246 : _GEN_9698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9700 = 10'hf7 == _T_25 ? ram_247 : _GEN_9699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9701 = 10'hf8 == _T_25 ? ram_248 : _GEN_9700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9702 = 10'hf9 == _T_25 ? ram_249 : _GEN_9701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9703 = 10'hfa == _T_25 ? ram_250 : _GEN_9702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9704 = 10'hfb == _T_25 ? ram_251 : _GEN_9703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9705 = 10'hfc == _T_25 ? ram_252 : _GEN_9704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9706 = 10'hfd == _T_25 ? ram_253 : _GEN_9705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9707 = 10'hfe == _T_25 ? ram_254 : _GEN_9706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9708 = 10'hff == _T_25 ? ram_255 : _GEN_9707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9709 = 10'h100 == _T_25 ? ram_256 : _GEN_9708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9710 = 10'h101 == _T_25 ? ram_257 : _GEN_9709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9711 = 10'h102 == _T_25 ? ram_258 : _GEN_9710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9712 = 10'h103 == _T_25 ? ram_259 : _GEN_9711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9713 = 10'h104 == _T_25 ? ram_260 : _GEN_9712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9714 = 10'h105 == _T_25 ? ram_261 : _GEN_9713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9715 = 10'h106 == _T_25 ? ram_262 : _GEN_9714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9716 = 10'h107 == _T_25 ? ram_263 : _GEN_9715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9717 = 10'h108 == _T_25 ? ram_264 : _GEN_9716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9718 = 10'h109 == _T_25 ? ram_265 : _GEN_9717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9719 = 10'h10a == _T_25 ? ram_266 : _GEN_9718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9720 = 10'h10b == _T_25 ? ram_267 : _GEN_9719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9721 = 10'h10c == _T_25 ? ram_268 : _GEN_9720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9722 = 10'h10d == _T_25 ? ram_269 : _GEN_9721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9723 = 10'h10e == _T_25 ? ram_270 : _GEN_9722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9724 = 10'h10f == _T_25 ? ram_271 : _GEN_9723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9725 = 10'h110 == _T_25 ? ram_272 : _GEN_9724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9726 = 10'h111 == _T_25 ? ram_273 : _GEN_9725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9727 = 10'h112 == _T_25 ? ram_274 : _GEN_9726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9728 = 10'h113 == _T_25 ? ram_275 : _GEN_9727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9729 = 10'h114 == _T_25 ? ram_276 : _GEN_9728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9730 = 10'h115 == _T_25 ? ram_277 : _GEN_9729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9731 = 10'h116 == _T_25 ? ram_278 : _GEN_9730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9732 = 10'h117 == _T_25 ? ram_279 : _GEN_9731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9733 = 10'h118 == _T_25 ? ram_280 : _GEN_9732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9734 = 10'h119 == _T_25 ? ram_281 : _GEN_9733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9735 = 10'h11a == _T_25 ? ram_282 : _GEN_9734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9736 = 10'h11b == _T_25 ? ram_283 : _GEN_9735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9737 = 10'h11c == _T_25 ? ram_284 : _GEN_9736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9738 = 10'h11d == _T_25 ? ram_285 : _GEN_9737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9739 = 10'h11e == _T_25 ? ram_286 : _GEN_9738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9740 = 10'h11f == _T_25 ? ram_287 : _GEN_9739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9741 = 10'h120 == _T_25 ? ram_288 : _GEN_9740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9742 = 10'h121 == _T_25 ? ram_289 : _GEN_9741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9743 = 10'h122 == _T_25 ? ram_290 : _GEN_9742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9744 = 10'h123 == _T_25 ? ram_291 : _GEN_9743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9745 = 10'h124 == _T_25 ? ram_292 : _GEN_9744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9746 = 10'h125 == _T_25 ? ram_293 : _GEN_9745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9747 = 10'h126 == _T_25 ? ram_294 : _GEN_9746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9748 = 10'h127 == _T_25 ? ram_295 : _GEN_9747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9749 = 10'h128 == _T_25 ? ram_296 : _GEN_9748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9750 = 10'h129 == _T_25 ? ram_297 : _GEN_9749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9751 = 10'h12a == _T_25 ? ram_298 : _GEN_9750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9752 = 10'h12b == _T_25 ? ram_299 : _GEN_9751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9753 = 10'h12c == _T_25 ? ram_300 : _GEN_9752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9754 = 10'h12d == _T_25 ? ram_301 : _GEN_9753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9755 = 10'h12e == _T_25 ? ram_302 : _GEN_9754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9756 = 10'h12f == _T_25 ? ram_303 : _GEN_9755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9757 = 10'h130 == _T_25 ? ram_304 : _GEN_9756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9758 = 10'h131 == _T_25 ? ram_305 : _GEN_9757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9759 = 10'h132 == _T_25 ? ram_306 : _GEN_9758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9760 = 10'h133 == _T_25 ? ram_307 : _GEN_9759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9761 = 10'h134 == _T_25 ? ram_308 : _GEN_9760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9762 = 10'h135 == _T_25 ? ram_309 : _GEN_9761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9763 = 10'h136 == _T_25 ? ram_310 : _GEN_9762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9764 = 10'h137 == _T_25 ? ram_311 : _GEN_9763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9765 = 10'h138 == _T_25 ? ram_312 : _GEN_9764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9766 = 10'h139 == _T_25 ? ram_313 : _GEN_9765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9767 = 10'h13a == _T_25 ? ram_314 : _GEN_9766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9768 = 10'h13b == _T_25 ? ram_315 : _GEN_9767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9769 = 10'h13c == _T_25 ? ram_316 : _GEN_9768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9770 = 10'h13d == _T_25 ? ram_317 : _GEN_9769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9771 = 10'h13e == _T_25 ? ram_318 : _GEN_9770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9772 = 10'h13f == _T_25 ? ram_319 : _GEN_9771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9773 = 10'h140 == _T_25 ? ram_320 : _GEN_9772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9774 = 10'h141 == _T_25 ? ram_321 : _GEN_9773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9775 = 10'h142 == _T_25 ? ram_322 : _GEN_9774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9776 = 10'h143 == _T_25 ? ram_323 : _GEN_9775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9777 = 10'h144 == _T_25 ? ram_324 : _GEN_9776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9778 = 10'h145 == _T_25 ? ram_325 : _GEN_9777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9779 = 10'h146 == _T_25 ? ram_326 : _GEN_9778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9780 = 10'h147 == _T_25 ? ram_327 : _GEN_9779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9781 = 10'h148 == _T_25 ? ram_328 : _GEN_9780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9782 = 10'h149 == _T_25 ? ram_329 : _GEN_9781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9783 = 10'h14a == _T_25 ? ram_330 : _GEN_9782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9784 = 10'h14b == _T_25 ? ram_331 : _GEN_9783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9785 = 10'h14c == _T_25 ? ram_332 : _GEN_9784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9786 = 10'h14d == _T_25 ? ram_333 : _GEN_9785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9787 = 10'h14e == _T_25 ? ram_334 : _GEN_9786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9788 = 10'h14f == _T_25 ? ram_335 : _GEN_9787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9789 = 10'h150 == _T_25 ? ram_336 : _GEN_9788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9790 = 10'h151 == _T_25 ? ram_337 : _GEN_9789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9791 = 10'h152 == _T_25 ? ram_338 : _GEN_9790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9792 = 10'h153 == _T_25 ? ram_339 : _GEN_9791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9793 = 10'h154 == _T_25 ? ram_340 : _GEN_9792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9794 = 10'h155 == _T_25 ? ram_341 : _GEN_9793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9795 = 10'h156 == _T_25 ? ram_342 : _GEN_9794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9796 = 10'h157 == _T_25 ? ram_343 : _GEN_9795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9797 = 10'h158 == _T_25 ? ram_344 : _GEN_9796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9798 = 10'h159 == _T_25 ? ram_345 : _GEN_9797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9799 = 10'h15a == _T_25 ? ram_346 : _GEN_9798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9800 = 10'h15b == _T_25 ? ram_347 : _GEN_9799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9801 = 10'h15c == _T_25 ? ram_348 : _GEN_9800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9802 = 10'h15d == _T_25 ? ram_349 : _GEN_9801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9803 = 10'h15e == _T_25 ? ram_350 : _GEN_9802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9804 = 10'h15f == _T_25 ? ram_351 : _GEN_9803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9805 = 10'h160 == _T_25 ? ram_352 : _GEN_9804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9806 = 10'h161 == _T_25 ? ram_353 : _GEN_9805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9807 = 10'h162 == _T_25 ? ram_354 : _GEN_9806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9808 = 10'h163 == _T_25 ? ram_355 : _GEN_9807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9809 = 10'h164 == _T_25 ? ram_356 : _GEN_9808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9810 = 10'h165 == _T_25 ? ram_357 : _GEN_9809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9811 = 10'h166 == _T_25 ? ram_358 : _GEN_9810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9812 = 10'h167 == _T_25 ? ram_359 : _GEN_9811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9813 = 10'h168 == _T_25 ? ram_360 : _GEN_9812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9814 = 10'h169 == _T_25 ? ram_361 : _GEN_9813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9815 = 10'h16a == _T_25 ? ram_362 : _GEN_9814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9816 = 10'h16b == _T_25 ? ram_363 : _GEN_9815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9817 = 10'h16c == _T_25 ? ram_364 : _GEN_9816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9818 = 10'h16d == _T_25 ? ram_365 : _GEN_9817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9819 = 10'h16e == _T_25 ? ram_366 : _GEN_9818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9820 = 10'h16f == _T_25 ? ram_367 : _GEN_9819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9821 = 10'h170 == _T_25 ? ram_368 : _GEN_9820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9822 = 10'h171 == _T_25 ? ram_369 : _GEN_9821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9823 = 10'h172 == _T_25 ? ram_370 : _GEN_9822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9824 = 10'h173 == _T_25 ? ram_371 : _GEN_9823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9825 = 10'h174 == _T_25 ? ram_372 : _GEN_9824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9826 = 10'h175 == _T_25 ? ram_373 : _GEN_9825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9827 = 10'h176 == _T_25 ? ram_374 : _GEN_9826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9828 = 10'h177 == _T_25 ? ram_375 : _GEN_9827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9829 = 10'h178 == _T_25 ? ram_376 : _GEN_9828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9830 = 10'h179 == _T_25 ? ram_377 : _GEN_9829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9831 = 10'h17a == _T_25 ? ram_378 : _GEN_9830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9832 = 10'h17b == _T_25 ? ram_379 : _GEN_9831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9833 = 10'h17c == _T_25 ? ram_380 : _GEN_9832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9834 = 10'h17d == _T_25 ? ram_381 : _GEN_9833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9835 = 10'h17e == _T_25 ? ram_382 : _GEN_9834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9836 = 10'h17f == _T_25 ? ram_383 : _GEN_9835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9837 = 10'h180 == _T_25 ? ram_384 : _GEN_9836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9838 = 10'h181 == _T_25 ? ram_385 : _GEN_9837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9839 = 10'h182 == _T_25 ? ram_386 : _GEN_9838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9840 = 10'h183 == _T_25 ? ram_387 : _GEN_9839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9841 = 10'h184 == _T_25 ? ram_388 : _GEN_9840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9842 = 10'h185 == _T_25 ? ram_389 : _GEN_9841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9843 = 10'h186 == _T_25 ? ram_390 : _GEN_9842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9844 = 10'h187 == _T_25 ? ram_391 : _GEN_9843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9845 = 10'h188 == _T_25 ? ram_392 : _GEN_9844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9846 = 10'h189 == _T_25 ? ram_393 : _GEN_9845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9847 = 10'h18a == _T_25 ? ram_394 : _GEN_9846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9848 = 10'h18b == _T_25 ? ram_395 : _GEN_9847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9849 = 10'h18c == _T_25 ? ram_396 : _GEN_9848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9850 = 10'h18d == _T_25 ? ram_397 : _GEN_9849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9851 = 10'h18e == _T_25 ? ram_398 : _GEN_9850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9852 = 10'h18f == _T_25 ? ram_399 : _GEN_9851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9853 = 10'h190 == _T_25 ? ram_400 : _GEN_9852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9854 = 10'h191 == _T_25 ? ram_401 : _GEN_9853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9855 = 10'h192 == _T_25 ? ram_402 : _GEN_9854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9856 = 10'h193 == _T_25 ? ram_403 : _GEN_9855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9857 = 10'h194 == _T_25 ? ram_404 : _GEN_9856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9858 = 10'h195 == _T_25 ? ram_405 : _GEN_9857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9859 = 10'h196 == _T_25 ? ram_406 : _GEN_9858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9860 = 10'h197 == _T_25 ? ram_407 : _GEN_9859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9861 = 10'h198 == _T_25 ? ram_408 : _GEN_9860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9862 = 10'h199 == _T_25 ? ram_409 : _GEN_9861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9863 = 10'h19a == _T_25 ? ram_410 : _GEN_9862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9864 = 10'h19b == _T_25 ? ram_411 : _GEN_9863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9865 = 10'h19c == _T_25 ? ram_412 : _GEN_9864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9866 = 10'h19d == _T_25 ? ram_413 : _GEN_9865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9867 = 10'h19e == _T_25 ? ram_414 : _GEN_9866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9868 = 10'h19f == _T_25 ? ram_415 : _GEN_9867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9869 = 10'h1a0 == _T_25 ? ram_416 : _GEN_9868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9870 = 10'h1a1 == _T_25 ? ram_417 : _GEN_9869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9871 = 10'h1a2 == _T_25 ? ram_418 : _GEN_9870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9872 = 10'h1a3 == _T_25 ? ram_419 : _GEN_9871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9873 = 10'h1a4 == _T_25 ? ram_420 : _GEN_9872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9874 = 10'h1a5 == _T_25 ? ram_421 : _GEN_9873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9875 = 10'h1a6 == _T_25 ? ram_422 : _GEN_9874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9876 = 10'h1a7 == _T_25 ? ram_423 : _GEN_9875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9877 = 10'h1a8 == _T_25 ? ram_424 : _GEN_9876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9878 = 10'h1a9 == _T_25 ? ram_425 : _GEN_9877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9879 = 10'h1aa == _T_25 ? ram_426 : _GEN_9878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9880 = 10'h1ab == _T_25 ? ram_427 : _GEN_9879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9881 = 10'h1ac == _T_25 ? ram_428 : _GEN_9880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9882 = 10'h1ad == _T_25 ? ram_429 : _GEN_9881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9883 = 10'h1ae == _T_25 ? ram_430 : _GEN_9882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9884 = 10'h1af == _T_25 ? ram_431 : _GEN_9883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9885 = 10'h1b0 == _T_25 ? ram_432 : _GEN_9884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9886 = 10'h1b1 == _T_25 ? ram_433 : _GEN_9885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9887 = 10'h1b2 == _T_25 ? ram_434 : _GEN_9886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9888 = 10'h1b3 == _T_25 ? ram_435 : _GEN_9887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9889 = 10'h1b4 == _T_25 ? ram_436 : _GEN_9888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9890 = 10'h1b5 == _T_25 ? ram_437 : _GEN_9889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9891 = 10'h1b6 == _T_25 ? ram_438 : _GEN_9890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9892 = 10'h1b7 == _T_25 ? ram_439 : _GEN_9891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9893 = 10'h1b8 == _T_25 ? ram_440 : _GEN_9892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9894 = 10'h1b9 == _T_25 ? ram_441 : _GEN_9893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9895 = 10'h1ba == _T_25 ? ram_442 : _GEN_9894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9896 = 10'h1bb == _T_25 ? ram_443 : _GEN_9895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9897 = 10'h1bc == _T_25 ? ram_444 : _GEN_9896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9898 = 10'h1bd == _T_25 ? ram_445 : _GEN_9897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9899 = 10'h1be == _T_25 ? ram_446 : _GEN_9898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9900 = 10'h1bf == _T_25 ? ram_447 : _GEN_9899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9901 = 10'h1c0 == _T_25 ? ram_448 : _GEN_9900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9902 = 10'h1c1 == _T_25 ? ram_449 : _GEN_9901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9903 = 10'h1c2 == _T_25 ? ram_450 : _GEN_9902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9904 = 10'h1c3 == _T_25 ? ram_451 : _GEN_9903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9905 = 10'h1c4 == _T_25 ? ram_452 : _GEN_9904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9906 = 10'h1c5 == _T_25 ? ram_453 : _GEN_9905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9907 = 10'h1c6 == _T_25 ? ram_454 : _GEN_9906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9908 = 10'h1c7 == _T_25 ? ram_455 : _GEN_9907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9909 = 10'h1c8 == _T_25 ? ram_456 : _GEN_9908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9910 = 10'h1c9 == _T_25 ? ram_457 : _GEN_9909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9911 = 10'h1ca == _T_25 ? ram_458 : _GEN_9910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9912 = 10'h1cb == _T_25 ? ram_459 : _GEN_9911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9913 = 10'h1cc == _T_25 ? ram_460 : _GEN_9912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9914 = 10'h1cd == _T_25 ? ram_461 : _GEN_9913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9915 = 10'h1ce == _T_25 ? ram_462 : _GEN_9914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9916 = 10'h1cf == _T_25 ? ram_463 : _GEN_9915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9917 = 10'h1d0 == _T_25 ? ram_464 : _GEN_9916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9918 = 10'h1d1 == _T_25 ? ram_465 : _GEN_9917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9919 = 10'h1d2 == _T_25 ? ram_466 : _GEN_9918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9920 = 10'h1d3 == _T_25 ? ram_467 : _GEN_9919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9921 = 10'h1d4 == _T_25 ? ram_468 : _GEN_9920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9922 = 10'h1d5 == _T_25 ? ram_469 : _GEN_9921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9923 = 10'h1d6 == _T_25 ? ram_470 : _GEN_9922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9924 = 10'h1d7 == _T_25 ? ram_471 : _GEN_9923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9925 = 10'h1d8 == _T_25 ? ram_472 : _GEN_9924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9926 = 10'h1d9 == _T_25 ? ram_473 : _GEN_9925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9927 = 10'h1da == _T_25 ? ram_474 : _GEN_9926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9928 = 10'h1db == _T_25 ? ram_475 : _GEN_9927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9929 = 10'h1dc == _T_25 ? ram_476 : _GEN_9928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9930 = 10'h1dd == _T_25 ? ram_477 : _GEN_9929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9931 = 10'h1de == _T_25 ? ram_478 : _GEN_9930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9932 = 10'h1df == _T_25 ? ram_479 : _GEN_9931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9933 = 10'h1e0 == _T_25 ? ram_480 : _GEN_9932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9934 = 10'h1e1 == _T_25 ? ram_481 : _GEN_9933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9935 = 10'h1e2 == _T_25 ? ram_482 : _GEN_9934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9936 = 10'h1e3 == _T_25 ? ram_483 : _GEN_9935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9937 = 10'h1e4 == _T_25 ? ram_484 : _GEN_9936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9938 = 10'h1e5 == _T_25 ? ram_485 : _GEN_9937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9939 = 10'h1e6 == _T_25 ? ram_486 : _GEN_9938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9940 = 10'h1e7 == _T_25 ? ram_487 : _GEN_9939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9941 = 10'h1e8 == _T_25 ? ram_488 : _GEN_9940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9942 = 10'h1e9 == _T_25 ? ram_489 : _GEN_9941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9943 = 10'h1ea == _T_25 ? ram_490 : _GEN_9942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9944 = 10'h1eb == _T_25 ? ram_491 : _GEN_9943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9945 = 10'h1ec == _T_25 ? ram_492 : _GEN_9944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9946 = 10'h1ed == _T_25 ? ram_493 : _GEN_9945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9947 = 10'h1ee == _T_25 ? ram_494 : _GEN_9946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9948 = 10'h1ef == _T_25 ? ram_495 : _GEN_9947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9949 = 10'h1f0 == _T_25 ? ram_496 : _GEN_9948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9950 = 10'h1f1 == _T_25 ? ram_497 : _GEN_9949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9951 = 10'h1f2 == _T_25 ? ram_498 : _GEN_9950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9952 = 10'h1f3 == _T_25 ? ram_499 : _GEN_9951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9953 = 10'h1f4 == _T_25 ? ram_500 : _GEN_9952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9954 = 10'h1f5 == _T_25 ? ram_501 : _GEN_9953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9955 = 10'h1f6 == _T_25 ? ram_502 : _GEN_9954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9956 = 10'h1f7 == _T_25 ? ram_503 : _GEN_9955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9957 = 10'h1f8 == _T_25 ? ram_504 : _GEN_9956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9958 = 10'h1f9 == _T_25 ? ram_505 : _GEN_9957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9959 = 10'h1fa == _T_25 ? ram_506 : _GEN_9958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9960 = 10'h1fb == _T_25 ? ram_507 : _GEN_9959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9961 = 10'h1fc == _T_25 ? ram_508 : _GEN_9960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9962 = 10'h1fd == _T_25 ? ram_509 : _GEN_9961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9963 = 10'h1fe == _T_25 ? ram_510 : _GEN_9962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9964 = 10'h1ff == _T_25 ? ram_511 : _GEN_9963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9965 = 10'h200 == _T_25 ? ram_512 : _GEN_9964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9966 = 10'h201 == _T_25 ? ram_513 : _GEN_9965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9967 = 10'h202 == _T_25 ? ram_514 : _GEN_9966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9968 = 10'h203 == _T_25 ? ram_515 : _GEN_9967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9969 = 10'h204 == _T_25 ? ram_516 : _GEN_9968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9970 = 10'h205 == _T_25 ? ram_517 : _GEN_9969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9971 = 10'h206 == _T_25 ? ram_518 : _GEN_9970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9972 = 10'h207 == _T_25 ? ram_519 : _GEN_9971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9973 = 10'h208 == _T_25 ? ram_520 : _GEN_9972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9974 = 10'h209 == _T_25 ? ram_521 : _GEN_9973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9975 = 10'h20a == _T_25 ? ram_522 : _GEN_9974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9976 = 10'h20b == _T_25 ? ram_523 : _GEN_9975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_9977 = 10'h20c == _T_25 ? ram_524 : _GEN_9976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19079 = {{8190'd0}, _GEN_9977}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_259 = _GEN_19079 ^ _ram_T_258; // @[vga.scala 64:41]
  wire [287:0] _GEN_9978 = 10'h0 == _T_25 ? _ram_T_259[287:0] : _GEN_8928; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9979 = 10'h1 == _T_25 ? _ram_T_259[287:0] : _GEN_8929; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9980 = 10'h2 == _T_25 ? _ram_T_259[287:0] : _GEN_8930; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9981 = 10'h3 == _T_25 ? _ram_T_259[287:0] : _GEN_8931; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9982 = 10'h4 == _T_25 ? _ram_T_259[287:0] : _GEN_8932; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9983 = 10'h5 == _T_25 ? _ram_T_259[287:0] : _GEN_8933; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9984 = 10'h6 == _T_25 ? _ram_T_259[287:0] : _GEN_8934; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9985 = 10'h7 == _T_25 ? _ram_T_259[287:0] : _GEN_8935; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9986 = 10'h8 == _T_25 ? _ram_T_259[287:0] : _GEN_8936; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9987 = 10'h9 == _T_25 ? _ram_T_259[287:0] : _GEN_8937; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9988 = 10'ha == _T_25 ? _ram_T_259[287:0] : _GEN_8938; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9989 = 10'hb == _T_25 ? _ram_T_259[287:0] : _GEN_8939; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9990 = 10'hc == _T_25 ? _ram_T_259[287:0] : _GEN_8940; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9991 = 10'hd == _T_25 ? _ram_T_259[287:0] : _GEN_8941; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9992 = 10'he == _T_25 ? _ram_T_259[287:0] : _GEN_8942; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9993 = 10'hf == _T_25 ? _ram_T_259[287:0] : _GEN_8943; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9994 = 10'h10 == _T_25 ? _ram_T_259[287:0] : _GEN_8944; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9995 = 10'h11 == _T_25 ? _ram_T_259[287:0] : _GEN_8945; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9996 = 10'h12 == _T_25 ? _ram_T_259[287:0] : _GEN_8946; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9997 = 10'h13 == _T_25 ? _ram_T_259[287:0] : _GEN_8947; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9998 = 10'h14 == _T_25 ? _ram_T_259[287:0] : _GEN_8948; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_9999 = 10'h15 == _T_25 ? _ram_T_259[287:0] : _GEN_8949; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10000 = 10'h16 == _T_25 ? _ram_T_259[287:0] : _GEN_8950; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10001 = 10'h17 == _T_25 ? _ram_T_259[287:0] : _GEN_8951; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10002 = 10'h18 == _T_25 ? _ram_T_259[287:0] : _GEN_8952; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10003 = 10'h19 == _T_25 ? _ram_T_259[287:0] : _GEN_8953; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10004 = 10'h1a == _T_25 ? _ram_T_259[287:0] : _GEN_8954; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10005 = 10'h1b == _T_25 ? _ram_T_259[287:0] : _GEN_8955; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10006 = 10'h1c == _T_25 ? _ram_T_259[287:0] : _GEN_8956; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10007 = 10'h1d == _T_25 ? _ram_T_259[287:0] : _GEN_8957; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10008 = 10'h1e == _T_25 ? _ram_T_259[287:0] : _GEN_8958; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10009 = 10'h1f == _T_25 ? _ram_T_259[287:0] : _GEN_8959; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10010 = 10'h20 == _T_25 ? _ram_T_259[287:0] : _GEN_8960; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10011 = 10'h21 == _T_25 ? _ram_T_259[287:0] : _GEN_8961; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10012 = 10'h22 == _T_25 ? _ram_T_259[287:0] : _GEN_8962; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10013 = 10'h23 == _T_25 ? _ram_T_259[287:0] : _GEN_8963; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10014 = 10'h24 == _T_25 ? _ram_T_259[287:0] : _GEN_8964; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10015 = 10'h25 == _T_25 ? _ram_T_259[287:0] : _GEN_8965; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10016 = 10'h26 == _T_25 ? _ram_T_259[287:0] : _GEN_8966; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10017 = 10'h27 == _T_25 ? _ram_T_259[287:0] : _GEN_8967; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10018 = 10'h28 == _T_25 ? _ram_T_259[287:0] : _GEN_8968; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10019 = 10'h29 == _T_25 ? _ram_T_259[287:0] : _GEN_8969; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10020 = 10'h2a == _T_25 ? _ram_T_259[287:0] : _GEN_8970; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10021 = 10'h2b == _T_25 ? _ram_T_259[287:0] : _GEN_8971; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10022 = 10'h2c == _T_25 ? _ram_T_259[287:0] : _GEN_8972; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10023 = 10'h2d == _T_25 ? _ram_T_259[287:0] : _GEN_8973; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10024 = 10'h2e == _T_25 ? _ram_T_259[287:0] : _GEN_8974; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10025 = 10'h2f == _T_25 ? _ram_T_259[287:0] : _GEN_8975; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10026 = 10'h30 == _T_25 ? _ram_T_259[287:0] : _GEN_8976; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10027 = 10'h31 == _T_25 ? _ram_T_259[287:0] : _GEN_8977; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10028 = 10'h32 == _T_25 ? _ram_T_259[287:0] : _GEN_8978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10029 = 10'h33 == _T_25 ? _ram_T_259[287:0] : _GEN_8979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10030 = 10'h34 == _T_25 ? _ram_T_259[287:0] : _GEN_8980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10031 = 10'h35 == _T_25 ? _ram_T_259[287:0] : _GEN_8981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10032 = 10'h36 == _T_25 ? _ram_T_259[287:0] : _GEN_8982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10033 = 10'h37 == _T_25 ? _ram_T_259[287:0] : _GEN_8983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10034 = 10'h38 == _T_25 ? _ram_T_259[287:0] : _GEN_8984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10035 = 10'h39 == _T_25 ? _ram_T_259[287:0] : _GEN_8985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10036 = 10'h3a == _T_25 ? _ram_T_259[287:0] : _GEN_8986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10037 = 10'h3b == _T_25 ? _ram_T_259[287:0] : _GEN_8987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10038 = 10'h3c == _T_25 ? _ram_T_259[287:0] : _GEN_8988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10039 = 10'h3d == _T_25 ? _ram_T_259[287:0] : _GEN_8989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10040 = 10'h3e == _T_25 ? _ram_T_259[287:0] : _GEN_8990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10041 = 10'h3f == _T_25 ? _ram_T_259[287:0] : _GEN_8991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10042 = 10'h40 == _T_25 ? _ram_T_259[287:0] : _GEN_8992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10043 = 10'h41 == _T_25 ? _ram_T_259[287:0] : _GEN_8993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10044 = 10'h42 == _T_25 ? _ram_T_259[287:0] : _GEN_8994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10045 = 10'h43 == _T_25 ? _ram_T_259[287:0] : _GEN_8995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10046 = 10'h44 == _T_25 ? _ram_T_259[287:0] : _GEN_8996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10047 = 10'h45 == _T_25 ? _ram_T_259[287:0] : _GEN_8997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10048 = 10'h46 == _T_25 ? _ram_T_259[287:0] : _GEN_8998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10049 = 10'h47 == _T_25 ? _ram_T_259[287:0] : _GEN_8999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10050 = 10'h48 == _T_25 ? _ram_T_259[287:0] : _GEN_9000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10051 = 10'h49 == _T_25 ? _ram_T_259[287:0] : _GEN_9001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10052 = 10'h4a == _T_25 ? _ram_T_259[287:0] : _GEN_9002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10053 = 10'h4b == _T_25 ? _ram_T_259[287:0] : _GEN_9003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10054 = 10'h4c == _T_25 ? _ram_T_259[287:0] : _GEN_9004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10055 = 10'h4d == _T_25 ? _ram_T_259[287:0] : _GEN_9005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10056 = 10'h4e == _T_25 ? _ram_T_259[287:0] : _GEN_9006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10057 = 10'h4f == _T_25 ? _ram_T_259[287:0] : _GEN_9007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10058 = 10'h50 == _T_25 ? _ram_T_259[287:0] : _GEN_9008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10059 = 10'h51 == _T_25 ? _ram_T_259[287:0] : _GEN_9009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10060 = 10'h52 == _T_25 ? _ram_T_259[287:0] : _GEN_9010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10061 = 10'h53 == _T_25 ? _ram_T_259[287:0] : _GEN_9011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10062 = 10'h54 == _T_25 ? _ram_T_259[287:0] : _GEN_9012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10063 = 10'h55 == _T_25 ? _ram_T_259[287:0] : _GEN_9013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10064 = 10'h56 == _T_25 ? _ram_T_259[287:0] : _GEN_9014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10065 = 10'h57 == _T_25 ? _ram_T_259[287:0] : _GEN_9015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10066 = 10'h58 == _T_25 ? _ram_T_259[287:0] : _GEN_9016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10067 = 10'h59 == _T_25 ? _ram_T_259[287:0] : _GEN_9017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10068 = 10'h5a == _T_25 ? _ram_T_259[287:0] : _GEN_9018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10069 = 10'h5b == _T_25 ? _ram_T_259[287:0] : _GEN_9019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10070 = 10'h5c == _T_25 ? _ram_T_259[287:0] : _GEN_9020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10071 = 10'h5d == _T_25 ? _ram_T_259[287:0] : _GEN_9021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10072 = 10'h5e == _T_25 ? _ram_T_259[287:0] : _GEN_9022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10073 = 10'h5f == _T_25 ? _ram_T_259[287:0] : _GEN_9023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10074 = 10'h60 == _T_25 ? _ram_T_259[287:0] : _GEN_9024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10075 = 10'h61 == _T_25 ? _ram_T_259[287:0] : _GEN_9025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10076 = 10'h62 == _T_25 ? _ram_T_259[287:0] : _GEN_9026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10077 = 10'h63 == _T_25 ? _ram_T_259[287:0] : _GEN_9027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10078 = 10'h64 == _T_25 ? _ram_T_259[287:0] : _GEN_9028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10079 = 10'h65 == _T_25 ? _ram_T_259[287:0] : _GEN_9029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10080 = 10'h66 == _T_25 ? _ram_T_259[287:0] : _GEN_9030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10081 = 10'h67 == _T_25 ? _ram_T_259[287:0] : _GEN_9031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10082 = 10'h68 == _T_25 ? _ram_T_259[287:0] : _GEN_9032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10083 = 10'h69 == _T_25 ? _ram_T_259[287:0] : _GEN_9033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10084 = 10'h6a == _T_25 ? _ram_T_259[287:0] : _GEN_9034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10085 = 10'h6b == _T_25 ? _ram_T_259[287:0] : _GEN_9035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10086 = 10'h6c == _T_25 ? _ram_T_259[287:0] : _GEN_9036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10087 = 10'h6d == _T_25 ? _ram_T_259[287:0] : _GEN_9037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10088 = 10'h6e == _T_25 ? _ram_T_259[287:0] : _GEN_9038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10089 = 10'h6f == _T_25 ? _ram_T_259[287:0] : _GEN_9039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10090 = 10'h70 == _T_25 ? _ram_T_259[287:0] : _GEN_9040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10091 = 10'h71 == _T_25 ? _ram_T_259[287:0] : _GEN_9041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10092 = 10'h72 == _T_25 ? _ram_T_259[287:0] : _GEN_9042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10093 = 10'h73 == _T_25 ? _ram_T_259[287:0] : _GEN_9043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10094 = 10'h74 == _T_25 ? _ram_T_259[287:0] : _GEN_9044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10095 = 10'h75 == _T_25 ? _ram_T_259[287:0] : _GEN_9045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10096 = 10'h76 == _T_25 ? _ram_T_259[287:0] : _GEN_9046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10097 = 10'h77 == _T_25 ? _ram_T_259[287:0] : _GEN_9047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10098 = 10'h78 == _T_25 ? _ram_T_259[287:0] : _GEN_9048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10099 = 10'h79 == _T_25 ? _ram_T_259[287:0] : _GEN_9049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10100 = 10'h7a == _T_25 ? _ram_T_259[287:0] : _GEN_9050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10101 = 10'h7b == _T_25 ? _ram_T_259[287:0] : _GEN_9051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10102 = 10'h7c == _T_25 ? _ram_T_259[287:0] : _GEN_9052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10103 = 10'h7d == _T_25 ? _ram_T_259[287:0] : _GEN_9053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10104 = 10'h7e == _T_25 ? _ram_T_259[287:0] : _GEN_9054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10105 = 10'h7f == _T_25 ? _ram_T_259[287:0] : _GEN_9055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10106 = 10'h80 == _T_25 ? _ram_T_259[287:0] : _GEN_9056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10107 = 10'h81 == _T_25 ? _ram_T_259[287:0] : _GEN_9057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10108 = 10'h82 == _T_25 ? _ram_T_259[287:0] : _GEN_9058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10109 = 10'h83 == _T_25 ? _ram_T_259[287:0] : _GEN_9059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10110 = 10'h84 == _T_25 ? _ram_T_259[287:0] : _GEN_9060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10111 = 10'h85 == _T_25 ? _ram_T_259[287:0] : _GEN_9061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10112 = 10'h86 == _T_25 ? _ram_T_259[287:0] : _GEN_9062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10113 = 10'h87 == _T_25 ? _ram_T_259[287:0] : _GEN_9063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10114 = 10'h88 == _T_25 ? _ram_T_259[287:0] : _GEN_9064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10115 = 10'h89 == _T_25 ? _ram_T_259[287:0] : _GEN_9065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10116 = 10'h8a == _T_25 ? _ram_T_259[287:0] : _GEN_9066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10117 = 10'h8b == _T_25 ? _ram_T_259[287:0] : _GEN_9067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10118 = 10'h8c == _T_25 ? _ram_T_259[287:0] : _GEN_9068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10119 = 10'h8d == _T_25 ? _ram_T_259[287:0] : _GEN_9069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10120 = 10'h8e == _T_25 ? _ram_T_259[287:0] : _GEN_9070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10121 = 10'h8f == _T_25 ? _ram_T_259[287:0] : _GEN_9071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10122 = 10'h90 == _T_25 ? _ram_T_259[287:0] : _GEN_9072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10123 = 10'h91 == _T_25 ? _ram_T_259[287:0] : _GEN_9073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10124 = 10'h92 == _T_25 ? _ram_T_259[287:0] : _GEN_9074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10125 = 10'h93 == _T_25 ? _ram_T_259[287:0] : _GEN_9075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10126 = 10'h94 == _T_25 ? _ram_T_259[287:0] : _GEN_9076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10127 = 10'h95 == _T_25 ? _ram_T_259[287:0] : _GEN_9077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10128 = 10'h96 == _T_25 ? _ram_T_259[287:0] : _GEN_9078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10129 = 10'h97 == _T_25 ? _ram_T_259[287:0] : _GEN_9079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10130 = 10'h98 == _T_25 ? _ram_T_259[287:0] : _GEN_9080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10131 = 10'h99 == _T_25 ? _ram_T_259[287:0] : _GEN_9081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10132 = 10'h9a == _T_25 ? _ram_T_259[287:0] : _GEN_9082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10133 = 10'h9b == _T_25 ? _ram_T_259[287:0] : _GEN_9083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10134 = 10'h9c == _T_25 ? _ram_T_259[287:0] : _GEN_9084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10135 = 10'h9d == _T_25 ? _ram_T_259[287:0] : _GEN_9085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10136 = 10'h9e == _T_25 ? _ram_T_259[287:0] : _GEN_9086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10137 = 10'h9f == _T_25 ? _ram_T_259[287:0] : _GEN_9087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10138 = 10'ha0 == _T_25 ? _ram_T_259[287:0] : _GEN_9088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10139 = 10'ha1 == _T_25 ? _ram_T_259[287:0] : _GEN_9089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10140 = 10'ha2 == _T_25 ? _ram_T_259[287:0] : _GEN_9090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10141 = 10'ha3 == _T_25 ? _ram_T_259[287:0] : _GEN_9091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10142 = 10'ha4 == _T_25 ? _ram_T_259[287:0] : _GEN_9092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10143 = 10'ha5 == _T_25 ? _ram_T_259[287:0] : _GEN_9093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10144 = 10'ha6 == _T_25 ? _ram_T_259[287:0] : _GEN_9094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10145 = 10'ha7 == _T_25 ? _ram_T_259[287:0] : _GEN_9095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10146 = 10'ha8 == _T_25 ? _ram_T_259[287:0] : _GEN_9096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10147 = 10'ha9 == _T_25 ? _ram_T_259[287:0] : _GEN_9097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10148 = 10'haa == _T_25 ? _ram_T_259[287:0] : _GEN_9098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10149 = 10'hab == _T_25 ? _ram_T_259[287:0] : _GEN_9099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10150 = 10'hac == _T_25 ? _ram_T_259[287:0] : _GEN_9100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10151 = 10'had == _T_25 ? _ram_T_259[287:0] : _GEN_9101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10152 = 10'hae == _T_25 ? _ram_T_259[287:0] : _GEN_9102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10153 = 10'haf == _T_25 ? _ram_T_259[287:0] : _GEN_9103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10154 = 10'hb0 == _T_25 ? _ram_T_259[287:0] : _GEN_9104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10155 = 10'hb1 == _T_25 ? _ram_T_259[287:0] : _GEN_9105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10156 = 10'hb2 == _T_25 ? _ram_T_259[287:0] : _GEN_9106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10157 = 10'hb3 == _T_25 ? _ram_T_259[287:0] : _GEN_9107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10158 = 10'hb4 == _T_25 ? _ram_T_259[287:0] : _GEN_9108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10159 = 10'hb5 == _T_25 ? _ram_T_259[287:0] : _GEN_9109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10160 = 10'hb6 == _T_25 ? _ram_T_259[287:0] : _GEN_9110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10161 = 10'hb7 == _T_25 ? _ram_T_259[287:0] : _GEN_9111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10162 = 10'hb8 == _T_25 ? _ram_T_259[287:0] : _GEN_9112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10163 = 10'hb9 == _T_25 ? _ram_T_259[287:0] : _GEN_9113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10164 = 10'hba == _T_25 ? _ram_T_259[287:0] : _GEN_9114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10165 = 10'hbb == _T_25 ? _ram_T_259[287:0] : _GEN_9115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10166 = 10'hbc == _T_25 ? _ram_T_259[287:0] : _GEN_9116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10167 = 10'hbd == _T_25 ? _ram_T_259[287:0] : _GEN_9117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10168 = 10'hbe == _T_25 ? _ram_T_259[287:0] : _GEN_9118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10169 = 10'hbf == _T_25 ? _ram_T_259[287:0] : _GEN_9119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10170 = 10'hc0 == _T_25 ? _ram_T_259[287:0] : _GEN_9120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10171 = 10'hc1 == _T_25 ? _ram_T_259[287:0] : _GEN_9121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10172 = 10'hc2 == _T_25 ? _ram_T_259[287:0] : _GEN_9122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10173 = 10'hc3 == _T_25 ? _ram_T_259[287:0] : _GEN_9123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10174 = 10'hc4 == _T_25 ? _ram_T_259[287:0] : _GEN_9124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10175 = 10'hc5 == _T_25 ? _ram_T_259[287:0] : _GEN_9125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10176 = 10'hc6 == _T_25 ? _ram_T_259[287:0] : _GEN_9126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10177 = 10'hc7 == _T_25 ? _ram_T_259[287:0] : _GEN_9127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10178 = 10'hc8 == _T_25 ? _ram_T_259[287:0] : _GEN_9128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10179 = 10'hc9 == _T_25 ? _ram_T_259[287:0] : _GEN_9129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10180 = 10'hca == _T_25 ? _ram_T_259[287:0] : _GEN_9130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10181 = 10'hcb == _T_25 ? _ram_T_259[287:0] : _GEN_9131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10182 = 10'hcc == _T_25 ? _ram_T_259[287:0] : _GEN_9132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10183 = 10'hcd == _T_25 ? _ram_T_259[287:0] : _GEN_9133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10184 = 10'hce == _T_25 ? _ram_T_259[287:0] : _GEN_9134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10185 = 10'hcf == _T_25 ? _ram_T_259[287:0] : _GEN_9135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10186 = 10'hd0 == _T_25 ? _ram_T_259[287:0] : _GEN_9136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10187 = 10'hd1 == _T_25 ? _ram_T_259[287:0] : _GEN_9137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10188 = 10'hd2 == _T_25 ? _ram_T_259[287:0] : _GEN_9138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10189 = 10'hd3 == _T_25 ? _ram_T_259[287:0] : _GEN_9139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10190 = 10'hd4 == _T_25 ? _ram_T_259[287:0] : _GEN_9140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10191 = 10'hd5 == _T_25 ? _ram_T_259[287:0] : _GEN_9141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10192 = 10'hd6 == _T_25 ? _ram_T_259[287:0] : _GEN_9142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10193 = 10'hd7 == _T_25 ? _ram_T_259[287:0] : _GEN_9143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10194 = 10'hd8 == _T_25 ? _ram_T_259[287:0] : _GEN_9144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10195 = 10'hd9 == _T_25 ? _ram_T_259[287:0] : _GEN_9145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10196 = 10'hda == _T_25 ? _ram_T_259[287:0] : _GEN_9146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10197 = 10'hdb == _T_25 ? _ram_T_259[287:0] : _GEN_9147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10198 = 10'hdc == _T_25 ? _ram_T_259[287:0] : _GEN_9148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10199 = 10'hdd == _T_25 ? _ram_T_259[287:0] : _GEN_9149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10200 = 10'hde == _T_25 ? _ram_T_259[287:0] : _GEN_9150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10201 = 10'hdf == _T_25 ? _ram_T_259[287:0] : _GEN_9151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10202 = 10'he0 == _T_25 ? _ram_T_259[287:0] : _GEN_9152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10203 = 10'he1 == _T_25 ? _ram_T_259[287:0] : _GEN_9153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10204 = 10'he2 == _T_25 ? _ram_T_259[287:0] : _GEN_9154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10205 = 10'he3 == _T_25 ? _ram_T_259[287:0] : _GEN_9155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10206 = 10'he4 == _T_25 ? _ram_T_259[287:0] : _GEN_9156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10207 = 10'he5 == _T_25 ? _ram_T_259[287:0] : _GEN_9157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10208 = 10'he6 == _T_25 ? _ram_T_259[287:0] : _GEN_9158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10209 = 10'he7 == _T_25 ? _ram_T_259[287:0] : _GEN_9159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10210 = 10'he8 == _T_25 ? _ram_T_259[287:0] : _GEN_9160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10211 = 10'he9 == _T_25 ? _ram_T_259[287:0] : _GEN_9161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10212 = 10'hea == _T_25 ? _ram_T_259[287:0] : _GEN_9162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10213 = 10'heb == _T_25 ? _ram_T_259[287:0] : _GEN_9163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10214 = 10'hec == _T_25 ? _ram_T_259[287:0] : _GEN_9164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10215 = 10'hed == _T_25 ? _ram_T_259[287:0] : _GEN_9165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10216 = 10'hee == _T_25 ? _ram_T_259[287:0] : _GEN_9166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10217 = 10'hef == _T_25 ? _ram_T_259[287:0] : _GEN_9167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10218 = 10'hf0 == _T_25 ? _ram_T_259[287:0] : _GEN_9168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10219 = 10'hf1 == _T_25 ? _ram_T_259[287:0] : _GEN_9169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10220 = 10'hf2 == _T_25 ? _ram_T_259[287:0] : _GEN_9170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10221 = 10'hf3 == _T_25 ? _ram_T_259[287:0] : _GEN_9171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10222 = 10'hf4 == _T_25 ? _ram_T_259[287:0] : _GEN_9172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10223 = 10'hf5 == _T_25 ? _ram_T_259[287:0] : _GEN_9173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10224 = 10'hf6 == _T_25 ? _ram_T_259[287:0] : _GEN_9174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10225 = 10'hf7 == _T_25 ? _ram_T_259[287:0] : _GEN_9175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10226 = 10'hf8 == _T_25 ? _ram_T_259[287:0] : _GEN_9176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10227 = 10'hf9 == _T_25 ? _ram_T_259[287:0] : _GEN_9177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10228 = 10'hfa == _T_25 ? _ram_T_259[287:0] : _GEN_9178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10229 = 10'hfb == _T_25 ? _ram_T_259[287:0] : _GEN_9179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10230 = 10'hfc == _T_25 ? _ram_T_259[287:0] : _GEN_9180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10231 = 10'hfd == _T_25 ? _ram_T_259[287:0] : _GEN_9181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10232 = 10'hfe == _T_25 ? _ram_T_259[287:0] : _GEN_9182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10233 = 10'hff == _T_25 ? _ram_T_259[287:0] : _GEN_9183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10234 = 10'h100 == _T_25 ? _ram_T_259[287:0] : _GEN_9184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10235 = 10'h101 == _T_25 ? _ram_T_259[287:0] : _GEN_9185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10236 = 10'h102 == _T_25 ? _ram_T_259[287:0] : _GEN_9186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10237 = 10'h103 == _T_25 ? _ram_T_259[287:0] : _GEN_9187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10238 = 10'h104 == _T_25 ? _ram_T_259[287:0] : _GEN_9188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10239 = 10'h105 == _T_25 ? _ram_T_259[287:0] : _GEN_9189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10240 = 10'h106 == _T_25 ? _ram_T_259[287:0] : _GEN_9190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10241 = 10'h107 == _T_25 ? _ram_T_259[287:0] : _GEN_9191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10242 = 10'h108 == _T_25 ? _ram_T_259[287:0] : _GEN_9192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10243 = 10'h109 == _T_25 ? _ram_T_259[287:0] : _GEN_9193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10244 = 10'h10a == _T_25 ? _ram_T_259[287:0] : _GEN_9194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10245 = 10'h10b == _T_25 ? _ram_T_259[287:0] : _GEN_9195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10246 = 10'h10c == _T_25 ? _ram_T_259[287:0] : _GEN_9196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10247 = 10'h10d == _T_25 ? _ram_T_259[287:0] : _GEN_9197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10248 = 10'h10e == _T_25 ? _ram_T_259[287:0] : _GEN_9198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10249 = 10'h10f == _T_25 ? _ram_T_259[287:0] : _GEN_9199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10250 = 10'h110 == _T_25 ? _ram_T_259[287:0] : _GEN_9200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10251 = 10'h111 == _T_25 ? _ram_T_259[287:0] : _GEN_9201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10252 = 10'h112 == _T_25 ? _ram_T_259[287:0] : _GEN_9202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10253 = 10'h113 == _T_25 ? _ram_T_259[287:0] : _GEN_9203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10254 = 10'h114 == _T_25 ? _ram_T_259[287:0] : _GEN_9204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10255 = 10'h115 == _T_25 ? _ram_T_259[287:0] : _GEN_9205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10256 = 10'h116 == _T_25 ? _ram_T_259[287:0] : _GEN_9206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10257 = 10'h117 == _T_25 ? _ram_T_259[287:0] : _GEN_9207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10258 = 10'h118 == _T_25 ? _ram_T_259[287:0] : _GEN_9208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10259 = 10'h119 == _T_25 ? _ram_T_259[287:0] : _GEN_9209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10260 = 10'h11a == _T_25 ? _ram_T_259[287:0] : _GEN_9210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10261 = 10'h11b == _T_25 ? _ram_T_259[287:0] : _GEN_9211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10262 = 10'h11c == _T_25 ? _ram_T_259[287:0] : _GEN_9212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10263 = 10'h11d == _T_25 ? _ram_T_259[287:0] : _GEN_9213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10264 = 10'h11e == _T_25 ? _ram_T_259[287:0] : _GEN_9214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10265 = 10'h11f == _T_25 ? _ram_T_259[287:0] : _GEN_9215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10266 = 10'h120 == _T_25 ? _ram_T_259[287:0] : _GEN_9216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10267 = 10'h121 == _T_25 ? _ram_T_259[287:0] : _GEN_9217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10268 = 10'h122 == _T_25 ? _ram_T_259[287:0] : _GEN_9218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10269 = 10'h123 == _T_25 ? _ram_T_259[287:0] : _GEN_9219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10270 = 10'h124 == _T_25 ? _ram_T_259[287:0] : _GEN_9220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10271 = 10'h125 == _T_25 ? _ram_T_259[287:0] : _GEN_9221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10272 = 10'h126 == _T_25 ? _ram_T_259[287:0] : _GEN_9222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10273 = 10'h127 == _T_25 ? _ram_T_259[287:0] : _GEN_9223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10274 = 10'h128 == _T_25 ? _ram_T_259[287:0] : _GEN_9224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10275 = 10'h129 == _T_25 ? _ram_T_259[287:0] : _GEN_9225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10276 = 10'h12a == _T_25 ? _ram_T_259[287:0] : _GEN_9226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10277 = 10'h12b == _T_25 ? _ram_T_259[287:0] : _GEN_9227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10278 = 10'h12c == _T_25 ? _ram_T_259[287:0] : _GEN_9228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10279 = 10'h12d == _T_25 ? _ram_T_259[287:0] : _GEN_9229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10280 = 10'h12e == _T_25 ? _ram_T_259[287:0] : _GEN_9230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10281 = 10'h12f == _T_25 ? _ram_T_259[287:0] : _GEN_9231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10282 = 10'h130 == _T_25 ? _ram_T_259[287:0] : _GEN_9232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10283 = 10'h131 == _T_25 ? _ram_T_259[287:0] : _GEN_9233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10284 = 10'h132 == _T_25 ? _ram_T_259[287:0] : _GEN_9234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10285 = 10'h133 == _T_25 ? _ram_T_259[287:0] : _GEN_9235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10286 = 10'h134 == _T_25 ? _ram_T_259[287:0] : _GEN_9236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10287 = 10'h135 == _T_25 ? _ram_T_259[287:0] : _GEN_9237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10288 = 10'h136 == _T_25 ? _ram_T_259[287:0] : _GEN_9238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10289 = 10'h137 == _T_25 ? _ram_T_259[287:0] : _GEN_9239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10290 = 10'h138 == _T_25 ? _ram_T_259[287:0] : _GEN_9240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10291 = 10'h139 == _T_25 ? _ram_T_259[287:0] : _GEN_9241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10292 = 10'h13a == _T_25 ? _ram_T_259[287:0] : _GEN_9242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10293 = 10'h13b == _T_25 ? _ram_T_259[287:0] : _GEN_9243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10294 = 10'h13c == _T_25 ? _ram_T_259[287:0] : _GEN_9244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10295 = 10'h13d == _T_25 ? _ram_T_259[287:0] : _GEN_9245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10296 = 10'h13e == _T_25 ? _ram_T_259[287:0] : _GEN_9246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10297 = 10'h13f == _T_25 ? _ram_T_259[287:0] : _GEN_9247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10298 = 10'h140 == _T_25 ? _ram_T_259[287:0] : _GEN_9248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10299 = 10'h141 == _T_25 ? _ram_T_259[287:0] : _GEN_9249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10300 = 10'h142 == _T_25 ? _ram_T_259[287:0] : _GEN_9250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10301 = 10'h143 == _T_25 ? _ram_T_259[287:0] : _GEN_9251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10302 = 10'h144 == _T_25 ? _ram_T_259[287:0] : _GEN_9252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10303 = 10'h145 == _T_25 ? _ram_T_259[287:0] : _GEN_9253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10304 = 10'h146 == _T_25 ? _ram_T_259[287:0] : _GEN_9254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10305 = 10'h147 == _T_25 ? _ram_T_259[287:0] : _GEN_9255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10306 = 10'h148 == _T_25 ? _ram_T_259[287:0] : _GEN_9256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10307 = 10'h149 == _T_25 ? _ram_T_259[287:0] : _GEN_9257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10308 = 10'h14a == _T_25 ? _ram_T_259[287:0] : _GEN_9258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10309 = 10'h14b == _T_25 ? _ram_T_259[287:0] : _GEN_9259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10310 = 10'h14c == _T_25 ? _ram_T_259[287:0] : _GEN_9260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10311 = 10'h14d == _T_25 ? _ram_T_259[287:0] : _GEN_9261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10312 = 10'h14e == _T_25 ? _ram_T_259[287:0] : _GEN_9262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10313 = 10'h14f == _T_25 ? _ram_T_259[287:0] : _GEN_9263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10314 = 10'h150 == _T_25 ? _ram_T_259[287:0] : _GEN_9264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10315 = 10'h151 == _T_25 ? _ram_T_259[287:0] : _GEN_9265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10316 = 10'h152 == _T_25 ? _ram_T_259[287:0] : _GEN_9266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10317 = 10'h153 == _T_25 ? _ram_T_259[287:0] : _GEN_9267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10318 = 10'h154 == _T_25 ? _ram_T_259[287:0] : _GEN_9268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10319 = 10'h155 == _T_25 ? _ram_T_259[287:0] : _GEN_9269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10320 = 10'h156 == _T_25 ? _ram_T_259[287:0] : _GEN_9270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10321 = 10'h157 == _T_25 ? _ram_T_259[287:0] : _GEN_9271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10322 = 10'h158 == _T_25 ? _ram_T_259[287:0] : _GEN_9272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10323 = 10'h159 == _T_25 ? _ram_T_259[287:0] : _GEN_9273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10324 = 10'h15a == _T_25 ? _ram_T_259[287:0] : _GEN_9274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10325 = 10'h15b == _T_25 ? _ram_T_259[287:0] : _GEN_9275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10326 = 10'h15c == _T_25 ? _ram_T_259[287:0] : _GEN_9276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10327 = 10'h15d == _T_25 ? _ram_T_259[287:0] : _GEN_9277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10328 = 10'h15e == _T_25 ? _ram_T_259[287:0] : _GEN_9278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10329 = 10'h15f == _T_25 ? _ram_T_259[287:0] : _GEN_9279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10330 = 10'h160 == _T_25 ? _ram_T_259[287:0] : _GEN_9280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10331 = 10'h161 == _T_25 ? _ram_T_259[287:0] : _GEN_9281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10332 = 10'h162 == _T_25 ? _ram_T_259[287:0] : _GEN_9282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10333 = 10'h163 == _T_25 ? _ram_T_259[287:0] : _GEN_9283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10334 = 10'h164 == _T_25 ? _ram_T_259[287:0] : _GEN_9284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10335 = 10'h165 == _T_25 ? _ram_T_259[287:0] : _GEN_9285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10336 = 10'h166 == _T_25 ? _ram_T_259[287:0] : _GEN_9286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10337 = 10'h167 == _T_25 ? _ram_T_259[287:0] : _GEN_9287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10338 = 10'h168 == _T_25 ? _ram_T_259[287:0] : _GEN_9288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10339 = 10'h169 == _T_25 ? _ram_T_259[287:0] : _GEN_9289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10340 = 10'h16a == _T_25 ? _ram_T_259[287:0] : _GEN_9290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10341 = 10'h16b == _T_25 ? _ram_T_259[287:0] : _GEN_9291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10342 = 10'h16c == _T_25 ? _ram_T_259[287:0] : _GEN_9292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10343 = 10'h16d == _T_25 ? _ram_T_259[287:0] : _GEN_9293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10344 = 10'h16e == _T_25 ? _ram_T_259[287:0] : _GEN_9294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10345 = 10'h16f == _T_25 ? _ram_T_259[287:0] : _GEN_9295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10346 = 10'h170 == _T_25 ? _ram_T_259[287:0] : _GEN_9296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10347 = 10'h171 == _T_25 ? _ram_T_259[287:0] : _GEN_9297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10348 = 10'h172 == _T_25 ? _ram_T_259[287:0] : _GEN_9298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10349 = 10'h173 == _T_25 ? _ram_T_259[287:0] : _GEN_9299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10350 = 10'h174 == _T_25 ? _ram_T_259[287:0] : _GEN_9300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10351 = 10'h175 == _T_25 ? _ram_T_259[287:0] : _GEN_9301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10352 = 10'h176 == _T_25 ? _ram_T_259[287:0] : _GEN_9302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10353 = 10'h177 == _T_25 ? _ram_T_259[287:0] : _GEN_9303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10354 = 10'h178 == _T_25 ? _ram_T_259[287:0] : _GEN_9304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10355 = 10'h179 == _T_25 ? _ram_T_259[287:0] : _GEN_9305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10356 = 10'h17a == _T_25 ? _ram_T_259[287:0] : _GEN_9306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10357 = 10'h17b == _T_25 ? _ram_T_259[287:0] : _GEN_9307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10358 = 10'h17c == _T_25 ? _ram_T_259[287:0] : _GEN_9308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10359 = 10'h17d == _T_25 ? _ram_T_259[287:0] : _GEN_9309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10360 = 10'h17e == _T_25 ? _ram_T_259[287:0] : _GEN_9310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10361 = 10'h17f == _T_25 ? _ram_T_259[287:0] : _GEN_9311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10362 = 10'h180 == _T_25 ? _ram_T_259[287:0] : _GEN_9312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10363 = 10'h181 == _T_25 ? _ram_T_259[287:0] : _GEN_9313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10364 = 10'h182 == _T_25 ? _ram_T_259[287:0] : _GEN_9314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10365 = 10'h183 == _T_25 ? _ram_T_259[287:0] : _GEN_9315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10366 = 10'h184 == _T_25 ? _ram_T_259[287:0] : _GEN_9316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10367 = 10'h185 == _T_25 ? _ram_T_259[287:0] : _GEN_9317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10368 = 10'h186 == _T_25 ? _ram_T_259[287:0] : _GEN_9318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10369 = 10'h187 == _T_25 ? _ram_T_259[287:0] : _GEN_9319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10370 = 10'h188 == _T_25 ? _ram_T_259[287:0] : _GEN_9320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10371 = 10'h189 == _T_25 ? _ram_T_259[287:0] : _GEN_9321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10372 = 10'h18a == _T_25 ? _ram_T_259[287:0] : _GEN_9322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10373 = 10'h18b == _T_25 ? _ram_T_259[287:0] : _GEN_9323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10374 = 10'h18c == _T_25 ? _ram_T_259[287:0] : _GEN_9324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10375 = 10'h18d == _T_25 ? _ram_T_259[287:0] : _GEN_9325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10376 = 10'h18e == _T_25 ? _ram_T_259[287:0] : _GEN_9326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10377 = 10'h18f == _T_25 ? _ram_T_259[287:0] : _GEN_9327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10378 = 10'h190 == _T_25 ? _ram_T_259[287:0] : _GEN_9328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10379 = 10'h191 == _T_25 ? _ram_T_259[287:0] : _GEN_9329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10380 = 10'h192 == _T_25 ? _ram_T_259[287:0] : _GEN_9330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10381 = 10'h193 == _T_25 ? _ram_T_259[287:0] : _GEN_9331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10382 = 10'h194 == _T_25 ? _ram_T_259[287:0] : _GEN_9332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10383 = 10'h195 == _T_25 ? _ram_T_259[287:0] : _GEN_9333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10384 = 10'h196 == _T_25 ? _ram_T_259[287:0] : _GEN_9334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10385 = 10'h197 == _T_25 ? _ram_T_259[287:0] : _GEN_9335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10386 = 10'h198 == _T_25 ? _ram_T_259[287:0] : _GEN_9336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10387 = 10'h199 == _T_25 ? _ram_T_259[287:0] : _GEN_9337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10388 = 10'h19a == _T_25 ? _ram_T_259[287:0] : _GEN_9338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10389 = 10'h19b == _T_25 ? _ram_T_259[287:0] : _GEN_9339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10390 = 10'h19c == _T_25 ? _ram_T_259[287:0] : _GEN_9340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10391 = 10'h19d == _T_25 ? _ram_T_259[287:0] : _GEN_9341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10392 = 10'h19e == _T_25 ? _ram_T_259[287:0] : _GEN_9342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10393 = 10'h19f == _T_25 ? _ram_T_259[287:0] : _GEN_9343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10394 = 10'h1a0 == _T_25 ? _ram_T_259[287:0] : _GEN_9344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10395 = 10'h1a1 == _T_25 ? _ram_T_259[287:0] : _GEN_9345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10396 = 10'h1a2 == _T_25 ? _ram_T_259[287:0] : _GEN_9346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10397 = 10'h1a3 == _T_25 ? _ram_T_259[287:0] : _GEN_9347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10398 = 10'h1a4 == _T_25 ? _ram_T_259[287:0] : _GEN_9348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10399 = 10'h1a5 == _T_25 ? _ram_T_259[287:0] : _GEN_9349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10400 = 10'h1a6 == _T_25 ? _ram_T_259[287:0] : _GEN_9350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10401 = 10'h1a7 == _T_25 ? _ram_T_259[287:0] : _GEN_9351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10402 = 10'h1a8 == _T_25 ? _ram_T_259[287:0] : _GEN_9352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10403 = 10'h1a9 == _T_25 ? _ram_T_259[287:0] : _GEN_9353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10404 = 10'h1aa == _T_25 ? _ram_T_259[287:0] : _GEN_9354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10405 = 10'h1ab == _T_25 ? _ram_T_259[287:0] : _GEN_9355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10406 = 10'h1ac == _T_25 ? _ram_T_259[287:0] : _GEN_9356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10407 = 10'h1ad == _T_25 ? _ram_T_259[287:0] : _GEN_9357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10408 = 10'h1ae == _T_25 ? _ram_T_259[287:0] : _GEN_9358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10409 = 10'h1af == _T_25 ? _ram_T_259[287:0] : _GEN_9359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10410 = 10'h1b0 == _T_25 ? _ram_T_259[287:0] : _GEN_9360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10411 = 10'h1b1 == _T_25 ? _ram_T_259[287:0] : _GEN_9361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10412 = 10'h1b2 == _T_25 ? _ram_T_259[287:0] : _GEN_9362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10413 = 10'h1b3 == _T_25 ? _ram_T_259[287:0] : _GEN_9363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10414 = 10'h1b4 == _T_25 ? _ram_T_259[287:0] : _GEN_9364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10415 = 10'h1b5 == _T_25 ? _ram_T_259[287:0] : _GEN_9365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10416 = 10'h1b6 == _T_25 ? _ram_T_259[287:0] : _GEN_9366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10417 = 10'h1b7 == _T_25 ? _ram_T_259[287:0] : _GEN_9367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10418 = 10'h1b8 == _T_25 ? _ram_T_259[287:0] : _GEN_9368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10419 = 10'h1b9 == _T_25 ? _ram_T_259[287:0] : _GEN_9369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10420 = 10'h1ba == _T_25 ? _ram_T_259[287:0] : _GEN_9370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10421 = 10'h1bb == _T_25 ? _ram_T_259[287:0] : _GEN_9371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10422 = 10'h1bc == _T_25 ? _ram_T_259[287:0] : _GEN_9372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10423 = 10'h1bd == _T_25 ? _ram_T_259[287:0] : _GEN_9373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10424 = 10'h1be == _T_25 ? _ram_T_259[287:0] : _GEN_9374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10425 = 10'h1bf == _T_25 ? _ram_T_259[287:0] : _GEN_9375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10426 = 10'h1c0 == _T_25 ? _ram_T_259[287:0] : _GEN_9376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10427 = 10'h1c1 == _T_25 ? _ram_T_259[287:0] : _GEN_9377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10428 = 10'h1c2 == _T_25 ? _ram_T_259[287:0] : _GEN_9378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10429 = 10'h1c3 == _T_25 ? _ram_T_259[287:0] : _GEN_9379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10430 = 10'h1c4 == _T_25 ? _ram_T_259[287:0] : _GEN_9380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10431 = 10'h1c5 == _T_25 ? _ram_T_259[287:0] : _GEN_9381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10432 = 10'h1c6 == _T_25 ? _ram_T_259[287:0] : _GEN_9382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10433 = 10'h1c7 == _T_25 ? _ram_T_259[287:0] : _GEN_9383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10434 = 10'h1c8 == _T_25 ? _ram_T_259[287:0] : _GEN_9384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10435 = 10'h1c9 == _T_25 ? _ram_T_259[287:0] : _GEN_9385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10436 = 10'h1ca == _T_25 ? _ram_T_259[287:0] : _GEN_9386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10437 = 10'h1cb == _T_25 ? _ram_T_259[287:0] : _GEN_9387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10438 = 10'h1cc == _T_25 ? _ram_T_259[287:0] : _GEN_9388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10439 = 10'h1cd == _T_25 ? _ram_T_259[287:0] : _GEN_9389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10440 = 10'h1ce == _T_25 ? _ram_T_259[287:0] : _GEN_9390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10441 = 10'h1cf == _T_25 ? _ram_T_259[287:0] : _GEN_9391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10442 = 10'h1d0 == _T_25 ? _ram_T_259[287:0] : _GEN_9392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10443 = 10'h1d1 == _T_25 ? _ram_T_259[287:0] : _GEN_9393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10444 = 10'h1d2 == _T_25 ? _ram_T_259[287:0] : _GEN_9394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10445 = 10'h1d3 == _T_25 ? _ram_T_259[287:0] : _GEN_9395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10446 = 10'h1d4 == _T_25 ? _ram_T_259[287:0] : _GEN_9396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10447 = 10'h1d5 == _T_25 ? _ram_T_259[287:0] : _GEN_9397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10448 = 10'h1d6 == _T_25 ? _ram_T_259[287:0] : _GEN_9398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10449 = 10'h1d7 == _T_25 ? _ram_T_259[287:0] : _GEN_9399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10450 = 10'h1d8 == _T_25 ? _ram_T_259[287:0] : _GEN_9400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10451 = 10'h1d9 == _T_25 ? _ram_T_259[287:0] : _GEN_9401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10452 = 10'h1da == _T_25 ? _ram_T_259[287:0] : _GEN_9402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10453 = 10'h1db == _T_25 ? _ram_T_259[287:0] : _GEN_9403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10454 = 10'h1dc == _T_25 ? _ram_T_259[287:0] : _GEN_9404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10455 = 10'h1dd == _T_25 ? _ram_T_259[287:0] : _GEN_9405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10456 = 10'h1de == _T_25 ? _ram_T_259[287:0] : _GEN_9406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10457 = 10'h1df == _T_25 ? _ram_T_259[287:0] : _GEN_9407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10458 = 10'h1e0 == _T_25 ? _ram_T_259[287:0] : _GEN_9408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10459 = 10'h1e1 == _T_25 ? _ram_T_259[287:0] : _GEN_9409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10460 = 10'h1e2 == _T_25 ? _ram_T_259[287:0] : _GEN_9410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10461 = 10'h1e3 == _T_25 ? _ram_T_259[287:0] : _GEN_9411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10462 = 10'h1e4 == _T_25 ? _ram_T_259[287:0] : _GEN_9412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10463 = 10'h1e5 == _T_25 ? _ram_T_259[287:0] : _GEN_9413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10464 = 10'h1e6 == _T_25 ? _ram_T_259[287:0] : _GEN_9414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10465 = 10'h1e7 == _T_25 ? _ram_T_259[287:0] : _GEN_9415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10466 = 10'h1e8 == _T_25 ? _ram_T_259[287:0] : _GEN_9416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10467 = 10'h1e9 == _T_25 ? _ram_T_259[287:0] : _GEN_9417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10468 = 10'h1ea == _T_25 ? _ram_T_259[287:0] : _GEN_9418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10469 = 10'h1eb == _T_25 ? _ram_T_259[287:0] : _GEN_9419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10470 = 10'h1ec == _T_25 ? _ram_T_259[287:0] : _GEN_9420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10471 = 10'h1ed == _T_25 ? _ram_T_259[287:0] : _GEN_9421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10472 = 10'h1ee == _T_25 ? _ram_T_259[287:0] : _GEN_9422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10473 = 10'h1ef == _T_25 ? _ram_T_259[287:0] : _GEN_9423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10474 = 10'h1f0 == _T_25 ? _ram_T_259[287:0] : _GEN_9424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10475 = 10'h1f1 == _T_25 ? _ram_T_259[287:0] : _GEN_9425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10476 = 10'h1f2 == _T_25 ? _ram_T_259[287:0] : _GEN_9426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10477 = 10'h1f3 == _T_25 ? _ram_T_259[287:0] : _GEN_9427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10478 = 10'h1f4 == _T_25 ? _ram_T_259[287:0] : _GEN_9428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10479 = 10'h1f5 == _T_25 ? _ram_T_259[287:0] : _GEN_9429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10480 = 10'h1f6 == _T_25 ? _ram_T_259[287:0] : _GEN_9430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10481 = 10'h1f7 == _T_25 ? _ram_T_259[287:0] : _GEN_9431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10482 = 10'h1f8 == _T_25 ? _ram_T_259[287:0] : _GEN_9432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10483 = 10'h1f9 == _T_25 ? _ram_T_259[287:0] : _GEN_9433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10484 = 10'h1fa == _T_25 ? _ram_T_259[287:0] : _GEN_9434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10485 = 10'h1fb == _T_25 ? _ram_T_259[287:0] : _GEN_9435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10486 = 10'h1fc == _T_25 ? _ram_T_259[287:0] : _GEN_9436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10487 = 10'h1fd == _T_25 ? _ram_T_259[287:0] : _GEN_9437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10488 = 10'h1fe == _T_25 ? _ram_T_259[287:0] : _GEN_9438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10489 = 10'h1ff == _T_25 ? _ram_T_259[287:0] : _GEN_9439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10490 = 10'h200 == _T_25 ? _ram_T_259[287:0] : _GEN_9440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10491 = 10'h201 == _T_25 ? _ram_T_259[287:0] : _GEN_9441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10492 = 10'h202 == _T_25 ? _ram_T_259[287:0] : _GEN_9442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10493 = 10'h203 == _T_25 ? _ram_T_259[287:0] : _GEN_9443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10494 = 10'h204 == _T_25 ? _ram_T_259[287:0] : _GEN_9444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10495 = 10'h205 == _T_25 ? _ram_T_259[287:0] : _GEN_9445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10496 = 10'h206 == _T_25 ? _ram_T_259[287:0] : _GEN_9446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10497 = 10'h207 == _T_25 ? _ram_T_259[287:0] : _GEN_9447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10498 = 10'h208 == _T_25 ? _ram_T_259[287:0] : _GEN_9448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10499 = 10'h209 == _T_25 ? _ram_T_259[287:0] : _GEN_9449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10500 = 10'h20a == _T_25 ? _ram_T_259[287:0] : _GEN_9450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10501 = 10'h20b == _T_25 ? _ram_T_259[287:0] : _GEN_9451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_10502 = 10'h20c == _T_25 ? _ram_T_259[287:0] : _GEN_9452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_27 = h + 10'ha; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_10 = vga_mem_ram_MPORT_90_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_10 = vga_mem_ram_MPORT_91_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_10 = vga_mem_ram_MPORT_92_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_10 = vga_mem_ram_MPORT_93_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_10 = vga_mem_ram_MPORT_94_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_10 = vga_mem_ram_MPORT_95_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_10 = vga_mem_ram_MPORT_96_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_10 = vga_mem_ram_MPORT_97_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_10 = vga_mem_ram_MPORT_98_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_280 = {278'h0,ram_hi_hi_hi_lo_10,ram_hi_hi_lo_10,ram_hi_lo_hi_10,ram_hi_lo_lo_10,
    ram_lo_hi_hi_hi_10,ram_lo_hi_hi_lo_10,ram_lo_hi_lo_10,ram_lo_lo_hi_10,ram_lo_lo_lo_10}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19080 = {{8191'd0}, _ram_T_280}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_284 = _GEN_19080 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_10504 = 10'h1 == _T_27 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10505 = 10'h2 == _T_27 ? ram_2 : _GEN_10504; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10506 = 10'h3 == _T_27 ? ram_3 : _GEN_10505; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10507 = 10'h4 == _T_27 ? ram_4 : _GEN_10506; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10508 = 10'h5 == _T_27 ? ram_5 : _GEN_10507; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10509 = 10'h6 == _T_27 ? ram_6 : _GEN_10508; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10510 = 10'h7 == _T_27 ? ram_7 : _GEN_10509; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10511 = 10'h8 == _T_27 ? ram_8 : _GEN_10510; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10512 = 10'h9 == _T_27 ? ram_9 : _GEN_10511; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10513 = 10'ha == _T_27 ? ram_10 : _GEN_10512; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10514 = 10'hb == _T_27 ? ram_11 : _GEN_10513; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10515 = 10'hc == _T_27 ? ram_12 : _GEN_10514; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10516 = 10'hd == _T_27 ? ram_13 : _GEN_10515; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10517 = 10'he == _T_27 ? ram_14 : _GEN_10516; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10518 = 10'hf == _T_27 ? ram_15 : _GEN_10517; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10519 = 10'h10 == _T_27 ? ram_16 : _GEN_10518; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10520 = 10'h11 == _T_27 ? ram_17 : _GEN_10519; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10521 = 10'h12 == _T_27 ? ram_18 : _GEN_10520; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10522 = 10'h13 == _T_27 ? ram_19 : _GEN_10521; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10523 = 10'h14 == _T_27 ? ram_20 : _GEN_10522; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10524 = 10'h15 == _T_27 ? ram_21 : _GEN_10523; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10525 = 10'h16 == _T_27 ? ram_22 : _GEN_10524; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10526 = 10'h17 == _T_27 ? ram_23 : _GEN_10525; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10527 = 10'h18 == _T_27 ? ram_24 : _GEN_10526; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10528 = 10'h19 == _T_27 ? ram_25 : _GEN_10527; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10529 = 10'h1a == _T_27 ? ram_26 : _GEN_10528; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10530 = 10'h1b == _T_27 ? ram_27 : _GEN_10529; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10531 = 10'h1c == _T_27 ? ram_28 : _GEN_10530; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10532 = 10'h1d == _T_27 ? ram_29 : _GEN_10531; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10533 = 10'h1e == _T_27 ? ram_30 : _GEN_10532; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10534 = 10'h1f == _T_27 ? ram_31 : _GEN_10533; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10535 = 10'h20 == _T_27 ? ram_32 : _GEN_10534; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10536 = 10'h21 == _T_27 ? ram_33 : _GEN_10535; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10537 = 10'h22 == _T_27 ? ram_34 : _GEN_10536; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10538 = 10'h23 == _T_27 ? ram_35 : _GEN_10537; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10539 = 10'h24 == _T_27 ? ram_36 : _GEN_10538; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10540 = 10'h25 == _T_27 ? ram_37 : _GEN_10539; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10541 = 10'h26 == _T_27 ? ram_38 : _GEN_10540; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10542 = 10'h27 == _T_27 ? ram_39 : _GEN_10541; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10543 = 10'h28 == _T_27 ? ram_40 : _GEN_10542; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10544 = 10'h29 == _T_27 ? ram_41 : _GEN_10543; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10545 = 10'h2a == _T_27 ? ram_42 : _GEN_10544; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10546 = 10'h2b == _T_27 ? ram_43 : _GEN_10545; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10547 = 10'h2c == _T_27 ? ram_44 : _GEN_10546; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10548 = 10'h2d == _T_27 ? ram_45 : _GEN_10547; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10549 = 10'h2e == _T_27 ? ram_46 : _GEN_10548; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10550 = 10'h2f == _T_27 ? ram_47 : _GEN_10549; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10551 = 10'h30 == _T_27 ? ram_48 : _GEN_10550; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10552 = 10'h31 == _T_27 ? ram_49 : _GEN_10551; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10553 = 10'h32 == _T_27 ? ram_50 : _GEN_10552; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10554 = 10'h33 == _T_27 ? ram_51 : _GEN_10553; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10555 = 10'h34 == _T_27 ? ram_52 : _GEN_10554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10556 = 10'h35 == _T_27 ? ram_53 : _GEN_10555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10557 = 10'h36 == _T_27 ? ram_54 : _GEN_10556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10558 = 10'h37 == _T_27 ? ram_55 : _GEN_10557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10559 = 10'h38 == _T_27 ? ram_56 : _GEN_10558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10560 = 10'h39 == _T_27 ? ram_57 : _GEN_10559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10561 = 10'h3a == _T_27 ? ram_58 : _GEN_10560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10562 = 10'h3b == _T_27 ? ram_59 : _GEN_10561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10563 = 10'h3c == _T_27 ? ram_60 : _GEN_10562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10564 = 10'h3d == _T_27 ? ram_61 : _GEN_10563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10565 = 10'h3e == _T_27 ? ram_62 : _GEN_10564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10566 = 10'h3f == _T_27 ? ram_63 : _GEN_10565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10567 = 10'h40 == _T_27 ? ram_64 : _GEN_10566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10568 = 10'h41 == _T_27 ? ram_65 : _GEN_10567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10569 = 10'h42 == _T_27 ? ram_66 : _GEN_10568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10570 = 10'h43 == _T_27 ? ram_67 : _GEN_10569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10571 = 10'h44 == _T_27 ? ram_68 : _GEN_10570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10572 = 10'h45 == _T_27 ? ram_69 : _GEN_10571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10573 = 10'h46 == _T_27 ? ram_70 : _GEN_10572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10574 = 10'h47 == _T_27 ? ram_71 : _GEN_10573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10575 = 10'h48 == _T_27 ? ram_72 : _GEN_10574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10576 = 10'h49 == _T_27 ? ram_73 : _GEN_10575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10577 = 10'h4a == _T_27 ? ram_74 : _GEN_10576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10578 = 10'h4b == _T_27 ? ram_75 : _GEN_10577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10579 = 10'h4c == _T_27 ? ram_76 : _GEN_10578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10580 = 10'h4d == _T_27 ? ram_77 : _GEN_10579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10581 = 10'h4e == _T_27 ? ram_78 : _GEN_10580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10582 = 10'h4f == _T_27 ? ram_79 : _GEN_10581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10583 = 10'h50 == _T_27 ? ram_80 : _GEN_10582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10584 = 10'h51 == _T_27 ? ram_81 : _GEN_10583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10585 = 10'h52 == _T_27 ? ram_82 : _GEN_10584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10586 = 10'h53 == _T_27 ? ram_83 : _GEN_10585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10587 = 10'h54 == _T_27 ? ram_84 : _GEN_10586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10588 = 10'h55 == _T_27 ? ram_85 : _GEN_10587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10589 = 10'h56 == _T_27 ? ram_86 : _GEN_10588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10590 = 10'h57 == _T_27 ? ram_87 : _GEN_10589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10591 = 10'h58 == _T_27 ? ram_88 : _GEN_10590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10592 = 10'h59 == _T_27 ? ram_89 : _GEN_10591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10593 = 10'h5a == _T_27 ? ram_90 : _GEN_10592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10594 = 10'h5b == _T_27 ? ram_91 : _GEN_10593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10595 = 10'h5c == _T_27 ? ram_92 : _GEN_10594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10596 = 10'h5d == _T_27 ? ram_93 : _GEN_10595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10597 = 10'h5e == _T_27 ? ram_94 : _GEN_10596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10598 = 10'h5f == _T_27 ? ram_95 : _GEN_10597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10599 = 10'h60 == _T_27 ? ram_96 : _GEN_10598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10600 = 10'h61 == _T_27 ? ram_97 : _GEN_10599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10601 = 10'h62 == _T_27 ? ram_98 : _GEN_10600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10602 = 10'h63 == _T_27 ? ram_99 : _GEN_10601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10603 = 10'h64 == _T_27 ? ram_100 : _GEN_10602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10604 = 10'h65 == _T_27 ? ram_101 : _GEN_10603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10605 = 10'h66 == _T_27 ? ram_102 : _GEN_10604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10606 = 10'h67 == _T_27 ? ram_103 : _GEN_10605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10607 = 10'h68 == _T_27 ? ram_104 : _GEN_10606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10608 = 10'h69 == _T_27 ? ram_105 : _GEN_10607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10609 = 10'h6a == _T_27 ? ram_106 : _GEN_10608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10610 = 10'h6b == _T_27 ? ram_107 : _GEN_10609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10611 = 10'h6c == _T_27 ? ram_108 : _GEN_10610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10612 = 10'h6d == _T_27 ? ram_109 : _GEN_10611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10613 = 10'h6e == _T_27 ? ram_110 : _GEN_10612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10614 = 10'h6f == _T_27 ? ram_111 : _GEN_10613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10615 = 10'h70 == _T_27 ? ram_112 : _GEN_10614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10616 = 10'h71 == _T_27 ? ram_113 : _GEN_10615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10617 = 10'h72 == _T_27 ? ram_114 : _GEN_10616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10618 = 10'h73 == _T_27 ? ram_115 : _GEN_10617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10619 = 10'h74 == _T_27 ? ram_116 : _GEN_10618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10620 = 10'h75 == _T_27 ? ram_117 : _GEN_10619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10621 = 10'h76 == _T_27 ? ram_118 : _GEN_10620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10622 = 10'h77 == _T_27 ? ram_119 : _GEN_10621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10623 = 10'h78 == _T_27 ? ram_120 : _GEN_10622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10624 = 10'h79 == _T_27 ? ram_121 : _GEN_10623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10625 = 10'h7a == _T_27 ? ram_122 : _GEN_10624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10626 = 10'h7b == _T_27 ? ram_123 : _GEN_10625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10627 = 10'h7c == _T_27 ? ram_124 : _GEN_10626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10628 = 10'h7d == _T_27 ? ram_125 : _GEN_10627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10629 = 10'h7e == _T_27 ? ram_126 : _GEN_10628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10630 = 10'h7f == _T_27 ? ram_127 : _GEN_10629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10631 = 10'h80 == _T_27 ? ram_128 : _GEN_10630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10632 = 10'h81 == _T_27 ? ram_129 : _GEN_10631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10633 = 10'h82 == _T_27 ? ram_130 : _GEN_10632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10634 = 10'h83 == _T_27 ? ram_131 : _GEN_10633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10635 = 10'h84 == _T_27 ? ram_132 : _GEN_10634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10636 = 10'h85 == _T_27 ? ram_133 : _GEN_10635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10637 = 10'h86 == _T_27 ? ram_134 : _GEN_10636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10638 = 10'h87 == _T_27 ? ram_135 : _GEN_10637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10639 = 10'h88 == _T_27 ? ram_136 : _GEN_10638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10640 = 10'h89 == _T_27 ? ram_137 : _GEN_10639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10641 = 10'h8a == _T_27 ? ram_138 : _GEN_10640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10642 = 10'h8b == _T_27 ? ram_139 : _GEN_10641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10643 = 10'h8c == _T_27 ? ram_140 : _GEN_10642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10644 = 10'h8d == _T_27 ? ram_141 : _GEN_10643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10645 = 10'h8e == _T_27 ? ram_142 : _GEN_10644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10646 = 10'h8f == _T_27 ? ram_143 : _GEN_10645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10647 = 10'h90 == _T_27 ? ram_144 : _GEN_10646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10648 = 10'h91 == _T_27 ? ram_145 : _GEN_10647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10649 = 10'h92 == _T_27 ? ram_146 : _GEN_10648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10650 = 10'h93 == _T_27 ? ram_147 : _GEN_10649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10651 = 10'h94 == _T_27 ? ram_148 : _GEN_10650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10652 = 10'h95 == _T_27 ? ram_149 : _GEN_10651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10653 = 10'h96 == _T_27 ? ram_150 : _GEN_10652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10654 = 10'h97 == _T_27 ? ram_151 : _GEN_10653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10655 = 10'h98 == _T_27 ? ram_152 : _GEN_10654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10656 = 10'h99 == _T_27 ? ram_153 : _GEN_10655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10657 = 10'h9a == _T_27 ? ram_154 : _GEN_10656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10658 = 10'h9b == _T_27 ? ram_155 : _GEN_10657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10659 = 10'h9c == _T_27 ? ram_156 : _GEN_10658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10660 = 10'h9d == _T_27 ? ram_157 : _GEN_10659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10661 = 10'h9e == _T_27 ? ram_158 : _GEN_10660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10662 = 10'h9f == _T_27 ? ram_159 : _GEN_10661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10663 = 10'ha0 == _T_27 ? ram_160 : _GEN_10662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10664 = 10'ha1 == _T_27 ? ram_161 : _GEN_10663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10665 = 10'ha2 == _T_27 ? ram_162 : _GEN_10664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10666 = 10'ha3 == _T_27 ? ram_163 : _GEN_10665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10667 = 10'ha4 == _T_27 ? ram_164 : _GEN_10666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10668 = 10'ha5 == _T_27 ? ram_165 : _GEN_10667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10669 = 10'ha6 == _T_27 ? ram_166 : _GEN_10668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10670 = 10'ha7 == _T_27 ? ram_167 : _GEN_10669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10671 = 10'ha8 == _T_27 ? ram_168 : _GEN_10670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10672 = 10'ha9 == _T_27 ? ram_169 : _GEN_10671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10673 = 10'haa == _T_27 ? ram_170 : _GEN_10672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10674 = 10'hab == _T_27 ? ram_171 : _GEN_10673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10675 = 10'hac == _T_27 ? ram_172 : _GEN_10674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10676 = 10'had == _T_27 ? ram_173 : _GEN_10675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10677 = 10'hae == _T_27 ? ram_174 : _GEN_10676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10678 = 10'haf == _T_27 ? ram_175 : _GEN_10677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10679 = 10'hb0 == _T_27 ? ram_176 : _GEN_10678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10680 = 10'hb1 == _T_27 ? ram_177 : _GEN_10679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10681 = 10'hb2 == _T_27 ? ram_178 : _GEN_10680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10682 = 10'hb3 == _T_27 ? ram_179 : _GEN_10681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10683 = 10'hb4 == _T_27 ? ram_180 : _GEN_10682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10684 = 10'hb5 == _T_27 ? ram_181 : _GEN_10683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10685 = 10'hb6 == _T_27 ? ram_182 : _GEN_10684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10686 = 10'hb7 == _T_27 ? ram_183 : _GEN_10685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10687 = 10'hb8 == _T_27 ? ram_184 : _GEN_10686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10688 = 10'hb9 == _T_27 ? ram_185 : _GEN_10687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10689 = 10'hba == _T_27 ? ram_186 : _GEN_10688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10690 = 10'hbb == _T_27 ? ram_187 : _GEN_10689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10691 = 10'hbc == _T_27 ? ram_188 : _GEN_10690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10692 = 10'hbd == _T_27 ? ram_189 : _GEN_10691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10693 = 10'hbe == _T_27 ? ram_190 : _GEN_10692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10694 = 10'hbf == _T_27 ? ram_191 : _GEN_10693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10695 = 10'hc0 == _T_27 ? ram_192 : _GEN_10694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10696 = 10'hc1 == _T_27 ? ram_193 : _GEN_10695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10697 = 10'hc2 == _T_27 ? ram_194 : _GEN_10696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10698 = 10'hc3 == _T_27 ? ram_195 : _GEN_10697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10699 = 10'hc4 == _T_27 ? ram_196 : _GEN_10698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10700 = 10'hc5 == _T_27 ? ram_197 : _GEN_10699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10701 = 10'hc6 == _T_27 ? ram_198 : _GEN_10700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10702 = 10'hc7 == _T_27 ? ram_199 : _GEN_10701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10703 = 10'hc8 == _T_27 ? ram_200 : _GEN_10702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10704 = 10'hc9 == _T_27 ? ram_201 : _GEN_10703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10705 = 10'hca == _T_27 ? ram_202 : _GEN_10704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10706 = 10'hcb == _T_27 ? ram_203 : _GEN_10705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10707 = 10'hcc == _T_27 ? ram_204 : _GEN_10706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10708 = 10'hcd == _T_27 ? ram_205 : _GEN_10707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10709 = 10'hce == _T_27 ? ram_206 : _GEN_10708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10710 = 10'hcf == _T_27 ? ram_207 : _GEN_10709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10711 = 10'hd0 == _T_27 ? ram_208 : _GEN_10710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10712 = 10'hd1 == _T_27 ? ram_209 : _GEN_10711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10713 = 10'hd2 == _T_27 ? ram_210 : _GEN_10712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10714 = 10'hd3 == _T_27 ? ram_211 : _GEN_10713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10715 = 10'hd4 == _T_27 ? ram_212 : _GEN_10714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10716 = 10'hd5 == _T_27 ? ram_213 : _GEN_10715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10717 = 10'hd6 == _T_27 ? ram_214 : _GEN_10716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10718 = 10'hd7 == _T_27 ? ram_215 : _GEN_10717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10719 = 10'hd8 == _T_27 ? ram_216 : _GEN_10718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10720 = 10'hd9 == _T_27 ? ram_217 : _GEN_10719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10721 = 10'hda == _T_27 ? ram_218 : _GEN_10720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10722 = 10'hdb == _T_27 ? ram_219 : _GEN_10721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10723 = 10'hdc == _T_27 ? ram_220 : _GEN_10722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10724 = 10'hdd == _T_27 ? ram_221 : _GEN_10723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10725 = 10'hde == _T_27 ? ram_222 : _GEN_10724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10726 = 10'hdf == _T_27 ? ram_223 : _GEN_10725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10727 = 10'he0 == _T_27 ? ram_224 : _GEN_10726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10728 = 10'he1 == _T_27 ? ram_225 : _GEN_10727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10729 = 10'he2 == _T_27 ? ram_226 : _GEN_10728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10730 = 10'he3 == _T_27 ? ram_227 : _GEN_10729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10731 = 10'he4 == _T_27 ? ram_228 : _GEN_10730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10732 = 10'he5 == _T_27 ? ram_229 : _GEN_10731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10733 = 10'he6 == _T_27 ? ram_230 : _GEN_10732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10734 = 10'he7 == _T_27 ? ram_231 : _GEN_10733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10735 = 10'he8 == _T_27 ? ram_232 : _GEN_10734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10736 = 10'he9 == _T_27 ? ram_233 : _GEN_10735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10737 = 10'hea == _T_27 ? ram_234 : _GEN_10736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10738 = 10'heb == _T_27 ? ram_235 : _GEN_10737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10739 = 10'hec == _T_27 ? ram_236 : _GEN_10738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10740 = 10'hed == _T_27 ? ram_237 : _GEN_10739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10741 = 10'hee == _T_27 ? ram_238 : _GEN_10740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10742 = 10'hef == _T_27 ? ram_239 : _GEN_10741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10743 = 10'hf0 == _T_27 ? ram_240 : _GEN_10742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10744 = 10'hf1 == _T_27 ? ram_241 : _GEN_10743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10745 = 10'hf2 == _T_27 ? ram_242 : _GEN_10744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10746 = 10'hf3 == _T_27 ? ram_243 : _GEN_10745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10747 = 10'hf4 == _T_27 ? ram_244 : _GEN_10746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10748 = 10'hf5 == _T_27 ? ram_245 : _GEN_10747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10749 = 10'hf6 == _T_27 ? ram_246 : _GEN_10748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10750 = 10'hf7 == _T_27 ? ram_247 : _GEN_10749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10751 = 10'hf8 == _T_27 ? ram_248 : _GEN_10750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10752 = 10'hf9 == _T_27 ? ram_249 : _GEN_10751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10753 = 10'hfa == _T_27 ? ram_250 : _GEN_10752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10754 = 10'hfb == _T_27 ? ram_251 : _GEN_10753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10755 = 10'hfc == _T_27 ? ram_252 : _GEN_10754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10756 = 10'hfd == _T_27 ? ram_253 : _GEN_10755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10757 = 10'hfe == _T_27 ? ram_254 : _GEN_10756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10758 = 10'hff == _T_27 ? ram_255 : _GEN_10757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10759 = 10'h100 == _T_27 ? ram_256 : _GEN_10758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10760 = 10'h101 == _T_27 ? ram_257 : _GEN_10759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10761 = 10'h102 == _T_27 ? ram_258 : _GEN_10760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10762 = 10'h103 == _T_27 ? ram_259 : _GEN_10761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10763 = 10'h104 == _T_27 ? ram_260 : _GEN_10762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10764 = 10'h105 == _T_27 ? ram_261 : _GEN_10763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10765 = 10'h106 == _T_27 ? ram_262 : _GEN_10764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10766 = 10'h107 == _T_27 ? ram_263 : _GEN_10765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10767 = 10'h108 == _T_27 ? ram_264 : _GEN_10766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10768 = 10'h109 == _T_27 ? ram_265 : _GEN_10767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10769 = 10'h10a == _T_27 ? ram_266 : _GEN_10768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10770 = 10'h10b == _T_27 ? ram_267 : _GEN_10769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10771 = 10'h10c == _T_27 ? ram_268 : _GEN_10770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10772 = 10'h10d == _T_27 ? ram_269 : _GEN_10771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10773 = 10'h10e == _T_27 ? ram_270 : _GEN_10772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10774 = 10'h10f == _T_27 ? ram_271 : _GEN_10773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10775 = 10'h110 == _T_27 ? ram_272 : _GEN_10774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10776 = 10'h111 == _T_27 ? ram_273 : _GEN_10775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10777 = 10'h112 == _T_27 ? ram_274 : _GEN_10776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10778 = 10'h113 == _T_27 ? ram_275 : _GEN_10777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10779 = 10'h114 == _T_27 ? ram_276 : _GEN_10778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10780 = 10'h115 == _T_27 ? ram_277 : _GEN_10779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10781 = 10'h116 == _T_27 ? ram_278 : _GEN_10780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10782 = 10'h117 == _T_27 ? ram_279 : _GEN_10781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10783 = 10'h118 == _T_27 ? ram_280 : _GEN_10782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10784 = 10'h119 == _T_27 ? ram_281 : _GEN_10783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10785 = 10'h11a == _T_27 ? ram_282 : _GEN_10784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10786 = 10'h11b == _T_27 ? ram_283 : _GEN_10785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10787 = 10'h11c == _T_27 ? ram_284 : _GEN_10786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10788 = 10'h11d == _T_27 ? ram_285 : _GEN_10787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10789 = 10'h11e == _T_27 ? ram_286 : _GEN_10788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10790 = 10'h11f == _T_27 ? ram_287 : _GEN_10789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10791 = 10'h120 == _T_27 ? ram_288 : _GEN_10790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10792 = 10'h121 == _T_27 ? ram_289 : _GEN_10791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10793 = 10'h122 == _T_27 ? ram_290 : _GEN_10792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10794 = 10'h123 == _T_27 ? ram_291 : _GEN_10793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10795 = 10'h124 == _T_27 ? ram_292 : _GEN_10794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10796 = 10'h125 == _T_27 ? ram_293 : _GEN_10795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10797 = 10'h126 == _T_27 ? ram_294 : _GEN_10796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10798 = 10'h127 == _T_27 ? ram_295 : _GEN_10797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10799 = 10'h128 == _T_27 ? ram_296 : _GEN_10798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10800 = 10'h129 == _T_27 ? ram_297 : _GEN_10799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10801 = 10'h12a == _T_27 ? ram_298 : _GEN_10800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10802 = 10'h12b == _T_27 ? ram_299 : _GEN_10801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10803 = 10'h12c == _T_27 ? ram_300 : _GEN_10802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10804 = 10'h12d == _T_27 ? ram_301 : _GEN_10803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10805 = 10'h12e == _T_27 ? ram_302 : _GEN_10804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10806 = 10'h12f == _T_27 ? ram_303 : _GEN_10805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10807 = 10'h130 == _T_27 ? ram_304 : _GEN_10806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10808 = 10'h131 == _T_27 ? ram_305 : _GEN_10807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10809 = 10'h132 == _T_27 ? ram_306 : _GEN_10808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10810 = 10'h133 == _T_27 ? ram_307 : _GEN_10809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10811 = 10'h134 == _T_27 ? ram_308 : _GEN_10810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10812 = 10'h135 == _T_27 ? ram_309 : _GEN_10811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10813 = 10'h136 == _T_27 ? ram_310 : _GEN_10812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10814 = 10'h137 == _T_27 ? ram_311 : _GEN_10813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10815 = 10'h138 == _T_27 ? ram_312 : _GEN_10814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10816 = 10'h139 == _T_27 ? ram_313 : _GEN_10815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10817 = 10'h13a == _T_27 ? ram_314 : _GEN_10816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10818 = 10'h13b == _T_27 ? ram_315 : _GEN_10817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10819 = 10'h13c == _T_27 ? ram_316 : _GEN_10818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10820 = 10'h13d == _T_27 ? ram_317 : _GEN_10819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10821 = 10'h13e == _T_27 ? ram_318 : _GEN_10820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10822 = 10'h13f == _T_27 ? ram_319 : _GEN_10821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10823 = 10'h140 == _T_27 ? ram_320 : _GEN_10822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10824 = 10'h141 == _T_27 ? ram_321 : _GEN_10823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10825 = 10'h142 == _T_27 ? ram_322 : _GEN_10824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10826 = 10'h143 == _T_27 ? ram_323 : _GEN_10825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10827 = 10'h144 == _T_27 ? ram_324 : _GEN_10826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10828 = 10'h145 == _T_27 ? ram_325 : _GEN_10827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10829 = 10'h146 == _T_27 ? ram_326 : _GEN_10828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10830 = 10'h147 == _T_27 ? ram_327 : _GEN_10829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10831 = 10'h148 == _T_27 ? ram_328 : _GEN_10830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10832 = 10'h149 == _T_27 ? ram_329 : _GEN_10831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10833 = 10'h14a == _T_27 ? ram_330 : _GEN_10832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10834 = 10'h14b == _T_27 ? ram_331 : _GEN_10833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10835 = 10'h14c == _T_27 ? ram_332 : _GEN_10834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10836 = 10'h14d == _T_27 ? ram_333 : _GEN_10835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10837 = 10'h14e == _T_27 ? ram_334 : _GEN_10836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10838 = 10'h14f == _T_27 ? ram_335 : _GEN_10837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10839 = 10'h150 == _T_27 ? ram_336 : _GEN_10838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10840 = 10'h151 == _T_27 ? ram_337 : _GEN_10839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10841 = 10'h152 == _T_27 ? ram_338 : _GEN_10840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10842 = 10'h153 == _T_27 ? ram_339 : _GEN_10841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10843 = 10'h154 == _T_27 ? ram_340 : _GEN_10842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10844 = 10'h155 == _T_27 ? ram_341 : _GEN_10843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10845 = 10'h156 == _T_27 ? ram_342 : _GEN_10844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10846 = 10'h157 == _T_27 ? ram_343 : _GEN_10845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10847 = 10'h158 == _T_27 ? ram_344 : _GEN_10846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10848 = 10'h159 == _T_27 ? ram_345 : _GEN_10847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10849 = 10'h15a == _T_27 ? ram_346 : _GEN_10848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10850 = 10'h15b == _T_27 ? ram_347 : _GEN_10849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10851 = 10'h15c == _T_27 ? ram_348 : _GEN_10850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10852 = 10'h15d == _T_27 ? ram_349 : _GEN_10851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10853 = 10'h15e == _T_27 ? ram_350 : _GEN_10852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10854 = 10'h15f == _T_27 ? ram_351 : _GEN_10853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10855 = 10'h160 == _T_27 ? ram_352 : _GEN_10854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10856 = 10'h161 == _T_27 ? ram_353 : _GEN_10855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10857 = 10'h162 == _T_27 ? ram_354 : _GEN_10856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10858 = 10'h163 == _T_27 ? ram_355 : _GEN_10857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10859 = 10'h164 == _T_27 ? ram_356 : _GEN_10858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10860 = 10'h165 == _T_27 ? ram_357 : _GEN_10859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10861 = 10'h166 == _T_27 ? ram_358 : _GEN_10860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10862 = 10'h167 == _T_27 ? ram_359 : _GEN_10861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10863 = 10'h168 == _T_27 ? ram_360 : _GEN_10862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10864 = 10'h169 == _T_27 ? ram_361 : _GEN_10863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10865 = 10'h16a == _T_27 ? ram_362 : _GEN_10864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10866 = 10'h16b == _T_27 ? ram_363 : _GEN_10865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10867 = 10'h16c == _T_27 ? ram_364 : _GEN_10866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10868 = 10'h16d == _T_27 ? ram_365 : _GEN_10867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10869 = 10'h16e == _T_27 ? ram_366 : _GEN_10868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10870 = 10'h16f == _T_27 ? ram_367 : _GEN_10869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10871 = 10'h170 == _T_27 ? ram_368 : _GEN_10870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10872 = 10'h171 == _T_27 ? ram_369 : _GEN_10871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10873 = 10'h172 == _T_27 ? ram_370 : _GEN_10872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10874 = 10'h173 == _T_27 ? ram_371 : _GEN_10873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10875 = 10'h174 == _T_27 ? ram_372 : _GEN_10874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10876 = 10'h175 == _T_27 ? ram_373 : _GEN_10875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10877 = 10'h176 == _T_27 ? ram_374 : _GEN_10876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10878 = 10'h177 == _T_27 ? ram_375 : _GEN_10877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10879 = 10'h178 == _T_27 ? ram_376 : _GEN_10878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10880 = 10'h179 == _T_27 ? ram_377 : _GEN_10879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10881 = 10'h17a == _T_27 ? ram_378 : _GEN_10880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10882 = 10'h17b == _T_27 ? ram_379 : _GEN_10881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10883 = 10'h17c == _T_27 ? ram_380 : _GEN_10882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10884 = 10'h17d == _T_27 ? ram_381 : _GEN_10883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10885 = 10'h17e == _T_27 ? ram_382 : _GEN_10884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10886 = 10'h17f == _T_27 ? ram_383 : _GEN_10885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10887 = 10'h180 == _T_27 ? ram_384 : _GEN_10886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10888 = 10'h181 == _T_27 ? ram_385 : _GEN_10887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10889 = 10'h182 == _T_27 ? ram_386 : _GEN_10888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10890 = 10'h183 == _T_27 ? ram_387 : _GEN_10889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10891 = 10'h184 == _T_27 ? ram_388 : _GEN_10890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10892 = 10'h185 == _T_27 ? ram_389 : _GEN_10891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10893 = 10'h186 == _T_27 ? ram_390 : _GEN_10892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10894 = 10'h187 == _T_27 ? ram_391 : _GEN_10893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10895 = 10'h188 == _T_27 ? ram_392 : _GEN_10894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10896 = 10'h189 == _T_27 ? ram_393 : _GEN_10895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10897 = 10'h18a == _T_27 ? ram_394 : _GEN_10896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10898 = 10'h18b == _T_27 ? ram_395 : _GEN_10897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10899 = 10'h18c == _T_27 ? ram_396 : _GEN_10898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10900 = 10'h18d == _T_27 ? ram_397 : _GEN_10899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10901 = 10'h18e == _T_27 ? ram_398 : _GEN_10900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10902 = 10'h18f == _T_27 ? ram_399 : _GEN_10901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10903 = 10'h190 == _T_27 ? ram_400 : _GEN_10902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10904 = 10'h191 == _T_27 ? ram_401 : _GEN_10903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10905 = 10'h192 == _T_27 ? ram_402 : _GEN_10904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10906 = 10'h193 == _T_27 ? ram_403 : _GEN_10905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10907 = 10'h194 == _T_27 ? ram_404 : _GEN_10906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10908 = 10'h195 == _T_27 ? ram_405 : _GEN_10907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10909 = 10'h196 == _T_27 ? ram_406 : _GEN_10908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10910 = 10'h197 == _T_27 ? ram_407 : _GEN_10909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10911 = 10'h198 == _T_27 ? ram_408 : _GEN_10910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10912 = 10'h199 == _T_27 ? ram_409 : _GEN_10911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10913 = 10'h19a == _T_27 ? ram_410 : _GEN_10912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10914 = 10'h19b == _T_27 ? ram_411 : _GEN_10913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10915 = 10'h19c == _T_27 ? ram_412 : _GEN_10914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10916 = 10'h19d == _T_27 ? ram_413 : _GEN_10915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10917 = 10'h19e == _T_27 ? ram_414 : _GEN_10916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10918 = 10'h19f == _T_27 ? ram_415 : _GEN_10917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10919 = 10'h1a0 == _T_27 ? ram_416 : _GEN_10918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10920 = 10'h1a1 == _T_27 ? ram_417 : _GEN_10919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10921 = 10'h1a2 == _T_27 ? ram_418 : _GEN_10920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10922 = 10'h1a3 == _T_27 ? ram_419 : _GEN_10921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10923 = 10'h1a4 == _T_27 ? ram_420 : _GEN_10922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10924 = 10'h1a5 == _T_27 ? ram_421 : _GEN_10923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10925 = 10'h1a6 == _T_27 ? ram_422 : _GEN_10924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10926 = 10'h1a7 == _T_27 ? ram_423 : _GEN_10925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10927 = 10'h1a8 == _T_27 ? ram_424 : _GEN_10926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10928 = 10'h1a9 == _T_27 ? ram_425 : _GEN_10927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10929 = 10'h1aa == _T_27 ? ram_426 : _GEN_10928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10930 = 10'h1ab == _T_27 ? ram_427 : _GEN_10929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10931 = 10'h1ac == _T_27 ? ram_428 : _GEN_10930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10932 = 10'h1ad == _T_27 ? ram_429 : _GEN_10931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10933 = 10'h1ae == _T_27 ? ram_430 : _GEN_10932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10934 = 10'h1af == _T_27 ? ram_431 : _GEN_10933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10935 = 10'h1b0 == _T_27 ? ram_432 : _GEN_10934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10936 = 10'h1b1 == _T_27 ? ram_433 : _GEN_10935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10937 = 10'h1b2 == _T_27 ? ram_434 : _GEN_10936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10938 = 10'h1b3 == _T_27 ? ram_435 : _GEN_10937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10939 = 10'h1b4 == _T_27 ? ram_436 : _GEN_10938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10940 = 10'h1b5 == _T_27 ? ram_437 : _GEN_10939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10941 = 10'h1b6 == _T_27 ? ram_438 : _GEN_10940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10942 = 10'h1b7 == _T_27 ? ram_439 : _GEN_10941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10943 = 10'h1b8 == _T_27 ? ram_440 : _GEN_10942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10944 = 10'h1b9 == _T_27 ? ram_441 : _GEN_10943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10945 = 10'h1ba == _T_27 ? ram_442 : _GEN_10944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10946 = 10'h1bb == _T_27 ? ram_443 : _GEN_10945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10947 = 10'h1bc == _T_27 ? ram_444 : _GEN_10946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10948 = 10'h1bd == _T_27 ? ram_445 : _GEN_10947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10949 = 10'h1be == _T_27 ? ram_446 : _GEN_10948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10950 = 10'h1bf == _T_27 ? ram_447 : _GEN_10949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10951 = 10'h1c0 == _T_27 ? ram_448 : _GEN_10950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10952 = 10'h1c1 == _T_27 ? ram_449 : _GEN_10951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10953 = 10'h1c2 == _T_27 ? ram_450 : _GEN_10952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10954 = 10'h1c3 == _T_27 ? ram_451 : _GEN_10953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10955 = 10'h1c4 == _T_27 ? ram_452 : _GEN_10954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10956 = 10'h1c5 == _T_27 ? ram_453 : _GEN_10955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10957 = 10'h1c6 == _T_27 ? ram_454 : _GEN_10956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10958 = 10'h1c7 == _T_27 ? ram_455 : _GEN_10957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10959 = 10'h1c8 == _T_27 ? ram_456 : _GEN_10958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10960 = 10'h1c9 == _T_27 ? ram_457 : _GEN_10959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10961 = 10'h1ca == _T_27 ? ram_458 : _GEN_10960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10962 = 10'h1cb == _T_27 ? ram_459 : _GEN_10961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10963 = 10'h1cc == _T_27 ? ram_460 : _GEN_10962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10964 = 10'h1cd == _T_27 ? ram_461 : _GEN_10963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10965 = 10'h1ce == _T_27 ? ram_462 : _GEN_10964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10966 = 10'h1cf == _T_27 ? ram_463 : _GEN_10965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10967 = 10'h1d0 == _T_27 ? ram_464 : _GEN_10966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10968 = 10'h1d1 == _T_27 ? ram_465 : _GEN_10967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10969 = 10'h1d2 == _T_27 ? ram_466 : _GEN_10968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10970 = 10'h1d3 == _T_27 ? ram_467 : _GEN_10969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10971 = 10'h1d4 == _T_27 ? ram_468 : _GEN_10970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10972 = 10'h1d5 == _T_27 ? ram_469 : _GEN_10971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10973 = 10'h1d6 == _T_27 ? ram_470 : _GEN_10972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10974 = 10'h1d7 == _T_27 ? ram_471 : _GEN_10973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10975 = 10'h1d8 == _T_27 ? ram_472 : _GEN_10974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10976 = 10'h1d9 == _T_27 ? ram_473 : _GEN_10975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10977 = 10'h1da == _T_27 ? ram_474 : _GEN_10976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10978 = 10'h1db == _T_27 ? ram_475 : _GEN_10977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10979 = 10'h1dc == _T_27 ? ram_476 : _GEN_10978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10980 = 10'h1dd == _T_27 ? ram_477 : _GEN_10979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10981 = 10'h1de == _T_27 ? ram_478 : _GEN_10980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10982 = 10'h1df == _T_27 ? ram_479 : _GEN_10981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10983 = 10'h1e0 == _T_27 ? ram_480 : _GEN_10982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10984 = 10'h1e1 == _T_27 ? ram_481 : _GEN_10983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10985 = 10'h1e2 == _T_27 ? ram_482 : _GEN_10984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10986 = 10'h1e3 == _T_27 ? ram_483 : _GEN_10985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10987 = 10'h1e4 == _T_27 ? ram_484 : _GEN_10986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10988 = 10'h1e5 == _T_27 ? ram_485 : _GEN_10987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10989 = 10'h1e6 == _T_27 ? ram_486 : _GEN_10988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10990 = 10'h1e7 == _T_27 ? ram_487 : _GEN_10989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10991 = 10'h1e8 == _T_27 ? ram_488 : _GEN_10990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10992 = 10'h1e9 == _T_27 ? ram_489 : _GEN_10991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10993 = 10'h1ea == _T_27 ? ram_490 : _GEN_10992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10994 = 10'h1eb == _T_27 ? ram_491 : _GEN_10993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10995 = 10'h1ec == _T_27 ? ram_492 : _GEN_10994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10996 = 10'h1ed == _T_27 ? ram_493 : _GEN_10995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10997 = 10'h1ee == _T_27 ? ram_494 : _GEN_10996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10998 = 10'h1ef == _T_27 ? ram_495 : _GEN_10997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_10999 = 10'h1f0 == _T_27 ? ram_496 : _GEN_10998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11000 = 10'h1f1 == _T_27 ? ram_497 : _GEN_10999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11001 = 10'h1f2 == _T_27 ? ram_498 : _GEN_11000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11002 = 10'h1f3 == _T_27 ? ram_499 : _GEN_11001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11003 = 10'h1f4 == _T_27 ? ram_500 : _GEN_11002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11004 = 10'h1f5 == _T_27 ? ram_501 : _GEN_11003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11005 = 10'h1f6 == _T_27 ? ram_502 : _GEN_11004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11006 = 10'h1f7 == _T_27 ? ram_503 : _GEN_11005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11007 = 10'h1f8 == _T_27 ? ram_504 : _GEN_11006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11008 = 10'h1f9 == _T_27 ? ram_505 : _GEN_11007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11009 = 10'h1fa == _T_27 ? ram_506 : _GEN_11008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11010 = 10'h1fb == _T_27 ? ram_507 : _GEN_11009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11011 = 10'h1fc == _T_27 ? ram_508 : _GEN_11010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11012 = 10'h1fd == _T_27 ? ram_509 : _GEN_11011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11013 = 10'h1fe == _T_27 ? ram_510 : _GEN_11012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11014 = 10'h1ff == _T_27 ? ram_511 : _GEN_11013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11015 = 10'h200 == _T_27 ? ram_512 : _GEN_11014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11016 = 10'h201 == _T_27 ? ram_513 : _GEN_11015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11017 = 10'h202 == _T_27 ? ram_514 : _GEN_11016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11018 = 10'h203 == _T_27 ? ram_515 : _GEN_11017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11019 = 10'h204 == _T_27 ? ram_516 : _GEN_11018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11020 = 10'h205 == _T_27 ? ram_517 : _GEN_11019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11021 = 10'h206 == _T_27 ? ram_518 : _GEN_11020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11022 = 10'h207 == _T_27 ? ram_519 : _GEN_11021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11023 = 10'h208 == _T_27 ? ram_520 : _GEN_11022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11024 = 10'h209 == _T_27 ? ram_521 : _GEN_11023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11025 = 10'h20a == _T_27 ? ram_522 : _GEN_11024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11026 = 10'h20b == _T_27 ? ram_523 : _GEN_11025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11027 = 10'h20c == _T_27 ? ram_524 : _GEN_11026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19081 = {{8190'd0}, _GEN_11027}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_285 = _GEN_19081 ^ _ram_T_284; // @[vga.scala 64:41]
  wire [287:0] _GEN_11028 = 10'h0 == _T_27 ? _ram_T_285[287:0] : _GEN_9978; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11029 = 10'h1 == _T_27 ? _ram_T_285[287:0] : _GEN_9979; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11030 = 10'h2 == _T_27 ? _ram_T_285[287:0] : _GEN_9980; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11031 = 10'h3 == _T_27 ? _ram_T_285[287:0] : _GEN_9981; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11032 = 10'h4 == _T_27 ? _ram_T_285[287:0] : _GEN_9982; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11033 = 10'h5 == _T_27 ? _ram_T_285[287:0] : _GEN_9983; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11034 = 10'h6 == _T_27 ? _ram_T_285[287:0] : _GEN_9984; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11035 = 10'h7 == _T_27 ? _ram_T_285[287:0] : _GEN_9985; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11036 = 10'h8 == _T_27 ? _ram_T_285[287:0] : _GEN_9986; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11037 = 10'h9 == _T_27 ? _ram_T_285[287:0] : _GEN_9987; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11038 = 10'ha == _T_27 ? _ram_T_285[287:0] : _GEN_9988; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11039 = 10'hb == _T_27 ? _ram_T_285[287:0] : _GEN_9989; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11040 = 10'hc == _T_27 ? _ram_T_285[287:0] : _GEN_9990; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11041 = 10'hd == _T_27 ? _ram_T_285[287:0] : _GEN_9991; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11042 = 10'he == _T_27 ? _ram_T_285[287:0] : _GEN_9992; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11043 = 10'hf == _T_27 ? _ram_T_285[287:0] : _GEN_9993; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11044 = 10'h10 == _T_27 ? _ram_T_285[287:0] : _GEN_9994; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11045 = 10'h11 == _T_27 ? _ram_T_285[287:0] : _GEN_9995; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11046 = 10'h12 == _T_27 ? _ram_T_285[287:0] : _GEN_9996; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11047 = 10'h13 == _T_27 ? _ram_T_285[287:0] : _GEN_9997; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11048 = 10'h14 == _T_27 ? _ram_T_285[287:0] : _GEN_9998; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11049 = 10'h15 == _T_27 ? _ram_T_285[287:0] : _GEN_9999; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11050 = 10'h16 == _T_27 ? _ram_T_285[287:0] : _GEN_10000; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11051 = 10'h17 == _T_27 ? _ram_T_285[287:0] : _GEN_10001; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11052 = 10'h18 == _T_27 ? _ram_T_285[287:0] : _GEN_10002; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11053 = 10'h19 == _T_27 ? _ram_T_285[287:0] : _GEN_10003; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11054 = 10'h1a == _T_27 ? _ram_T_285[287:0] : _GEN_10004; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11055 = 10'h1b == _T_27 ? _ram_T_285[287:0] : _GEN_10005; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11056 = 10'h1c == _T_27 ? _ram_T_285[287:0] : _GEN_10006; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11057 = 10'h1d == _T_27 ? _ram_T_285[287:0] : _GEN_10007; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11058 = 10'h1e == _T_27 ? _ram_T_285[287:0] : _GEN_10008; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11059 = 10'h1f == _T_27 ? _ram_T_285[287:0] : _GEN_10009; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11060 = 10'h20 == _T_27 ? _ram_T_285[287:0] : _GEN_10010; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11061 = 10'h21 == _T_27 ? _ram_T_285[287:0] : _GEN_10011; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11062 = 10'h22 == _T_27 ? _ram_T_285[287:0] : _GEN_10012; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11063 = 10'h23 == _T_27 ? _ram_T_285[287:0] : _GEN_10013; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11064 = 10'h24 == _T_27 ? _ram_T_285[287:0] : _GEN_10014; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11065 = 10'h25 == _T_27 ? _ram_T_285[287:0] : _GEN_10015; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11066 = 10'h26 == _T_27 ? _ram_T_285[287:0] : _GEN_10016; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11067 = 10'h27 == _T_27 ? _ram_T_285[287:0] : _GEN_10017; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11068 = 10'h28 == _T_27 ? _ram_T_285[287:0] : _GEN_10018; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11069 = 10'h29 == _T_27 ? _ram_T_285[287:0] : _GEN_10019; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11070 = 10'h2a == _T_27 ? _ram_T_285[287:0] : _GEN_10020; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11071 = 10'h2b == _T_27 ? _ram_T_285[287:0] : _GEN_10021; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11072 = 10'h2c == _T_27 ? _ram_T_285[287:0] : _GEN_10022; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11073 = 10'h2d == _T_27 ? _ram_T_285[287:0] : _GEN_10023; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11074 = 10'h2e == _T_27 ? _ram_T_285[287:0] : _GEN_10024; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11075 = 10'h2f == _T_27 ? _ram_T_285[287:0] : _GEN_10025; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11076 = 10'h30 == _T_27 ? _ram_T_285[287:0] : _GEN_10026; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11077 = 10'h31 == _T_27 ? _ram_T_285[287:0] : _GEN_10027; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11078 = 10'h32 == _T_27 ? _ram_T_285[287:0] : _GEN_10028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11079 = 10'h33 == _T_27 ? _ram_T_285[287:0] : _GEN_10029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11080 = 10'h34 == _T_27 ? _ram_T_285[287:0] : _GEN_10030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11081 = 10'h35 == _T_27 ? _ram_T_285[287:0] : _GEN_10031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11082 = 10'h36 == _T_27 ? _ram_T_285[287:0] : _GEN_10032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11083 = 10'h37 == _T_27 ? _ram_T_285[287:0] : _GEN_10033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11084 = 10'h38 == _T_27 ? _ram_T_285[287:0] : _GEN_10034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11085 = 10'h39 == _T_27 ? _ram_T_285[287:0] : _GEN_10035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11086 = 10'h3a == _T_27 ? _ram_T_285[287:0] : _GEN_10036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11087 = 10'h3b == _T_27 ? _ram_T_285[287:0] : _GEN_10037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11088 = 10'h3c == _T_27 ? _ram_T_285[287:0] : _GEN_10038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11089 = 10'h3d == _T_27 ? _ram_T_285[287:0] : _GEN_10039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11090 = 10'h3e == _T_27 ? _ram_T_285[287:0] : _GEN_10040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11091 = 10'h3f == _T_27 ? _ram_T_285[287:0] : _GEN_10041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11092 = 10'h40 == _T_27 ? _ram_T_285[287:0] : _GEN_10042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11093 = 10'h41 == _T_27 ? _ram_T_285[287:0] : _GEN_10043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11094 = 10'h42 == _T_27 ? _ram_T_285[287:0] : _GEN_10044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11095 = 10'h43 == _T_27 ? _ram_T_285[287:0] : _GEN_10045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11096 = 10'h44 == _T_27 ? _ram_T_285[287:0] : _GEN_10046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11097 = 10'h45 == _T_27 ? _ram_T_285[287:0] : _GEN_10047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11098 = 10'h46 == _T_27 ? _ram_T_285[287:0] : _GEN_10048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11099 = 10'h47 == _T_27 ? _ram_T_285[287:0] : _GEN_10049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11100 = 10'h48 == _T_27 ? _ram_T_285[287:0] : _GEN_10050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11101 = 10'h49 == _T_27 ? _ram_T_285[287:0] : _GEN_10051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11102 = 10'h4a == _T_27 ? _ram_T_285[287:0] : _GEN_10052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11103 = 10'h4b == _T_27 ? _ram_T_285[287:0] : _GEN_10053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11104 = 10'h4c == _T_27 ? _ram_T_285[287:0] : _GEN_10054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11105 = 10'h4d == _T_27 ? _ram_T_285[287:0] : _GEN_10055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11106 = 10'h4e == _T_27 ? _ram_T_285[287:0] : _GEN_10056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11107 = 10'h4f == _T_27 ? _ram_T_285[287:0] : _GEN_10057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11108 = 10'h50 == _T_27 ? _ram_T_285[287:0] : _GEN_10058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11109 = 10'h51 == _T_27 ? _ram_T_285[287:0] : _GEN_10059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11110 = 10'h52 == _T_27 ? _ram_T_285[287:0] : _GEN_10060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11111 = 10'h53 == _T_27 ? _ram_T_285[287:0] : _GEN_10061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11112 = 10'h54 == _T_27 ? _ram_T_285[287:0] : _GEN_10062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11113 = 10'h55 == _T_27 ? _ram_T_285[287:0] : _GEN_10063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11114 = 10'h56 == _T_27 ? _ram_T_285[287:0] : _GEN_10064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11115 = 10'h57 == _T_27 ? _ram_T_285[287:0] : _GEN_10065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11116 = 10'h58 == _T_27 ? _ram_T_285[287:0] : _GEN_10066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11117 = 10'h59 == _T_27 ? _ram_T_285[287:0] : _GEN_10067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11118 = 10'h5a == _T_27 ? _ram_T_285[287:0] : _GEN_10068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11119 = 10'h5b == _T_27 ? _ram_T_285[287:0] : _GEN_10069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11120 = 10'h5c == _T_27 ? _ram_T_285[287:0] : _GEN_10070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11121 = 10'h5d == _T_27 ? _ram_T_285[287:0] : _GEN_10071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11122 = 10'h5e == _T_27 ? _ram_T_285[287:0] : _GEN_10072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11123 = 10'h5f == _T_27 ? _ram_T_285[287:0] : _GEN_10073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11124 = 10'h60 == _T_27 ? _ram_T_285[287:0] : _GEN_10074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11125 = 10'h61 == _T_27 ? _ram_T_285[287:0] : _GEN_10075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11126 = 10'h62 == _T_27 ? _ram_T_285[287:0] : _GEN_10076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11127 = 10'h63 == _T_27 ? _ram_T_285[287:0] : _GEN_10077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11128 = 10'h64 == _T_27 ? _ram_T_285[287:0] : _GEN_10078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11129 = 10'h65 == _T_27 ? _ram_T_285[287:0] : _GEN_10079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11130 = 10'h66 == _T_27 ? _ram_T_285[287:0] : _GEN_10080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11131 = 10'h67 == _T_27 ? _ram_T_285[287:0] : _GEN_10081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11132 = 10'h68 == _T_27 ? _ram_T_285[287:0] : _GEN_10082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11133 = 10'h69 == _T_27 ? _ram_T_285[287:0] : _GEN_10083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11134 = 10'h6a == _T_27 ? _ram_T_285[287:0] : _GEN_10084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11135 = 10'h6b == _T_27 ? _ram_T_285[287:0] : _GEN_10085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11136 = 10'h6c == _T_27 ? _ram_T_285[287:0] : _GEN_10086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11137 = 10'h6d == _T_27 ? _ram_T_285[287:0] : _GEN_10087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11138 = 10'h6e == _T_27 ? _ram_T_285[287:0] : _GEN_10088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11139 = 10'h6f == _T_27 ? _ram_T_285[287:0] : _GEN_10089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11140 = 10'h70 == _T_27 ? _ram_T_285[287:0] : _GEN_10090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11141 = 10'h71 == _T_27 ? _ram_T_285[287:0] : _GEN_10091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11142 = 10'h72 == _T_27 ? _ram_T_285[287:0] : _GEN_10092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11143 = 10'h73 == _T_27 ? _ram_T_285[287:0] : _GEN_10093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11144 = 10'h74 == _T_27 ? _ram_T_285[287:0] : _GEN_10094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11145 = 10'h75 == _T_27 ? _ram_T_285[287:0] : _GEN_10095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11146 = 10'h76 == _T_27 ? _ram_T_285[287:0] : _GEN_10096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11147 = 10'h77 == _T_27 ? _ram_T_285[287:0] : _GEN_10097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11148 = 10'h78 == _T_27 ? _ram_T_285[287:0] : _GEN_10098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11149 = 10'h79 == _T_27 ? _ram_T_285[287:0] : _GEN_10099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11150 = 10'h7a == _T_27 ? _ram_T_285[287:0] : _GEN_10100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11151 = 10'h7b == _T_27 ? _ram_T_285[287:0] : _GEN_10101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11152 = 10'h7c == _T_27 ? _ram_T_285[287:0] : _GEN_10102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11153 = 10'h7d == _T_27 ? _ram_T_285[287:0] : _GEN_10103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11154 = 10'h7e == _T_27 ? _ram_T_285[287:0] : _GEN_10104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11155 = 10'h7f == _T_27 ? _ram_T_285[287:0] : _GEN_10105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11156 = 10'h80 == _T_27 ? _ram_T_285[287:0] : _GEN_10106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11157 = 10'h81 == _T_27 ? _ram_T_285[287:0] : _GEN_10107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11158 = 10'h82 == _T_27 ? _ram_T_285[287:0] : _GEN_10108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11159 = 10'h83 == _T_27 ? _ram_T_285[287:0] : _GEN_10109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11160 = 10'h84 == _T_27 ? _ram_T_285[287:0] : _GEN_10110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11161 = 10'h85 == _T_27 ? _ram_T_285[287:0] : _GEN_10111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11162 = 10'h86 == _T_27 ? _ram_T_285[287:0] : _GEN_10112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11163 = 10'h87 == _T_27 ? _ram_T_285[287:0] : _GEN_10113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11164 = 10'h88 == _T_27 ? _ram_T_285[287:0] : _GEN_10114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11165 = 10'h89 == _T_27 ? _ram_T_285[287:0] : _GEN_10115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11166 = 10'h8a == _T_27 ? _ram_T_285[287:0] : _GEN_10116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11167 = 10'h8b == _T_27 ? _ram_T_285[287:0] : _GEN_10117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11168 = 10'h8c == _T_27 ? _ram_T_285[287:0] : _GEN_10118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11169 = 10'h8d == _T_27 ? _ram_T_285[287:0] : _GEN_10119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11170 = 10'h8e == _T_27 ? _ram_T_285[287:0] : _GEN_10120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11171 = 10'h8f == _T_27 ? _ram_T_285[287:0] : _GEN_10121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11172 = 10'h90 == _T_27 ? _ram_T_285[287:0] : _GEN_10122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11173 = 10'h91 == _T_27 ? _ram_T_285[287:0] : _GEN_10123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11174 = 10'h92 == _T_27 ? _ram_T_285[287:0] : _GEN_10124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11175 = 10'h93 == _T_27 ? _ram_T_285[287:0] : _GEN_10125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11176 = 10'h94 == _T_27 ? _ram_T_285[287:0] : _GEN_10126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11177 = 10'h95 == _T_27 ? _ram_T_285[287:0] : _GEN_10127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11178 = 10'h96 == _T_27 ? _ram_T_285[287:0] : _GEN_10128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11179 = 10'h97 == _T_27 ? _ram_T_285[287:0] : _GEN_10129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11180 = 10'h98 == _T_27 ? _ram_T_285[287:0] : _GEN_10130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11181 = 10'h99 == _T_27 ? _ram_T_285[287:0] : _GEN_10131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11182 = 10'h9a == _T_27 ? _ram_T_285[287:0] : _GEN_10132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11183 = 10'h9b == _T_27 ? _ram_T_285[287:0] : _GEN_10133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11184 = 10'h9c == _T_27 ? _ram_T_285[287:0] : _GEN_10134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11185 = 10'h9d == _T_27 ? _ram_T_285[287:0] : _GEN_10135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11186 = 10'h9e == _T_27 ? _ram_T_285[287:0] : _GEN_10136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11187 = 10'h9f == _T_27 ? _ram_T_285[287:0] : _GEN_10137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11188 = 10'ha0 == _T_27 ? _ram_T_285[287:0] : _GEN_10138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11189 = 10'ha1 == _T_27 ? _ram_T_285[287:0] : _GEN_10139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11190 = 10'ha2 == _T_27 ? _ram_T_285[287:0] : _GEN_10140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11191 = 10'ha3 == _T_27 ? _ram_T_285[287:0] : _GEN_10141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11192 = 10'ha4 == _T_27 ? _ram_T_285[287:0] : _GEN_10142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11193 = 10'ha5 == _T_27 ? _ram_T_285[287:0] : _GEN_10143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11194 = 10'ha6 == _T_27 ? _ram_T_285[287:0] : _GEN_10144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11195 = 10'ha7 == _T_27 ? _ram_T_285[287:0] : _GEN_10145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11196 = 10'ha8 == _T_27 ? _ram_T_285[287:0] : _GEN_10146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11197 = 10'ha9 == _T_27 ? _ram_T_285[287:0] : _GEN_10147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11198 = 10'haa == _T_27 ? _ram_T_285[287:0] : _GEN_10148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11199 = 10'hab == _T_27 ? _ram_T_285[287:0] : _GEN_10149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11200 = 10'hac == _T_27 ? _ram_T_285[287:0] : _GEN_10150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11201 = 10'had == _T_27 ? _ram_T_285[287:0] : _GEN_10151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11202 = 10'hae == _T_27 ? _ram_T_285[287:0] : _GEN_10152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11203 = 10'haf == _T_27 ? _ram_T_285[287:0] : _GEN_10153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11204 = 10'hb0 == _T_27 ? _ram_T_285[287:0] : _GEN_10154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11205 = 10'hb1 == _T_27 ? _ram_T_285[287:0] : _GEN_10155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11206 = 10'hb2 == _T_27 ? _ram_T_285[287:0] : _GEN_10156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11207 = 10'hb3 == _T_27 ? _ram_T_285[287:0] : _GEN_10157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11208 = 10'hb4 == _T_27 ? _ram_T_285[287:0] : _GEN_10158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11209 = 10'hb5 == _T_27 ? _ram_T_285[287:0] : _GEN_10159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11210 = 10'hb6 == _T_27 ? _ram_T_285[287:0] : _GEN_10160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11211 = 10'hb7 == _T_27 ? _ram_T_285[287:0] : _GEN_10161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11212 = 10'hb8 == _T_27 ? _ram_T_285[287:0] : _GEN_10162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11213 = 10'hb9 == _T_27 ? _ram_T_285[287:0] : _GEN_10163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11214 = 10'hba == _T_27 ? _ram_T_285[287:0] : _GEN_10164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11215 = 10'hbb == _T_27 ? _ram_T_285[287:0] : _GEN_10165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11216 = 10'hbc == _T_27 ? _ram_T_285[287:0] : _GEN_10166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11217 = 10'hbd == _T_27 ? _ram_T_285[287:0] : _GEN_10167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11218 = 10'hbe == _T_27 ? _ram_T_285[287:0] : _GEN_10168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11219 = 10'hbf == _T_27 ? _ram_T_285[287:0] : _GEN_10169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11220 = 10'hc0 == _T_27 ? _ram_T_285[287:0] : _GEN_10170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11221 = 10'hc1 == _T_27 ? _ram_T_285[287:0] : _GEN_10171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11222 = 10'hc2 == _T_27 ? _ram_T_285[287:0] : _GEN_10172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11223 = 10'hc3 == _T_27 ? _ram_T_285[287:0] : _GEN_10173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11224 = 10'hc4 == _T_27 ? _ram_T_285[287:0] : _GEN_10174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11225 = 10'hc5 == _T_27 ? _ram_T_285[287:0] : _GEN_10175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11226 = 10'hc6 == _T_27 ? _ram_T_285[287:0] : _GEN_10176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11227 = 10'hc7 == _T_27 ? _ram_T_285[287:0] : _GEN_10177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11228 = 10'hc8 == _T_27 ? _ram_T_285[287:0] : _GEN_10178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11229 = 10'hc9 == _T_27 ? _ram_T_285[287:0] : _GEN_10179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11230 = 10'hca == _T_27 ? _ram_T_285[287:0] : _GEN_10180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11231 = 10'hcb == _T_27 ? _ram_T_285[287:0] : _GEN_10181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11232 = 10'hcc == _T_27 ? _ram_T_285[287:0] : _GEN_10182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11233 = 10'hcd == _T_27 ? _ram_T_285[287:0] : _GEN_10183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11234 = 10'hce == _T_27 ? _ram_T_285[287:0] : _GEN_10184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11235 = 10'hcf == _T_27 ? _ram_T_285[287:0] : _GEN_10185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11236 = 10'hd0 == _T_27 ? _ram_T_285[287:0] : _GEN_10186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11237 = 10'hd1 == _T_27 ? _ram_T_285[287:0] : _GEN_10187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11238 = 10'hd2 == _T_27 ? _ram_T_285[287:0] : _GEN_10188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11239 = 10'hd3 == _T_27 ? _ram_T_285[287:0] : _GEN_10189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11240 = 10'hd4 == _T_27 ? _ram_T_285[287:0] : _GEN_10190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11241 = 10'hd5 == _T_27 ? _ram_T_285[287:0] : _GEN_10191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11242 = 10'hd6 == _T_27 ? _ram_T_285[287:0] : _GEN_10192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11243 = 10'hd7 == _T_27 ? _ram_T_285[287:0] : _GEN_10193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11244 = 10'hd8 == _T_27 ? _ram_T_285[287:0] : _GEN_10194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11245 = 10'hd9 == _T_27 ? _ram_T_285[287:0] : _GEN_10195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11246 = 10'hda == _T_27 ? _ram_T_285[287:0] : _GEN_10196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11247 = 10'hdb == _T_27 ? _ram_T_285[287:0] : _GEN_10197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11248 = 10'hdc == _T_27 ? _ram_T_285[287:0] : _GEN_10198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11249 = 10'hdd == _T_27 ? _ram_T_285[287:0] : _GEN_10199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11250 = 10'hde == _T_27 ? _ram_T_285[287:0] : _GEN_10200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11251 = 10'hdf == _T_27 ? _ram_T_285[287:0] : _GEN_10201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11252 = 10'he0 == _T_27 ? _ram_T_285[287:0] : _GEN_10202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11253 = 10'he1 == _T_27 ? _ram_T_285[287:0] : _GEN_10203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11254 = 10'he2 == _T_27 ? _ram_T_285[287:0] : _GEN_10204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11255 = 10'he3 == _T_27 ? _ram_T_285[287:0] : _GEN_10205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11256 = 10'he4 == _T_27 ? _ram_T_285[287:0] : _GEN_10206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11257 = 10'he5 == _T_27 ? _ram_T_285[287:0] : _GEN_10207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11258 = 10'he6 == _T_27 ? _ram_T_285[287:0] : _GEN_10208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11259 = 10'he7 == _T_27 ? _ram_T_285[287:0] : _GEN_10209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11260 = 10'he8 == _T_27 ? _ram_T_285[287:0] : _GEN_10210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11261 = 10'he9 == _T_27 ? _ram_T_285[287:0] : _GEN_10211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11262 = 10'hea == _T_27 ? _ram_T_285[287:0] : _GEN_10212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11263 = 10'heb == _T_27 ? _ram_T_285[287:0] : _GEN_10213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11264 = 10'hec == _T_27 ? _ram_T_285[287:0] : _GEN_10214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11265 = 10'hed == _T_27 ? _ram_T_285[287:0] : _GEN_10215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11266 = 10'hee == _T_27 ? _ram_T_285[287:0] : _GEN_10216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11267 = 10'hef == _T_27 ? _ram_T_285[287:0] : _GEN_10217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11268 = 10'hf0 == _T_27 ? _ram_T_285[287:0] : _GEN_10218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11269 = 10'hf1 == _T_27 ? _ram_T_285[287:0] : _GEN_10219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11270 = 10'hf2 == _T_27 ? _ram_T_285[287:0] : _GEN_10220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11271 = 10'hf3 == _T_27 ? _ram_T_285[287:0] : _GEN_10221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11272 = 10'hf4 == _T_27 ? _ram_T_285[287:0] : _GEN_10222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11273 = 10'hf5 == _T_27 ? _ram_T_285[287:0] : _GEN_10223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11274 = 10'hf6 == _T_27 ? _ram_T_285[287:0] : _GEN_10224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11275 = 10'hf7 == _T_27 ? _ram_T_285[287:0] : _GEN_10225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11276 = 10'hf8 == _T_27 ? _ram_T_285[287:0] : _GEN_10226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11277 = 10'hf9 == _T_27 ? _ram_T_285[287:0] : _GEN_10227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11278 = 10'hfa == _T_27 ? _ram_T_285[287:0] : _GEN_10228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11279 = 10'hfb == _T_27 ? _ram_T_285[287:0] : _GEN_10229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11280 = 10'hfc == _T_27 ? _ram_T_285[287:0] : _GEN_10230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11281 = 10'hfd == _T_27 ? _ram_T_285[287:0] : _GEN_10231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11282 = 10'hfe == _T_27 ? _ram_T_285[287:0] : _GEN_10232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11283 = 10'hff == _T_27 ? _ram_T_285[287:0] : _GEN_10233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11284 = 10'h100 == _T_27 ? _ram_T_285[287:0] : _GEN_10234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11285 = 10'h101 == _T_27 ? _ram_T_285[287:0] : _GEN_10235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11286 = 10'h102 == _T_27 ? _ram_T_285[287:0] : _GEN_10236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11287 = 10'h103 == _T_27 ? _ram_T_285[287:0] : _GEN_10237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11288 = 10'h104 == _T_27 ? _ram_T_285[287:0] : _GEN_10238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11289 = 10'h105 == _T_27 ? _ram_T_285[287:0] : _GEN_10239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11290 = 10'h106 == _T_27 ? _ram_T_285[287:0] : _GEN_10240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11291 = 10'h107 == _T_27 ? _ram_T_285[287:0] : _GEN_10241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11292 = 10'h108 == _T_27 ? _ram_T_285[287:0] : _GEN_10242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11293 = 10'h109 == _T_27 ? _ram_T_285[287:0] : _GEN_10243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11294 = 10'h10a == _T_27 ? _ram_T_285[287:0] : _GEN_10244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11295 = 10'h10b == _T_27 ? _ram_T_285[287:0] : _GEN_10245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11296 = 10'h10c == _T_27 ? _ram_T_285[287:0] : _GEN_10246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11297 = 10'h10d == _T_27 ? _ram_T_285[287:0] : _GEN_10247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11298 = 10'h10e == _T_27 ? _ram_T_285[287:0] : _GEN_10248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11299 = 10'h10f == _T_27 ? _ram_T_285[287:0] : _GEN_10249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11300 = 10'h110 == _T_27 ? _ram_T_285[287:0] : _GEN_10250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11301 = 10'h111 == _T_27 ? _ram_T_285[287:0] : _GEN_10251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11302 = 10'h112 == _T_27 ? _ram_T_285[287:0] : _GEN_10252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11303 = 10'h113 == _T_27 ? _ram_T_285[287:0] : _GEN_10253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11304 = 10'h114 == _T_27 ? _ram_T_285[287:0] : _GEN_10254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11305 = 10'h115 == _T_27 ? _ram_T_285[287:0] : _GEN_10255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11306 = 10'h116 == _T_27 ? _ram_T_285[287:0] : _GEN_10256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11307 = 10'h117 == _T_27 ? _ram_T_285[287:0] : _GEN_10257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11308 = 10'h118 == _T_27 ? _ram_T_285[287:0] : _GEN_10258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11309 = 10'h119 == _T_27 ? _ram_T_285[287:0] : _GEN_10259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11310 = 10'h11a == _T_27 ? _ram_T_285[287:0] : _GEN_10260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11311 = 10'h11b == _T_27 ? _ram_T_285[287:0] : _GEN_10261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11312 = 10'h11c == _T_27 ? _ram_T_285[287:0] : _GEN_10262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11313 = 10'h11d == _T_27 ? _ram_T_285[287:0] : _GEN_10263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11314 = 10'h11e == _T_27 ? _ram_T_285[287:0] : _GEN_10264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11315 = 10'h11f == _T_27 ? _ram_T_285[287:0] : _GEN_10265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11316 = 10'h120 == _T_27 ? _ram_T_285[287:0] : _GEN_10266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11317 = 10'h121 == _T_27 ? _ram_T_285[287:0] : _GEN_10267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11318 = 10'h122 == _T_27 ? _ram_T_285[287:0] : _GEN_10268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11319 = 10'h123 == _T_27 ? _ram_T_285[287:0] : _GEN_10269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11320 = 10'h124 == _T_27 ? _ram_T_285[287:0] : _GEN_10270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11321 = 10'h125 == _T_27 ? _ram_T_285[287:0] : _GEN_10271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11322 = 10'h126 == _T_27 ? _ram_T_285[287:0] : _GEN_10272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11323 = 10'h127 == _T_27 ? _ram_T_285[287:0] : _GEN_10273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11324 = 10'h128 == _T_27 ? _ram_T_285[287:0] : _GEN_10274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11325 = 10'h129 == _T_27 ? _ram_T_285[287:0] : _GEN_10275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11326 = 10'h12a == _T_27 ? _ram_T_285[287:0] : _GEN_10276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11327 = 10'h12b == _T_27 ? _ram_T_285[287:0] : _GEN_10277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11328 = 10'h12c == _T_27 ? _ram_T_285[287:0] : _GEN_10278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11329 = 10'h12d == _T_27 ? _ram_T_285[287:0] : _GEN_10279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11330 = 10'h12e == _T_27 ? _ram_T_285[287:0] : _GEN_10280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11331 = 10'h12f == _T_27 ? _ram_T_285[287:0] : _GEN_10281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11332 = 10'h130 == _T_27 ? _ram_T_285[287:0] : _GEN_10282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11333 = 10'h131 == _T_27 ? _ram_T_285[287:0] : _GEN_10283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11334 = 10'h132 == _T_27 ? _ram_T_285[287:0] : _GEN_10284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11335 = 10'h133 == _T_27 ? _ram_T_285[287:0] : _GEN_10285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11336 = 10'h134 == _T_27 ? _ram_T_285[287:0] : _GEN_10286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11337 = 10'h135 == _T_27 ? _ram_T_285[287:0] : _GEN_10287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11338 = 10'h136 == _T_27 ? _ram_T_285[287:0] : _GEN_10288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11339 = 10'h137 == _T_27 ? _ram_T_285[287:0] : _GEN_10289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11340 = 10'h138 == _T_27 ? _ram_T_285[287:0] : _GEN_10290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11341 = 10'h139 == _T_27 ? _ram_T_285[287:0] : _GEN_10291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11342 = 10'h13a == _T_27 ? _ram_T_285[287:0] : _GEN_10292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11343 = 10'h13b == _T_27 ? _ram_T_285[287:0] : _GEN_10293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11344 = 10'h13c == _T_27 ? _ram_T_285[287:0] : _GEN_10294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11345 = 10'h13d == _T_27 ? _ram_T_285[287:0] : _GEN_10295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11346 = 10'h13e == _T_27 ? _ram_T_285[287:0] : _GEN_10296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11347 = 10'h13f == _T_27 ? _ram_T_285[287:0] : _GEN_10297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11348 = 10'h140 == _T_27 ? _ram_T_285[287:0] : _GEN_10298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11349 = 10'h141 == _T_27 ? _ram_T_285[287:0] : _GEN_10299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11350 = 10'h142 == _T_27 ? _ram_T_285[287:0] : _GEN_10300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11351 = 10'h143 == _T_27 ? _ram_T_285[287:0] : _GEN_10301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11352 = 10'h144 == _T_27 ? _ram_T_285[287:0] : _GEN_10302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11353 = 10'h145 == _T_27 ? _ram_T_285[287:0] : _GEN_10303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11354 = 10'h146 == _T_27 ? _ram_T_285[287:0] : _GEN_10304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11355 = 10'h147 == _T_27 ? _ram_T_285[287:0] : _GEN_10305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11356 = 10'h148 == _T_27 ? _ram_T_285[287:0] : _GEN_10306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11357 = 10'h149 == _T_27 ? _ram_T_285[287:0] : _GEN_10307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11358 = 10'h14a == _T_27 ? _ram_T_285[287:0] : _GEN_10308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11359 = 10'h14b == _T_27 ? _ram_T_285[287:0] : _GEN_10309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11360 = 10'h14c == _T_27 ? _ram_T_285[287:0] : _GEN_10310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11361 = 10'h14d == _T_27 ? _ram_T_285[287:0] : _GEN_10311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11362 = 10'h14e == _T_27 ? _ram_T_285[287:0] : _GEN_10312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11363 = 10'h14f == _T_27 ? _ram_T_285[287:0] : _GEN_10313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11364 = 10'h150 == _T_27 ? _ram_T_285[287:0] : _GEN_10314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11365 = 10'h151 == _T_27 ? _ram_T_285[287:0] : _GEN_10315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11366 = 10'h152 == _T_27 ? _ram_T_285[287:0] : _GEN_10316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11367 = 10'h153 == _T_27 ? _ram_T_285[287:0] : _GEN_10317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11368 = 10'h154 == _T_27 ? _ram_T_285[287:0] : _GEN_10318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11369 = 10'h155 == _T_27 ? _ram_T_285[287:0] : _GEN_10319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11370 = 10'h156 == _T_27 ? _ram_T_285[287:0] : _GEN_10320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11371 = 10'h157 == _T_27 ? _ram_T_285[287:0] : _GEN_10321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11372 = 10'h158 == _T_27 ? _ram_T_285[287:0] : _GEN_10322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11373 = 10'h159 == _T_27 ? _ram_T_285[287:0] : _GEN_10323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11374 = 10'h15a == _T_27 ? _ram_T_285[287:0] : _GEN_10324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11375 = 10'h15b == _T_27 ? _ram_T_285[287:0] : _GEN_10325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11376 = 10'h15c == _T_27 ? _ram_T_285[287:0] : _GEN_10326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11377 = 10'h15d == _T_27 ? _ram_T_285[287:0] : _GEN_10327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11378 = 10'h15e == _T_27 ? _ram_T_285[287:0] : _GEN_10328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11379 = 10'h15f == _T_27 ? _ram_T_285[287:0] : _GEN_10329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11380 = 10'h160 == _T_27 ? _ram_T_285[287:0] : _GEN_10330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11381 = 10'h161 == _T_27 ? _ram_T_285[287:0] : _GEN_10331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11382 = 10'h162 == _T_27 ? _ram_T_285[287:0] : _GEN_10332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11383 = 10'h163 == _T_27 ? _ram_T_285[287:0] : _GEN_10333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11384 = 10'h164 == _T_27 ? _ram_T_285[287:0] : _GEN_10334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11385 = 10'h165 == _T_27 ? _ram_T_285[287:0] : _GEN_10335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11386 = 10'h166 == _T_27 ? _ram_T_285[287:0] : _GEN_10336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11387 = 10'h167 == _T_27 ? _ram_T_285[287:0] : _GEN_10337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11388 = 10'h168 == _T_27 ? _ram_T_285[287:0] : _GEN_10338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11389 = 10'h169 == _T_27 ? _ram_T_285[287:0] : _GEN_10339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11390 = 10'h16a == _T_27 ? _ram_T_285[287:0] : _GEN_10340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11391 = 10'h16b == _T_27 ? _ram_T_285[287:0] : _GEN_10341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11392 = 10'h16c == _T_27 ? _ram_T_285[287:0] : _GEN_10342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11393 = 10'h16d == _T_27 ? _ram_T_285[287:0] : _GEN_10343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11394 = 10'h16e == _T_27 ? _ram_T_285[287:0] : _GEN_10344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11395 = 10'h16f == _T_27 ? _ram_T_285[287:0] : _GEN_10345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11396 = 10'h170 == _T_27 ? _ram_T_285[287:0] : _GEN_10346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11397 = 10'h171 == _T_27 ? _ram_T_285[287:0] : _GEN_10347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11398 = 10'h172 == _T_27 ? _ram_T_285[287:0] : _GEN_10348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11399 = 10'h173 == _T_27 ? _ram_T_285[287:0] : _GEN_10349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11400 = 10'h174 == _T_27 ? _ram_T_285[287:0] : _GEN_10350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11401 = 10'h175 == _T_27 ? _ram_T_285[287:0] : _GEN_10351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11402 = 10'h176 == _T_27 ? _ram_T_285[287:0] : _GEN_10352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11403 = 10'h177 == _T_27 ? _ram_T_285[287:0] : _GEN_10353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11404 = 10'h178 == _T_27 ? _ram_T_285[287:0] : _GEN_10354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11405 = 10'h179 == _T_27 ? _ram_T_285[287:0] : _GEN_10355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11406 = 10'h17a == _T_27 ? _ram_T_285[287:0] : _GEN_10356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11407 = 10'h17b == _T_27 ? _ram_T_285[287:0] : _GEN_10357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11408 = 10'h17c == _T_27 ? _ram_T_285[287:0] : _GEN_10358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11409 = 10'h17d == _T_27 ? _ram_T_285[287:0] : _GEN_10359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11410 = 10'h17e == _T_27 ? _ram_T_285[287:0] : _GEN_10360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11411 = 10'h17f == _T_27 ? _ram_T_285[287:0] : _GEN_10361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11412 = 10'h180 == _T_27 ? _ram_T_285[287:0] : _GEN_10362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11413 = 10'h181 == _T_27 ? _ram_T_285[287:0] : _GEN_10363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11414 = 10'h182 == _T_27 ? _ram_T_285[287:0] : _GEN_10364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11415 = 10'h183 == _T_27 ? _ram_T_285[287:0] : _GEN_10365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11416 = 10'h184 == _T_27 ? _ram_T_285[287:0] : _GEN_10366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11417 = 10'h185 == _T_27 ? _ram_T_285[287:0] : _GEN_10367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11418 = 10'h186 == _T_27 ? _ram_T_285[287:0] : _GEN_10368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11419 = 10'h187 == _T_27 ? _ram_T_285[287:0] : _GEN_10369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11420 = 10'h188 == _T_27 ? _ram_T_285[287:0] : _GEN_10370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11421 = 10'h189 == _T_27 ? _ram_T_285[287:0] : _GEN_10371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11422 = 10'h18a == _T_27 ? _ram_T_285[287:0] : _GEN_10372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11423 = 10'h18b == _T_27 ? _ram_T_285[287:0] : _GEN_10373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11424 = 10'h18c == _T_27 ? _ram_T_285[287:0] : _GEN_10374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11425 = 10'h18d == _T_27 ? _ram_T_285[287:0] : _GEN_10375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11426 = 10'h18e == _T_27 ? _ram_T_285[287:0] : _GEN_10376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11427 = 10'h18f == _T_27 ? _ram_T_285[287:0] : _GEN_10377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11428 = 10'h190 == _T_27 ? _ram_T_285[287:0] : _GEN_10378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11429 = 10'h191 == _T_27 ? _ram_T_285[287:0] : _GEN_10379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11430 = 10'h192 == _T_27 ? _ram_T_285[287:0] : _GEN_10380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11431 = 10'h193 == _T_27 ? _ram_T_285[287:0] : _GEN_10381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11432 = 10'h194 == _T_27 ? _ram_T_285[287:0] : _GEN_10382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11433 = 10'h195 == _T_27 ? _ram_T_285[287:0] : _GEN_10383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11434 = 10'h196 == _T_27 ? _ram_T_285[287:0] : _GEN_10384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11435 = 10'h197 == _T_27 ? _ram_T_285[287:0] : _GEN_10385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11436 = 10'h198 == _T_27 ? _ram_T_285[287:0] : _GEN_10386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11437 = 10'h199 == _T_27 ? _ram_T_285[287:0] : _GEN_10387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11438 = 10'h19a == _T_27 ? _ram_T_285[287:0] : _GEN_10388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11439 = 10'h19b == _T_27 ? _ram_T_285[287:0] : _GEN_10389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11440 = 10'h19c == _T_27 ? _ram_T_285[287:0] : _GEN_10390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11441 = 10'h19d == _T_27 ? _ram_T_285[287:0] : _GEN_10391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11442 = 10'h19e == _T_27 ? _ram_T_285[287:0] : _GEN_10392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11443 = 10'h19f == _T_27 ? _ram_T_285[287:0] : _GEN_10393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11444 = 10'h1a0 == _T_27 ? _ram_T_285[287:0] : _GEN_10394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11445 = 10'h1a1 == _T_27 ? _ram_T_285[287:0] : _GEN_10395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11446 = 10'h1a2 == _T_27 ? _ram_T_285[287:0] : _GEN_10396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11447 = 10'h1a3 == _T_27 ? _ram_T_285[287:0] : _GEN_10397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11448 = 10'h1a4 == _T_27 ? _ram_T_285[287:0] : _GEN_10398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11449 = 10'h1a5 == _T_27 ? _ram_T_285[287:0] : _GEN_10399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11450 = 10'h1a6 == _T_27 ? _ram_T_285[287:0] : _GEN_10400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11451 = 10'h1a7 == _T_27 ? _ram_T_285[287:0] : _GEN_10401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11452 = 10'h1a8 == _T_27 ? _ram_T_285[287:0] : _GEN_10402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11453 = 10'h1a9 == _T_27 ? _ram_T_285[287:0] : _GEN_10403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11454 = 10'h1aa == _T_27 ? _ram_T_285[287:0] : _GEN_10404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11455 = 10'h1ab == _T_27 ? _ram_T_285[287:0] : _GEN_10405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11456 = 10'h1ac == _T_27 ? _ram_T_285[287:0] : _GEN_10406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11457 = 10'h1ad == _T_27 ? _ram_T_285[287:0] : _GEN_10407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11458 = 10'h1ae == _T_27 ? _ram_T_285[287:0] : _GEN_10408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11459 = 10'h1af == _T_27 ? _ram_T_285[287:0] : _GEN_10409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11460 = 10'h1b0 == _T_27 ? _ram_T_285[287:0] : _GEN_10410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11461 = 10'h1b1 == _T_27 ? _ram_T_285[287:0] : _GEN_10411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11462 = 10'h1b2 == _T_27 ? _ram_T_285[287:0] : _GEN_10412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11463 = 10'h1b3 == _T_27 ? _ram_T_285[287:0] : _GEN_10413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11464 = 10'h1b4 == _T_27 ? _ram_T_285[287:0] : _GEN_10414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11465 = 10'h1b5 == _T_27 ? _ram_T_285[287:0] : _GEN_10415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11466 = 10'h1b6 == _T_27 ? _ram_T_285[287:0] : _GEN_10416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11467 = 10'h1b7 == _T_27 ? _ram_T_285[287:0] : _GEN_10417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11468 = 10'h1b8 == _T_27 ? _ram_T_285[287:0] : _GEN_10418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11469 = 10'h1b9 == _T_27 ? _ram_T_285[287:0] : _GEN_10419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11470 = 10'h1ba == _T_27 ? _ram_T_285[287:0] : _GEN_10420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11471 = 10'h1bb == _T_27 ? _ram_T_285[287:0] : _GEN_10421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11472 = 10'h1bc == _T_27 ? _ram_T_285[287:0] : _GEN_10422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11473 = 10'h1bd == _T_27 ? _ram_T_285[287:0] : _GEN_10423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11474 = 10'h1be == _T_27 ? _ram_T_285[287:0] : _GEN_10424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11475 = 10'h1bf == _T_27 ? _ram_T_285[287:0] : _GEN_10425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11476 = 10'h1c0 == _T_27 ? _ram_T_285[287:0] : _GEN_10426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11477 = 10'h1c1 == _T_27 ? _ram_T_285[287:0] : _GEN_10427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11478 = 10'h1c2 == _T_27 ? _ram_T_285[287:0] : _GEN_10428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11479 = 10'h1c3 == _T_27 ? _ram_T_285[287:0] : _GEN_10429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11480 = 10'h1c4 == _T_27 ? _ram_T_285[287:0] : _GEN_10430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11481 = 10'h1c5 == _T_27 ? _ram_T_285[287:0] : _GEN_10431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11482 = 10'h1c6 == _T_27 ? _ram_T_285[287:0] : _GEN_10432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11483 = 10'h1c7 == _T_27 ? _ram_T_285[287:0] : _GEN_10433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11484 = 10'h1c8 == _T_27 ? _ram_T_285[287:0] : _GEN_10434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11485 = 10'h1c9 == _T_27 ? _ram_T_285[287:0] : _GEN_10435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11486 = 10'h1ca == _T_27 ? _ram_T_285[287:0] : _GEN_10436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11487 = 10'h1cb == _T_27 ? _ram_T_285[287:0] : _GEN_10437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11488 = 10'h1cc == _T_27 ? _ram_T_285[287:0] : _GEN_10438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11489 = 10'h1cd == _T_27 ? _ram_T_285[287:0] : _GEN_10439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11490 = 10'h1ce == _T_27 ? _ram_T_285[287:0] : _GEN_10440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11491 = 10'h1cf == _T_27 ? _ram_T_285[287:0] : _GEN_10441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11492 = 10'h1d0 == _T_27 ? _ram_T_285[287:0] : _GEN_10442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11493 = 10'h1d1 == _T_27 ? _ram_T_285[287:0] : _GEN_10443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11494 = 10'h1d2 == _T_27 ? _ram_T_285[287:0] : _GEN_10444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11495 = 10'h1d3 == _T_27 ? _ram_T_285[287:0] : _GEN_10445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11496 = 10'h1d4 == _T_27 ? _ram_T_285[287:0] : _GEN_10446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11497 = 10'h1d5 == _T_27 ? _ram_T_285[287:0] : _GEN_10447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11498 = 10'h1d6 == _T_27 ? _ram_T_285[287:0] : _GEN_10448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11499 = 10'h1d7 == _T_27 ? _ram_T_285[287:0] : _GEN_10449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11500 = 10'h1d8 == _T_27 ? _ram_T_285[287:0] : _GEN_10450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11501 = 10'h1d9 == _T_27 ? _ram_T_285[287:0] : _GEN_10451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11502 = 10'h1da == _T_27 ? _ram_T_285[287:0] : _GEN_10452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11503 = 10'h1db == _T_27 ? _ram_T_285[287:0] : _GEN_10453; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11504 = 10'h1dc == _T_27 ? _ram_T_285[287:0] : _GEN_10454; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11505 = 10'h1dd == _T_27 ? _ram_T_285[287:0] : _GEN_10455; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11506 = 10'h1de == _T_27 ? _ram_T_285[287:0] : _GEN_10456; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11507 = 10'h1df == _T_27 ? _ram_T_285[287:0] : _GEN_10457; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11508 = 10'h1e0 == _T_27 ? _ram_T_285[287:0] : _GEN_10458; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11509 = 10'h1e1 == _T_27 ? _ram_T_285[287:0] : _GEN_10459; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11510 = 10'h1e2 == _T_27 ? _ram_T_285[287:0] : _GEN_10460; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11511 = 10'h1e3 == _T_27 ? _ram_T_285[287:0] : _GEN_10461; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11512 = 10'h1e4 == _T_27 ? _ram_T_285[287:0] : _GEN_10462; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11513 = 10'h1e5 == _T_27 ? _ram_T_285[287:0] : _GEN_10463; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11514 = 10'h1e6 == _T_27 ? _ram_T_285[287:0] : _GEN_10464; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11515 = 10'h1e7 == _T_27 ? _ram_T_285[287:0] : _GEN_10465; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11516 = 10'h1e8 == _T_27 ? _ram_T_285[287:0] : _GEN_10466; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11517 = 10'h1e9 == _T_27 ? _ram_T_285[287:0] : _GEN_10467; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11518 = 10'h1ea == _T_27 ? _ram_T_285[287:0] : _GEN_10468; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11519 = 10'h1eb == _T_27 ? _ram_T_285[287:0] : _GEN_10469; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11520 = 10'h1ec == _T_27 ? _ram_T_285[287:0] : _GEN_10470; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11521 = 10'h1ed == _T_27 ? _ram_T_285[287:0] : _GEN_10471; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11522 = 10'h1ee == _T_27 ? _ram_T_285[287:0] : _GEN_10472; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11523 = 10'h1ef == _T_27 ? _ram_T_285[287:0] : _GEN_10473; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11524 = 10'h1f0 == _T_27 ? _ram_T_285[287:0] : _GEN_10474; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11525 = 10'h1f1 == _T_27 ? _ram_T_285[287:0] : _GEN_10475; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11526 = 10'h1f2 == _T_27 ? _ram_T_285[287:0] : _GEN_10476; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11527 = 10'h1f3 == _T_27 ? _ram_T_285[287:0] : _GEN_10477; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11528 = 10'h1f4 == _T_27 ? _ram_T_285[287:0] : _GEN_10478; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11529 = 10'h1f5 == _T_27 ? _ram_T_285[287:0] : _GEN_10479; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11530 = 10'h1f6 == _T_27 ? _ram_T_285[287:0] : _GEN_10480; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11531 = 10'h1f7 == _T_27 ? _ram_T_285[287:0] : _GEN_10481; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11532 = 10'h1f8 == _T_27 ? _ram_T_285[287:0] : _GEN_10482; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11533 = 10'h1f9 == _T_27 ? _ram_T_285[287:0] : _GEN_10483; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11534 = 10'h1fa == _T_27 ? _ram_T_285[287:0] : _GEN_10484; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11535 = 10'h1fb == _T_27 ? _ram_T_285[287:0] : _GEN_10485; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11536 = 10'h1fc == _T_27 ? _ram_T_285[287:0] : _GEN_10486; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11537 = 10'h1fd == _T_27 ? _ram_T_285[287:0] : _GEN_10487; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11538 = 10'h1fe == _T_27 ? _ram_T_285[287:0] : _GEN_10488; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11539 = 10'h1ff == _T_27 ? _ram_T_285[287:0] : _GEN_10489; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11540 = 10'h200 == _T_27 ? _ram_T_285[287:0] : _GEN_10490; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11541 = 10'h201 == _T_27 ? _ram_T_285[287:0] : _GEN_10491; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11542 = 10'h202 == _T_27 ? _ram_T_285[287:0] : _GEN_10492; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11543 = 10'h203 == _T_27 ? _ram_T_285[287:0] : _GEN_10493; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11544 = 10'h204 == _T_27 ? _ram_T_285[287:0] : _GEN_10494; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11545 = 10'h205 == _T_27 ? _ram_T_285[287:0] : _GEN_10495; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11546 = 10'h206 == _T_27 ? _ram_T_285[287:0] : _GEN_10496; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11547 = 10'h207 == _T_27 ? _ram_T_285[287:0] : _GEN_10497; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11548 = 10'h208 == _T_27 ? _ram_T_285[287:0] : _GEN_10498; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11549 = 10'h209 == _T_27 ? _ram_T_285[287:0] : _GEN_10499; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11550 = 10'h20a == _T_27 ? _ram_T_285[287:0] : _GEN_10500; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11551 = 10'h20b == _T_27 ? _ram_T_285[287:0] : _GEN_10501; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_11552 = 10'h20c == _T_27 ? _ram_T_285[287:0] : _GEN_10502; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_29 = h + 10'hb; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_11 = vga_mem_ram_MPORT_99_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_11 = vga_mem_ram_MPORT_100_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_11 = vga_mem_ram_MPORT_101_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_11 = vga_mem_ram_MPORT_102_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_11 = vga_mem_ram_MPORT_103_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_11 = vga_mem_ram_MPORT_104_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_11 = vga_mem_ram_MPORT_105_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_11 = vga_mem_ram_MPORT_106_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_11 = vga_mem_ram_MPORT_107_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_306 = {278'h0,ram_hi_hi_hi_lo_11,ram_hi_hi_lo_11,ram_hi_lo_hi_11,ram_hi_lo_lo_11,
    ram_lo_hi_hi_hi_11,ram_lo_hi_hi_lo_11,ram_lo_hi_lo_11,ram_lo_lo_hi_11,ram_lo_lo_lo_11}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19082 = {{8191'd0}, _ram_T_306}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_310 = _GEN_19082 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_11554 = 10'h1 == _T_29 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11555 = 10'h2 == _T_29 ? ram_2 : _GEN_11554; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11556 = 10'h3 == _T_29 ? ram_3 : _GEN_11555; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11557 = 10'h4 == _T_29 ? ram_4 : _GEN_11556; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11558 = 10'h5 == _T_29 ? ram_5 : _GEN_11557; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11559 = 10'h6 == _T_29 ? ram_6 : _GEN_11558; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11560 = 10'h7 == _T_29 ? ram_7 : _GEN_11559; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11561 = 10'h8 == _T_29 ? ram_8 : _GEN_11560; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11562 = 10'h9 == _T_29 ? ram_9 : _GEN_11561; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11563 = 10'ha == _T_29 ? ram_10 : _GEN_11562; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11564 = 10'hb == _T_29 ? ram_11 : _GEN_11563; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11565 = 10'hc == _T_29 ? ram_12 : _GEN_11564; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11566 = 10'hd == _T_29 ? ram_13 : _GEN_11565; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11567 = 10'he == _T_29 ? ram_14 : _GEN_11566; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11568 = 10'hf == _T_29 ? ram_15 : _GEN_11567; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11569 = 10'h10 == _T_29 ? ram_16 : _GEN_11568; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11570 = 10'h11 == _T_29 ? ram_17 : _GEN_11569; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11571 = 10'h12 == _T_29 ? ram_18 : _GEN_11570; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11572 = 10'h13 == _T_29 ? ram_19 : _GEN_11571; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11573 = 10'h14 == _T_29 ? ram_20 : _GEN_11572; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11574 = 10'h15 == _T_29 ? ram_21 : _GEN_11573; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11575 = 10'h16 == _T_29 ? ram_22 : _GEN_11574; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11576 = 10'h17 == _T_29 ? ram_23 : _GEN_11575; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11577 = 10'h18 == _T_29 ? ram_24 : _GEN_11576; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11578 = 10'h19 == _T_29 ? ram_25 : _GEN_11577; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11579 = 10'h1a == _T_29 ? ram_26 : _GEN_11578; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11580 = 10'h1b == _T_29 ? ram_27 : _GEN_11579; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11581 = 10'h1c == _T_29 ? ram_28 : _GEN_11580; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11582 = 10'h1d == _T_29 ? ram_29 : _GEN_11581; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11583 = 10'h1e == _T_29 ? ram_30 : _GEN_11582; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11584 = 10'h1f == _T_29 ? ram_31 : _GEN_11583; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11585 = 10'h20 == _T_29 ? ram_32 : _GEN_11584; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11586 = 10'h21 == _T_29 ? ram_33 : _GEN_11585; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11587 = 10'h22 == _T_29 ? ram_34 : _GEN_11586; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11588 = 10'h23 == _T_29 ? ram_35 : _GEN_11587; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11589 = 10'h24 == _T_29 ? ram_36 : _GEN_11588; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11590 = 10'h25 == _T_29 ? ram_37 : _GEN_11589; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11591 = 10'h26 == _T_29 ? ram_38 : _GEN_11590; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11592 = 10'h27 == _T_29 ? ram_39 : _GEN_11591; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11593 = 10'h28 == _T_29 ? ram_40 : _GEN_11592; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11594 = 10'h29 == _T_29 ? ram_41 : _GEN_11593; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11595 = 10'h2a == _T_29 ? ram_42 : _GEN_11594; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11596 = 10'h2b == _T_29 ? ram_43 : _GEN_11595; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11597 = 10'h2c == _T_29 ? ram_44 : _GEN_11596; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11598 = 10'h2d == _T_29 ? ram_45 : _GEN_11597; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11599 = 10'h2e == _T_29 ? ram_46 : _GEN_11598; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11600 = 10'h2f == _T_29 ? ram_47 : _GEN_11599; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11601 = 10'h30 == _T_29 ? ram_48 : _GEN_11600; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11602 = 10'h31 == _T_29 ? ram_49 : _GEN_11601; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11603 = 10'h32 == _T_29 ? ram_50 : _GEN_11602; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11604 = 10'h33 == _T_29 ? ram_51 : _GEN_11603; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11605 = 10'h34 == _T_29 ? ram_52 : _GEN_11604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11606 = 10'h35 == _T_29 ? ram_53 : _GEN_11605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11607 = 10'h36 == _T_29 ? ram_54 : _GEN_11606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11608 = 10'h37 == _T_29 ? ram_55 : _GEN_11607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11609 = 10'h38 == _T_29 ? ram_56 : _GEN_11608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11610 = 10'h39 == _T_29 ? ram_57 : _GEN_11609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11611 = 10'h3a == _T_29 ? ram_58 : _GEN_11610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11612 = 10'h3b == _T_29 ? ram_59 : _GEN_11611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11613 = 10'h3c == _T_29 ? ram_60 : _GEN_11612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11614 = 10'h3d == _T_29 ? ram_61 : _GEN_11613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11615 = 10'h3e == _T_29 ? ram_62 : _GEN_11614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11616 = 10'h3f == _T_29 ? ram_63 : _GEN_11615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11617 = 10'h40 == _T_29 ? ram_64 : _GEN_11616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11618 = 10'h41 == _T_29 ? ram_65 : _GEN_11617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11619 = 10'h42 == _T_29 ? ram_66 : _GEN_11618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11620 = 10'h43 == _T_29 ? ram_67 : _GEN_11619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11621 = 10'h44 == _T_29 ? ram_68 : _GEN_11620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11622 = 10'h45 == _T_29 ? ram_69 : _GEN_11621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11623 = 10'h46 == _T_29 ? ram_70 : _GEN_11622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11624 = 10'h47 == _T_29 ? ram_71 : _GEN_11623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11625 = 10'h48 == _T_29 ? ram_72 : _GEN_11624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11626 = 10'h49 == _T_29 ? ram_73 : _GEN_11625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11627 = 10'h4a == _T_29 ? ram_74 : _GEN_11626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11628 = 10'h4b == _T_29 ? ram_75 : _GEN_11627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11629 = 10'h4c == _T_29 ? ram_76 : _GEN_11628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11630 = 10'h4d == _T_29 ? ram_77 : _GEN_11629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11631 = 10'h4e == _T_29 ? ram_78 : _GEN_11630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11632 = 10'h4f == _T_29 ? ram_79 : _GEN_11631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11633 = 10'h50 == _T_29 ? ram_80 : _GEN_11632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11634 = 10'h51 == _T_29 ? ram_81 : _GEN_11633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11635 = 10'h52 == _T_29 ? ram_82 : _GEN_11634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11636 = 10'h53 == _T_29 ? ram_83 : _GEN_11635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11637 = 10'h54 == _T_29 ? ram_84 : _GEN_11636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11638 = 10'h55 == _T_29 ? ram_85 : _GEN_11637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11639 = 10'h56 == _T_29 ? ram_86 : _GEN_11638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11640 = 10'h57 == _T_29 ? ram_87 : _GEN_11639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11641 = 10'h58 == _T_29 ? ram_88 : _GEN_11640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11642 = 10'h59 == _T_29 ? ram_89 : _GEN_11641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11643 = 10'h5a == _T_29 ? ram_90 : _GEN_11642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11644 = 10'h5b == _T_29 ? ram_91 : _GEN_11643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11645 = 10'h5c == _T_29 ? ram_92 : _GEN_11644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11646 = 10'h5d == _T_29 ? ram_93 : _GEN_11645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11647 = 10'h5e == _T_29 ? ram_94 : _GEN_11646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11648 = 10'h5f == _T_29 ? ram_95 : _GEN_11647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11649 = 10'h60 == _T_29 ? ram_96 : _GEN_11648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11650 = 10'h61 == _T_29 ? ram_97 : _GEN_11649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11651 = 10'h62 == _T_29 ? ram_98 : _GEN_11650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11652 = 10'h63 == _T_29 ? ram_99 : _GEN_11651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11653 = 10'h64 == _T_29 ? ram_100 : _GEN_11652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11654 = 10'h65 == _T_29 ? ram_101 : _GEN_11653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11655 = 10'h66 == _T_29 ? ram_102 : _GEN_11654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11656 = 10'h67 == _T_29 ? ram_103 : _GEN_11655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11657 = 10'h68 == _T_29 ? ram_104 : _GEN_11656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11658 = 10'h69 == _T_29 ? ram_105 : _GEN_11657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11659 = 10'h6a == _T_29 ? ram_106 : _GEN_11658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11660 = 10'h6b == _T_29 ? ram_107 : _GEN_11659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11661 = 10'h6c == _T_29 ? ram_108 : _GEN_11660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11662 = 10'h6d == _T_29 ? ram_109 : _GEN_11661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11663 = 10'h6e == _T_29 ? ram_110 : _GEN_11662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11664 = 10'h6f == _T_29 ? ram_111 : _GEN_11663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11665 = 10'h70 == _T_29 ? ram_112 : _GEN_11664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11666 = 10'h71 == _T_29 ? ram_113 : _GEN_11665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11667 = 10'h72 == _T_29 ? ram_114 : _GEN_11666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11668 = 10'h73 == _T_29 ? ram_115 : _GEN_11667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11669 = 10'h74 == _T_29 ? ram_116 : _GEN_11668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11670 = 10'h75 == _T_29 ? ram_117 : _GEN_11669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11671 = 10'h76 == _T_29 ? ram_118 : _GEN_11670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11672 = 10'h77 == _T_29 ? ram_119 : _GEN_11671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11673 = 10'h78 == _T_29 ? ram_120 : _GEN_11672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11674 = 10'h79 == _T_29 ? ram_121 : _GEN_11673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11675 = 10'h7a == _T_29 ? ram_122 : _GEN_11674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11676 = 10'h7b == _T_29 ? ram_123 : _GEN_11675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11677 = 10'h7c == _T_29 ? ram_124 : _GEN_11676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11678 = 10'h7d == _T_29 ? ram_125 : _GEN_11677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11679 = 10'h7e == _T_29 ? ram_126 : _GEN_11678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11680 = 10'h7f == _T_29 ? ram_127 : _GEN_11679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11681 = 10'h80 == _T_29 ? ram_128 : _GEN_11680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11682 = 10'h81 == _T_29 ? ram_129 : _GEN_11681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11683 = 10'h82 == _T_29 ? ram_130 : _GEN_11682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11684 = 10'h83 == _T_29 ? ram_131 : _GEN_11683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11685 = 10'h84 == _T_29 ? ram_132 : _GEN_11684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11686 = 10'h85 == _T_29 ? ram_133 : _GEN_11685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11687 = 10'h86 == _T_29 ? ram_134 : _GEN_11686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11688 = 10'h87 == _T_29 ? ram_135 : _GEN_11687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11689 = 10'h88 == _T_29 ? ram_136 : _GEN_11688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11690 = 10'h89 == _T_29 ? ram_137 : _GEN_11689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11691 = 10'h8a == _T_29 ? ram_138 : _GEN_11690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11692 = 10'h8b == _T_29 ? ram_139 : _GEN_11691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11693 = 10'h8c == _T_29 ? ram_140 : _GEN_11692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11694 = 10'h8d == _T_29 ? ram_141 : _GEN_11693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11695 = 10'h8e == _T_29 ? ram_142 : _GEN_11694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11696 = 10'h8f == _T_29 ? ram_143 : _GEN_11695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11697 = 10'h90 == _T_29 ? ram_144 : _GEN_11696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11698 = 10'h91 == _T_29 ? ram_145 : _GEN_11697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11699 = 10'h92 == _T_29 ? ram_146 : _GEN_11698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11700 = 10'h93 == _T_29 ? ram_147 : _GEN_11699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11701 = 10'h94 == _T_29 ? ram_148 : _GEN_11700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11702 = 10'h95 == _T_29 ? ram_149 : _GEN_11701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11703 = 10'h96 == _T_29 ? ram_150 : _GEN_11702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11704 = 10'h97 == _T_29 ? ram_151 : _GEN_11703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11705 = 10'h98 == _T_29 ? ram_152 : _GEN_11704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11706 = 10'h99 == _T_29 ? ram_153 : _GEN_11705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11707 = 10'h9a == _T_29 ? ram_154 : _GEN_11706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11708 = 10'h9b == _T_29 ? ram_155 : _GEN_11707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11709 = 10'h9c == _T_29 ? ram_156 : _GEN_11708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11710 = 10'h9d == _T_29 ? ram_157 : _GEN_11709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11711 = 10'h9e == _T_29 ? ram_158 : _GEN_11710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11712 = 10'h9f == _T_29 ? ram_159 : _GEN_11711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11713 = 10'ha0 == _T_29 ? ram_160 : _GEN_11712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11714 = 10'ha1 == _T_29 ? ram_161 : _GEN_11713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11715 = 10'ha2 == _T_29 ? ram_162 : _GEN_11714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11716 = 10'ha3 == _T_29 ? ram_163 : _GEN_11715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11717 = 10'ha4 == _T_29 ? ram_164 : _GEN_11716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11718 = 10'ha5 == _T_29 ? ram_165 : _GEN_11717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11719 = 10'ha6 == _T_29 ? ram_166 : _GEN_11718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11720 = 10'ha7 == _T_29 ? ram_167 : _GEN_11719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11721 = 10'ha8 == _T_29 ? ram_168 : _GEN_11720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11722 = 10'ha9 == _T_29 ? ram_169 : _GEN_11721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11723 = 10'haa == _T_29 ? ram_170 : _GEN_11722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11724 = 10'hab == _T_29 ? ram_171 : _GEN_11723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11725 = 10'hac == _T_29 ? ram_172 : _GEN_11724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11726 = 10'had == _T_29 ? ram_173 : _GEN_11725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11727 = 10'hae == _T_29 ? ram_174 : _GEN_11726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11728 = 10'haf == _T_29 ? ram_175 : _GEN_11727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11729 = 10'hb0 == _T_29 ? ram_176 : _GEN_11728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11730 = 10'hb1 == _T_29 ? ram_177 : _GEN_11729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11731 = 10'hb2 == _T_29 ? ram_178 : _GEN_11730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11732 = 10'hb3 == _T_29 ? ram_179 : _GEN_11731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11733 = 10'hb4 == _T_29 ? ram_180 : _GEN_11732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11734 = 10'hb5 == _T_29 ? ram_181 : _GEN_11733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11735 = 10'hb6 == _T_29 ? ram_182 : _GEN_11734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11736 = 10'hb7 == _T_29 ? ram_183 : _GEN_11735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11737 = 10'hb8 == _T_29 ? ram_184 : _GEN_11736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11738 = 10'hb9 == _T_29 ? ram_185 : _GEN_11737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11739 = 10'hba == _T_29 ? ram_186 : _GEN_11738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11740 = 10'hbb == _T_29 ? ram_187 : _GEN_11739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11741 = 10'hbc == _T_29 ? ram_188 : _GEN_11740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11742 = 10'hbd == _T_29 ? ram_189 : _GEN_11741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11743 = 10'hbe == _T_29 ? ram_190 : _GEN_11742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11744 = 10'hbf == _T_29 ? ram_191 : _GEN_11743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11745 = 10'hc0 == _T_29 ? ram_192 : _GEN_11744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11746 = 10'hc1 == _T_29 ? ram_193 : _GEN_11745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11747 = 10'hc2 == _T_29 ? ram_194 : _GEN_11746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11748 = 10'hc3 == _T_29 ? ram_195 : _GEN_11747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11749 = 10'hc4 == _T_29 ? ram_196 : _GEN_11748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11750 = 10'hc5 == _T_29 ? ram_197 : _GEN_11749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11751 = 10'hc6 == _T_29 ? ram_198 : _GEN_11750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11752 = 10'hc7 == _T_29 ? ram_199 : _GEN_11751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11753 = 10'hc8 == _T_29 ? ram_200 : _GEN_11752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11754 = 10'hc9 == _T_29 ? ram_201 : _GEN_11753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11755 = 10'hca == _T_29 ? ram_202 : _GEN_11754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11756 = 10'hcb == _T_29 ? ram_203 : _GEN_11755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11757 = 10'hcc == _T_29 ? ram_204 : _GEN_11756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11758 = 10'hcd == _T_29 ? ram_205 : _GEN_11757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11759 = 10'hce == _T_29 ? ram_206 : _GEN_11758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11760 = 10'hcf == _T_29 ? ram_207 : _GEN_11759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11761 = 10'hd0 == _T_29 ? ram_208 : _GEN_11760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11762 = 10'hd1 == _T_29 ? ram_209 : _GEN_11761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11763 = 10'hd2 == _T_29 ? ram_210 : _GEN_11762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11764 = 10'hd3 == _T_29 ? ram_211 : _GEN_11763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11765 = 10'hd4 == _T_29 ? ram_212 : _GEN_11764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11766 = 10'hd5 == _T_29 ? ram_213 : _GEN_11765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11767 = 10'hd6 == _T_29 ? ram_214 : _GEN_11766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11768 = 10'hd7 == _T_29 ? ram_215 : _GEN_11767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11769 = 10'hd8 == _T_29 ? ram_216 : _GEN_11768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11770 = 10'hd9 == _T_29 ? ram_217 : _GEN_11769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11771 = 10'hda == _T_29 ? ram_218 : _GEN_11770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11772 = 10'hdb == _T_29 ? ram_219 : _GEN_11771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11773 = 10'hdc == _T_29 ? ram_220 : _GEN_11772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11774 = 10'hdd == _T_29 ? ram_221 : _GEN_11773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11775 = 10'hde == _T_29 ? ram_222 : _GEN_11774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11776 = 10'hdf == _T_29 ? ram_223 : _GEN_11775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11777 = 10'he0 == _T_29 ? ram_224 : _GEN_11776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11778 = 10'he1 == _T_29 ? ram_225 : _GEN_11777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11779 = 10'he2 == _T_29 ? ram_226 : _GEN_11778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11780 = 10'he3 == _T_29 ? ram_227 : _GEN_11779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11781 = 10'he4 == _T_29 ? ram_228 : _GEN_11780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11782 = 10'he5 == _T_29 ? ram_229 : _GEN_11781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11783 = 10'he6 == _T_29 ? ram_230 : _GEN_11782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11784 = 10'he7 == _T_29 ? ram_231 : _GEN_11783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11785 = 10'he8 == _T_29 ? ram_232 : _GEN_11784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11786 = 10'he9 == _T_29 ? ram_233 : _GEN_11785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11787 = 10'hea == _T_29 ? ram_234 : _GEN_11786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11788 = 10'heb == _T_29 ? ram_235 : _GEN_11787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11789 = 10'hec == _T_29 ? ram_236 : _GEN_11788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11790 = 10'hed == _T_29 ? ram_237 : _GEN_11789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11791 = 10'hee == _T_29 ? ram_238 : _GEN_11790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11792 = 10'hef == _T_29 ? ram_239 : _GEN_11791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11793 = 10'hf0 == _T_29 ? ram_240 : _GEN_11792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11794 = 10'hf1 == _T_29 ? ram_241 : _GEN_11793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11795 = 10'hf2 == _T_29 ? ram_242 : _GEN_11794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11796 = 10'hf3 == _T_29 ? ram_243 : _GEN_11795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11797 = 10'hf4 == _T_29 ? ram_244 : _GEN_11796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11798 = 10'hf5 == _T_29 ? ram_245 : _GEN_11797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11799 = 10'hf6 == _T_29 ? ram_246 : _GEN_11798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11800 = 10'hf7 == _T_29 ? ram_247 : _GEN_11799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11801 = 10'hf8 == _T_29 ? ram_248 : _GEN_11800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11802 = 10'hf9 == _T_29 ? ram_249 : _GEN_11801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11803 = 10'hfa == _T_29 ? ram_250 : _GEN_11802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11804 = 10'hfb == _T_29 ? ram_251 : _GEN_11803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11805 = 10'hfc == _T_29 ? ram_252 : _GEN_11804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11806 = 10'hfd == _T_29 ? ram_253 : _GEN_11805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11807 = 10'hfe == _T_29 ? ram_254 : _GEN_11806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11808 = 10'hff == _T_29 ? ram_255 : _GEN_11807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11809 = 10'h100 == _T_29 ? ram_256 : _GEN_11808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11810 = 10'h101 == _T_29 ? ram_257 : _GEN_11809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11811 = 10'h102 == _T_29 ? ram_258 : _GEN_11810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11812 = 10'h103 == _T_29 ? ram_259 : _GEN_11811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11813 = 10'h104 == _T_29 ? ram_260 : _GEN_11812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11814 = 10'h105 == _T_29 ? ram_261 : _GEN_11813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11815 = 10'h106 == _T_29 ? ram_262 : _GEN_11814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11816 = 10'h107 == _T_29 ? ram_263 : _GEN_11815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11817 = 10'h108 == _T_29 ? ram_264 : _GEN_11816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11818 = 10'h109 == _T_29 ? ram_265 : _GEN_11817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11819 = 10'h10a == _T_29 ? ram_266 : _GEN_11818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11820 = 10'h10b == _T_29 ? ram_267 : _GEN_11819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11821 = 10'h10c == _T_29 ? ram_268 : _GEN_11820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11822 = 10'h10d == _T_29 ? ram_269 : _GEN_11821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11823 = 10'h10e == _T_29 ? ram_270 : _GEN_11822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11824 = 10'h10f == _T_29 ? ram_271 : _GEN_11823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11825 = 10'h110 == _T_29 ? ram_272 : _GEN_11824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11826 = 10'h111 == _T_29 ? ram_273 : _GEN_11825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11827 = 10'h112 == _T_29 ? ram_274 : _GEN_11826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11828 = 10'h113 == _T_29 ? ram_275 : _GEN_11827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11829 = 10'h114 == _T_29 ? ram_276 : _GEN_11828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11830 = 10'h115 == _T_29 ? ram_277 : _GEN_11829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11831 = 10'h116 == _T_29 ? ram_278 : _GEN_11830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11832 = 10'h117 == _T_29 ? ram_279 : _GEN_11831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11833 = 10'h118 == _T_29 ? ram_280 : _GEN_11832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11834 = 10'h119 == _T_29 ? ram_281 : _GEN_11833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11835 = 10'h11a == _T_29 ? ram_282 : _GEN_11834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11836 = 10'h11b == _T_29 ? ram_283 : _GEN_11835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11837 = 10'h11c == _T_29 ? ram_284 : _GEN_11836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11838 = 10'h11d == _T_29 ? ram_285 : _GEN_11837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11839 = 10'h11e == _T_29 ? ram_286 : _GEN_11838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11840 = 10'h11f == _T_29 ? ram_287 : _GEN_11839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11841 = 10'h120 == _T_29 ? ram_288 : _GEN_11840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11842 = 10'h121 == _T_29 ? ram_289 : _GEN_11841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11843 = 10'h122 == _T_29 ? ram_290 : _GEN_11842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11844 = 10'h123 == _T_29 ? ram_291 : _GEN_11843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11845 = 10'h124 == _T_29 ? ram_292 : _GEN_11844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11846 = 10'h125 == _T_29 ? ram_293 : _GEN_11845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11847 = 10'h126 == _T_29 ? ram_294 : _GEN_11846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11848 = 10'h127 == _T_29 ? ram_295 : _GEN_11847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11849 = 10'h128 == _T_29 ? ram_296 : _GEN_11848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11850 = 10'h129 == _T_29 ? ram_297 : _GEN_11849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11851 = 10'h12a == _T_29 ? ram_298 : _GEN_11850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11852 = 10'h12b == _T_29 ? ram_299 : _GEN_11851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11853 = 10'h12c == _T_29 ? ram_300 : _GEN_11852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11854 = 10'h12d == _T_29 ? ram_301 : _GEN_11853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11855 = 10'h12e == _T_29 ? ram_302 : _GEN_11854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11856 = 10'h12f == _T_29 ? ram_303 : _GEN_11855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11857 = 10'h130 == _T_29 ? ram_304 : _GEN_11856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11858 = 10'h131 == _T_29 ? ram_305 : _GEN_11857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11859 = 10'h132 == _T_29 ? ram_306 : _GEN_11858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11860 = 10'h133 == _T_29 ? ram_307 : _GEN_11859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11861 = 10'h134 == _T_29 ? ram_308 : _GEN_11860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11862 = 10'h135 == _T_29 ? ram_309 : _GEN_11861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11863 = 10'h136 == _T_29 ? ram_310 : _GEN_11862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11864 = 10'h137 == _T_29 ? ram_311 : _GEN_11863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11865 = 10'h138 == _T_29 ? ram_312 : _GEN_11864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11866 = 10'h139 == _T_29 ? ram_313 : _GEN_11865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11867 = 10'h13a == _T_29 ? ram_314 : _GEN_11866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11868 = 10'h13b == _T_29 ? ram_315 : _GEN_11867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11869 = 10'h13c == _T_29 ? ram_316 : _GEN_11868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11870 = 10'h13d == _T_29 ? ram_317 : _GEN_11869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11871 = 10'h13e == _T_29 ? ram_318 : _GEN_11870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11872 = 10'h13f == _T_29 ? ram_319 : _GEN_11871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11873 = 10'h140 == _T_29 ? ram_320 : _GEN_11872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11874 = 10'h141 == _T_29 ? ram_321 : _GEN_11873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11875 = 10'h142 == _T_29 ? ram_322 : _GEN_11874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11876 = 10'h143 == _T_29 ? ram_323 : _GEN_11875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11877 = 10'h144 == _T_29 ? ram_324 : _GEN_11876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11878 = 10'h145 == _T_29 ? ram_325 : _GEN_11877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11879 = 10'h146 == _T_29 ? ram_326 : _GEN_11878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11880 = 10'h147 == _T_29 ? ram_327 : _GEN_11879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11881 = 10'h148 == _T_29 ? ram_328 : _GEN_11880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11882 = 10'h149 == _T_29 ? ram_329 : _GEN_11881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11883 = 10'h14a == _T_29 ? ram_330 : _GEN_11882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11884 = 10'h14b == _T_29 ? ram_331 : _GEN_11883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11885 = 10'h14c == _T_29 ? ram_332 : _GEN_11884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11886 = 10'h14d == _T_29 ? ram_333 : _GEN_11885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11887 = 10'h14e == _T_29 ? ram_334 : _GEN_11886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11888 = 10'h14f == _T_29 ? ram_335 : _GEN_11887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11889 = 10'h150 == _T_29 ? ram_336 : _GEN_11888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11890 = 10'h151 == _T_29 ? ram_337 : _GEN_11889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11891 = 10'h152 == _T_29 ? ram_338 : _GEN_11890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11892 = 10'h153 == _T_29 ? ram_339 : _GEN_11891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11893 = 10'h154 == _T_29 ? ram_340 : _GEN_11892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11894 = 10'h155 == _T_29 ? ram_341 : _GEN_11893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11895 = 10'h156 == _T_29 ? ram_342 : _GEN_11894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11896 = 10'h157 == _T_29 ? ram_343 : _GEN_11895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11897 = 10'h158 == _T_29 ? ram_344 : _GEN_11896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11898 = 10'h159 == _T_29 ? ram_345 : _GEN_11897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11899 = 10'h15a == _T_29 ? ram_346 : _GEN_11898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11900 = 10'h15b == _T_29 ? ram_347 : _GEN_11899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11901 = 10'h15c == _T_29 ? ram_348 : _GEN_11900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11902 = 10'h15d == _T_29 ? ram_349 : _GEN_11901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11903 = 10'h15e == _T_29 ? ram_350 : _GEN_11902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11904 = 10'h15f == _T_29 ? ram_351 : _GEN_11903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11905 = 10'h160 == _T_29 ? ram_352 : _GEN_11904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11906 = 10'h161 == _T_29 ? ram_353 : _GEN_11905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11907 = 10'h162 == _T_29 ? ram_354 : _GEN_11906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11908 = 10'h163 == _T_29 ? ram_355 : _GEN_11907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11909 = 10'h164 == _T_29 ? ram_356 : _GEN_11908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11910 = 10'h165 == _T_29 ? ram_357 : _GEN_11909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11911 = 10'h166 == _T_29 ? ram_358 : _GEN_11910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11912 = 10'h167 == _T_29 ? ram_359 : _GEN_11911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11913 = 10'h168 == _T_29 ? ram_360 : _GEN_11912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11914 = 10'h169 == _T_29 ? ram_361 : _GEN_11913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11915 = 10'h16a == _T_29 ? ram_362 : _GEN_11914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11916 = 10'h16b == _T_29 ? ram_363 : _GEN_11915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11917 = 10'h16c == _T_29 ? ram_364 : _GEN_11916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11918 = 10'h16d == _T_29 ? ram_365 : _GEN_11917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11919 = 10'h16e == _T_29 ? ram_366 : _GEN_11918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11920 = 10'h16f == _T_29 ? ram_367 : _GEN_11919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11921 = 10'h170 == _T_29 ? ram_368 : _GEN_11920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11922 = 10'h171 == _T_29 ? ram_369 : _GEN_11921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11923 = 10'h172 == _T_29 ? ram_370 : _GEN_11922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11924 = 10'h173 == _T_29 ? ram_371 : _GEN_11923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11925 = 10'h174 == _T_29 ? ram_372 : _GEN_11924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11926 = 10'h175 == _T_29 ? ram_373 : _GEN_11925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11927 = 10'h176 == _T_29 ? ram_374 : _GEN_11926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11928 = 10'h177 == _T_29 ? ram_375 : _GEN_11927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11929 = 10'h178 == _T_29 ? ram_376 : _GEN_11928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11930 = 10'h179 == _T_29 ? ram_377 : _GEN_11929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11931 = 10'h17a == _T_29 ? ram_378 : _GEN_11930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11932 = 10'h17b == _T_29 ? ram_379 : _GEN_11931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11933 = 10'h17c == _T_29 ? ram_380 : _GEN_11932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11934 = 10'h17d == _T_29 ? ram_381 : _GEN_11933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11935 = 10'h17e == _T_29 ? ram_382 : _GEN_11934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11936 = 10'h17f == _T_29 ? ram_383 : _GEN_11935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11937 = 10'h180 == _T_29 ? ram_384 : _GEN_11936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11938 = 10'h181 == _T_29 ? ram_385 : _GEN_11937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11939 = 10'h182 == _T_29 ? ram_386 : _GEN_11938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11940 = 10'h183 == _T_29 ? ram_387 : _GEN_11939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11941 = 10'h184 == _T_29 ? ram_388 : _GEN_11940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11942 = 10'h185 == _T_29 ? ram_389 : _GEN_11941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11943 = 10'h186 == _T_29 ? ram_390 : _GEN_11942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11944 = 10'h187 == _T_29 ? ram_391 : _GEN_11943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11945 = 10'h188 == _T_29 ? ram_392 : _GEN_11944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11946 = 10'h189 == _T_29 ? ram_393 : _GEN_11945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11947 = 10'h18a == _T_29 ? ram_394 : _GEN_11946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11948 = 10'h18b == _T_29 ? ram_395 : _GEN_11947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11949 = 10'h18c == _T_29 ? ram_396 : _GEN_11948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11950 = 10'h18d == _T_29 ? ram_397 : _GEN_11949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11951 = 10'h18e == _T_29 ? ram_398 : _GEN_11950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11952 = 10'h18f == _T_29 ? ram_399 : _GEN_11951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11953 = 10'h190 == _T_29 ? ram_400 : _GEN_11952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11954 = 10'h191 == _T_29 ? ram_401 : _GEN_11953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11955 = 10'h192 == _T_29 ? ram_402 : _GEN_11954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11956 = 10'h193 == _T_29 ? ram_403 : _GEN_11955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11957 = 10'h194 == _T_29 ? ram_404 : _GEN_11956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11958 = 10'h195 == _T_29 ? ram_405 : _GEN_11957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11959 = 10'h196 == _T_29 ? ram_406 : _GEN_11958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11960 = 10'h197 == _T_29 ? ram_407 : _GEN_11959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11961 = 10'h198 == _T_29 ? ram_408 : _GEN_11960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11962 = 10'h199 == _T_29 ? ram_409 : _GEN_11961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11963 = 10'h19a == _T_29 ? ram_410 : _GEN_11962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11964 = 10'h19b == _T_29 ? ram_411 : _GEN_11963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11965 = 10'h19c == _T_29 ? ram_412 : _GEN_11964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11966 = 10'h19d == _T_29 ? ram_413 : _GEN_11965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11967 = 10'h19e == _T_29 ? ram_414 : _GEN_11966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11968 = 10'h19f == _T_29 ? ram_415 : _GEN_11967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11969 = 10'h1a0 == _T_29 ? ram_416 : _GEN_11968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11970 = 10'h1a1 == _T_29 ? ram_417 : _GEN_11969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11971 = 10'h1a2 == _T_29 ? ram_418 : _GEN_11970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11972 = 10'h1a3 == _T_29 ? ram_419 : _GEN_11971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11973 = 10'h1a4 == _T_29 ? ram_420 : _GEN_11972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11974 = 10'h1a5 == _T_29 ? ram_421 : _GEN_11973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11975 = 10'h1a6 == _T_29 ? ram_422 : _GEN_11974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11976 = 10'h1a7 == _T_29 ? ram_423 : _GEN_11975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11977 = 10'h1a8 == _T_29 ? ram_424 : _GEN_11976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11978 = 10'h1a9 == _T_29 ? ram_425 : _GEN_11977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11979 = 10'h1aa == _T_29 ? ram_426 : _GEN_11978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11980 = 10'h1ab == _T_29 ? ram_427 : _GEN_11979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11981 = 10'h1ac == _T_29 ? ram_428 : _GEN_11980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11982 = 10'h1ad == _T_29 ? ram_429 : _GEN_11981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11983 = 10'h1ae == _T_29 ? ram_430 : _GEN_11982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11984 = 10'h1af == _T_29 ? ram_431 : _GEN_11983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11985 = 10'h1b0 == _T_29 ? ram_432 : _GEN_11984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11986 = 10'h1b1 == _T_29 ? ram_433 : _GEN_11985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11987 = 10'h1b2 == _T_29 ? ram_434 : _GEN_11986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11988 = 10'h1b3 == _T_29 ? ram_435 : _GEN_11987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11989 = 10'h1b4 == _T_29 ? ram_436 : _GEN_11988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11990 = 10'h1b5 == _T_29 ? ram_437 : _GEN_11989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11991 = 10'h1b6 == _T_29 ? ram_438 : _GEN_11990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11992 = 10'h1b7 == _T_29 ? ram_439 : _GEN_11991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11993 = 10'h1b8 == _T_29 ? ram_440 : _GEN_11992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11994 = 10'h1b9 == _T_29 ? ram_441 : _GEN_11993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11995 = 10'h1ba == _T_29 ? ram_442 : _GEN_11994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11996 = 10'h1bb == _T_29 ? ram_443 : _GEN_11995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11997 = 10'h1bc == _T_29 ? ram_444 : _GEN_11996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11998 = 10'h1bd == _T_29 ? ram_445 : _GEN_11997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_11999 = 10'h1be == _T_29 ? ram_446 : _GEN_11998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12000 = 10'h1bf == _T_29 ? ram_447 : _GEN_11999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12001 = 10'h1c0 == _T_29 ? ram_448 : _GEN_12000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12002 = 10'h1c1 == _T_29 ? ram_449 : _GEN_12001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12003 = 10'h1c2 == _T_29 ? ram_450 : _GEN_12002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12004 = 10'h1c3 == _T_29 ? ram_451 : _GEN_12003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12005 = 10'h1c4 == _T_29 ? ram_452 : _GEN_12004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12006 = 10'h1c5 == _T_29 ? ram_453 : _GEN_12005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12007 = 10'h1c6 == _T_29 ? ram_454 : _GEN_12006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12008 = 10'h1c7 == _T_29 ? ram_455 : _GEN_12007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12009 = 10'h1c8 == _T_29 ? ram_456 : _GEN_12008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12010 = 10'h1c9 == _T_29 ? ram_457 : _GEN_12009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12011 = 10'h1ca == _T_29 ? ram_458 : _GEN_12010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12012 = 10'h1cb == _T_29 ? ram_459 : _GEN_12011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12013 = 10'h1cc == _T_29 ? ram_460 : _GEN_12012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12014 = 10'h1cd == _T_29 ? ram_461 : _GEN_12013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12015 = 10'h1ce == _T_29 ? ram_462 : _GEN_12014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12016 = 10'h1cf == _T_29 ? ram_463 : _GEN_12015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12017 = 10'h1d0 == _T_29 ? ram_464 : _GEN_12016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12018 = 10'h1d1 == _T_29 ? ram_465 : _GEN_12017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12019 = 10'h1d2 == _T_29 ? ram_466 : _GEN_12018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12020 = 10'h1d3 == _T_29 ? ram_467 : _GEN_12019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12021 = 10'h1d4 == _T_29 ? ram_468 : _GEN_12020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12022 = 10'h1d5 == _T_29 ? ram_469 : _GEN_12021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12023 = 10'h1d6 == _T_29 ? ram_470 : _GEN_12022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12024 = 10'h1d7 == _T_29 ? ram_471 : _GEN_12023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12025 = 10'h1d8 == _T_29 ? ram_472 : _GEN_12024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12026 = 10'h1d9 == _T_29 ? ram_473 : _GEN_12025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12027 = 10'h1da == _T_29 ? ram_474 : _GEN_12026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12028 = 10'h1db == _T_29 ? ram_475 : _GEN_12027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12029 = 10'h1dc == _T_29 ? ram_476 : _GEN_12028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12030 = 10'h1dd == _T_29 ? ram_477 : _GEN_12029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12031 = 10'h1de == _T_29 ? ram_478 : _GEN_12030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12032 = 10'h1df == _T_29 ? ram_479 : _GEN_12031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12033 = 10'h1e0 == _T_29 ? ram_480 : _GEN_12032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12034 = 10'h1e1 == _T_29 ? ram_481 : _GEN_12033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12035 = 10'h1e2 == _T_29 ? ram_482 : _GEN_12034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12036 = 10'h1e3 == _T_29 ? ram_483 : _GEN_12035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12037 = 10'h1e4 == _T_29 ? ram_484 : _GEN_12036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12038 = 10'h1e5 == _T_29 ? ram_485 : _GEN_12037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12039 = 10'h1e6 == _T_29 ? ram_486 : _GEN_12038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12040 = 10'h1e7 == _T_29 ? ram_487 : _GEN_12039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12041 = 10'h1e8 == _T_29 ? ram_488 : _GEN_12040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12042 = 10'h1e9 == _T_29 ? ram_489 : _GEN_12041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12043 = 10'h1ea == _T_29 ? ram_490 : _GEN_12042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12044 = 10'h1eb == _T_29 ? ram_491 : _GEN_12043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12045 = 10'h1ec == _T_29 ? ram_492 : _GEN_12044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12046 = 10'h1ed == _T_29 ? ram_493 : _GEN_12045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12047 = 10'h1ee == _T_29 ? ram_494 : _GEN_12046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12048 = 10'h1ef == _T_29 ? ram_495 : _GEN_12047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12049 = 10'h1f0 == _T_29 ? ram_496 : _GEN_12048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12050 = 10'h1f1 == _T_29 ? ram_497 : _GEN_12049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12051 = 10'h1f2 == _T_29 ? ram_498 : _GEN_12050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12052 = 10'h1f3 == _T_29 ? ram_499 : _GEN_12051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12053 = 10'h1f4 == _T_29 ? ram_500 : _GEN_12052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12054 = 10'h1f5 == _T_29 ? ram_501 : _GEN_12053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12055 = 10'h1f6 == _T_29 ? ram_502 : _GEN_12054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12056 = 10'h1f7 == _T_29 ? ram_503 : _GEN_12055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12057 = 10'h1f8 == _T_29 ? ram_504 : _GEN_12056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12058 = 10'h1f9 == _T_29 ? ram_505 : _GEN_12057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12059 = 10'h1fa == _T_29 ? ram_506 : _GEN_12058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12060 = 10'h1fb == _T_29 ? ram_507 : _GEN_12059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12061 = 10'h1fc == _T_29 ? ram_508 : _GEN_12060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12062 = 10'h1fd == _T_29 ? ram_509 : _GEN_12061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12063 = 10'h1fe == _T_29 ? ram_510 : _GEN_12062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12064 = 10'h1ff == _T_29 ? ram_511 : _GEN_12063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12065 = 10'h200 == _T_29 ? ram_512 : _GEN_12064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12066 = 10'h201 == _T_29 ? ram_513 : _GEN_12065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12067 = 10'h202 == _T_29 ? ram_514 : _GEN_12066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12068 = 10'h203 == _T_29 ? ram_515 : _GEN_12067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12069 = 10'h204 == _T_29 ? ram_516 : _GEN_12068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12070 = 10'h205 == _T_29 ? ram_517 : _GEN_12069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12071 = 10'h206 == _T_29 ? ram_518 : _GEN_12070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12072 = 10'h207 == _T_29 ? ram_519 : _GEN_12071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12073 = 10'h208 == _T_29 ? ram_520 : _GEN_12072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12074 = 10'h209 == _T_29 ? ram_521 : _GEN_12073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12075 = 10'h20a == _T_29 ? ram_522 : _GEN_12074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12076 = 10'h20b == _T_29 ? ram_523 : _GEN_12075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12077 = 10'h20c == _T_29 ? ram_524 : _GEN_12076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19083 = {{8190'd0}, _GEN_12077}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_311 = _GEN_19083 ^ _ram_T_310; // @[vga.scala 64:41]
  wire [287:0] _GEN_12078 = 10'h0 == _T_29 ? _ram_T_311[287:0] : _GEN_11028; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12079 = 10'h1 == _T_29 ? _ram_T_311[287:0] : _GEN_11029; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12080 = 10'h2 == _T_29 ? _ram_T_311[287:0] : _GEN_11030; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12081 = 10'h3 == _T_29 ? _ram_T_311[287:0] : _GEN_11031; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12082 = 10'h4 == _T_29 ? _ram_T_311[287:0] : _GEN_11032; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12083 = 10'h5 == _T_29 ? _ram_T_311[287:0] : _GEN_11033; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12084 = 10'h6 == _T_29 ? _ram_T_311[287:0] : _GEN_11034; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12085 = 10'h7 == _T_29 ? _ram_T_311[287:0] : _GEN_11035; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12086 = 10'h8 == _T_29 ? _ram_T_311[287:0] : _GEN_11036; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12087 = 10'h9 == _T_29 ? _ram_T_311[287:0] : _GEN_11037; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12088 = 10'ha == _T_29 ? _ram_T_311[287:0] : _GEN_11038; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12089 = 10'hb == _T_29 ? _ram_T_311[287:0] : _GEN_11039; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12090 = 10'hc == _T_29 ? _ram_T_311[287:0] : _GEN_11040; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12091 = 10'hd == _T_29 ? _ram_T_311[287:0] : _GEN_11041; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12092 = 10'he == _T_29 ? _ram_T_311[287:0] : _GEN_11042; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12093 = 10'hf == _T_29 ? _ram_T_311[287:0] : _GEN_11043; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12094 = 10'h10 == _T_29 ? _ram_T_311[287:0] : _GEN_11044; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12095 = 10'h11 == _T_29 ? _ram_T_311[287:0] : _GEN_11045; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12096 = 10'h12 == _T_29 ? _ram_T_311[287:0] : _GEN_11046; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12097 = 10'h13 == _T_29 ? _ram_T_311[287:0] : _GEN_11047; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12098 = 10'h14 == _T_29 ? _ram_T_311[287:0] : _GEN_11048; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12099 = 10'h15 == _T_29 ? _ram_T_311[287:0] : _GEN_11049; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12100 = 10'h16 == _T_29 ? _ram_T_311[287:0] : _GEN_11050; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12101 = 10'h17 == _T_29 ? _ram_T_311[287:0] : _GEN_11051; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12102 = 10'h18 == _T_29 ? _ram_T_311[287:0] : _GEN_11052; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12103 = 10'h19 == _T_29 ? _ram_T_311[287:0] : _GEN_11053; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12104 = 10'h1a == _T_29 ? _ram_T_311[287:0] : _GEN_11054; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12105 = 10'h1b == _T_29 ? _ram_T_311[287:0] : _GEN_11055; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12106 = 10'h1c == _T_29 ? _ram_T_311[287:0] : _GEN_11056; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12107 = 10'h1d == _T_29 ? _ram_T_311[287:0] : _GEN_11057; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12108 = 10'h1e == _T_29 ? _ram_T_311[287:0] : _GEN_11058; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12109 = 10'h1f == _T_29 ? _ram_T_311[287:0] : _GEN_11059; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12110 = 10'h20 == _T_29 ? _ram_T_311[287:0] : _GEN_11060; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12111 = 10'h21 == _T_29 ? _ram_T_311[287:0] : _GEN_11061; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12112 = 10'h22 == _T_29 ? _ram_T_311[287:0] : _GEN_11062; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12113 = 10'h23 == _T_29 ? _ram_T_311[287:0] : _GEN_11063; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12114 = 10'h24 == _T_29 ? _ram_T_311[287:0] : _GEN_11064; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12115 = 10'h25 == _T_29 ? _ram_T_311[287:0] : _GEN_11065; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12116 = 10'h26 == _T_29 ? _ram_T_311[287:0] : _GEN_11066; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12117 = 10'h27 == _T_29 ? _ram_T_311[287:0] : _GEN_11067; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12118 = 10'h28 == _T_29 ? _ram_T_311[287:0] : _GEN_11068; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12119 = 10'h29 == _T_29 ? _ram_T_311[287:0] : _GEN_11069; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12120 = 10'h2a == _T_29 ? _ram_T_311[287:0] : _GEN_11070; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12121 = 10'h2b == _T_29 ? _ram_T_311[287:0] : _GEN_11071; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12122 = 10'h2c == _T_29 ? _ram_T_311[287:0] : _GEN_11072; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12123 = 10'h2d == _T_29 ? _ram_T_311[287:0] : _GEN_11073; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12124 = 10'h2e == _T_29 ? _ram_T_311[287:0] : _GEN_11074; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12125 = 10'h2f == _T_29 ? _ram_T_311[287:0] : _GEN_11075; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12126 = 10'h30 == _T_29 ? _ram_T_311[287:0] : _GEN_11076; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12127 = 10'h31 == _T_29 ? _ram_T_311[287:0] : _GEN_11077; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12128 = 10'h32 == _T_29 ? _ram_T_311[287:0] : _GEN_11078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12129 = 10'h33 == _T_29 ? _ram_T_311[287:0] : _GEN_11079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12130 = 10'h34 == _T_29 ? _ram_T_311[287:0] : _GEN_11080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12131 = 10'h35 == _T_29 ? _ram_T_311[287:0] : _GEN_11081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12132 = 10'h36 == _T_29 ? _ram_T_311[287:0] : _GEN_11082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12133 = 10'h37 == _T_29 ? _ram_T_311[287:0] : _GEN_11083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12134 = 10'h38 == _T_29 ? _ram_T_311[287:0] : _GEN_11084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12135 = 10'h39 == _T_29 ? _ram_T_311[287:0] : _GEN_11085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12136 = 10'h3a == _T_29 ? _ram_T_311[287:0] : _GEN_11086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12137 = 10'h3b == _T_29 ? _ram_T_311[287:0] : _GEN_11087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12138 = 10'h3c == _T_29 ? _ram_T_311[287:0] : _GEN_11088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12139 = 10'h3d == _T_29 ? _ram_T_311[287:0] : _GEN_11089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12140 = 10'h3e == _T_29 ? _ram_T_311[287:0] : _GEN_11090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12141 = 10'h3f == _T_29 ? _ram_T_311[287:0] : _GEN_11091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12142 = 10'h40 == _T_29 ? _ram_T_311[287:0] : _GEN_11092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12143 = 10'h41 == _T_29 ? _ram_T_311[287:0] : _GEN_11093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12144 = 10'h42 == _T_29 ? _ram_T_311[287:0] : _GEN_11094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12145 = 10'h43 == _T_29 ? _ram_T_311[287:0] : _GEN_11095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12146 = 10'h44 == _T_29 ? _ram_T_311[287:0] : _GEN_11096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12147 = 10'h45 == _T_29 ? _ram_T_311[287:0] : _GEN_11097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12148 = 10'h46 == _T_29 ? _ram_T_311[287:0] : _GEN_11098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12149 = 10'h47 == _T_29 ? _ram_T_311[287:0] : _GEN_11099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12150 = 10'h48 == _T_29 ? _ram_T_311[287:0] : _GEN_11100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12151 = 10'h49 == _T_29 ? _ram_T_311[287:0] : _GEN_11101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12152 = 10'h4a == _T_29 ? _ram_T_311[287:0] : _GEN_11102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12153 = 10'h4b == _T_29 ? _ram_T_311[287:0] : _GEN_11103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12154 = 10'h4c == _T_29 ? _ram_T_311[287:0] : _GEN_11104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12155 = 10'h4d == _T_29 ? _ram_T_311[287:0] : _GEN_11105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12156 = 10'h4e == _T_29 ? _ram_T_311[287:0] : _GEN_11106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12157 = 10'h4f == _T_29 ? _ram_T_311[287:0] : _GEN_11107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12158 = 10'h50 == _T_29 ? _ram_T_311[287:0] : _GEN_11108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12159 = 10'h51 == _T_29 ? _ram_T_311[287:0] : _GEN_11109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12160 = 10'h52 == _T_29 ? _ram_T_311[287:0] : _GEN_11110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12161 = 10'h53 == _T_29 ? _ram_T_311[287:0] : _GEN_11111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12162 = 10'h54 == _T_29 ? _ram_T_311[287:0] : _GEN_11112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12163 = 10'h55 == _T_29 ? _ram_T_311[287:0] : _GEN_11113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12164 = 10'h56 == _T_29 ? _ram_T_311[287:0] : _GEN_11114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12165 = 10'h57 == _T_29 ? _ram_T_311[287:0] : _GEN_11115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12166 = 10'h58 == _T_29 ? _ram_T_311[287:0] : _GEN_11116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12167 = 10'h59 == _T_29 ? _ram_T_311[287:0] : _GEN_11117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12168 = 10'h5a == _T_29 ? _ram_T_311[287:0] : _GEN_11118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12169 = 10'h5b == _T_29 ? _ram_T_311[287:0] : _GEN_11119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12170 = 10'h5c == _T_29 ? _ram_T_311[287:0] : _GEN_11120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12171 = 10'h5d == _T_29 ? _ram_T_311[287:0] : _GEN_11121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12172 = 10'h5e == _T_29 ? _ram_T_311[287:0] : _GEN_11122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12173 = 10'h5f == _T_29 ? _ram_T_311[287:0] : _GEN_11123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12174 = 10'h60 == _T_29 ? _ram_T_311[287:0] : _GEN_11124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12175 = 10'h61 == _T_29 ? _ram_T_311[287:0] : _GEN_11125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12176 = 10'h62 == _T_29 ? _ram_T_311[287:0] : _GEN_11126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12177 = 10'h63 == _T_29 ? _ram_T_311[287:0] : _GEN_11127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12178 = 10'h64 == _T_29 ? _ram_T_311[287:0] : _GEN_11128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12179 = 10'h65 == _T_29 ? _ram_T_311[287:0] : _GEN_11129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12180 = 10'h66 == _T_29 ? _ram_T_311[287:0] : _GEN_11130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12181 = 10'h67 == _T_29 ? _ram_T_311[287:0] : _GEN_11131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12182 = 10'h68 == _T_29 ? _ram_T_311[287:0] : _GEN_11132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12183 = 10'h69 == _T_29 ? _ram_T_311[287:0] : _GEN_11133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12184 = 10'h6a == _T_29 ? _ram_T_311[287:0] : _GEN_11134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12185 = 10'h6b == _T_29 ? _ram_T_311[287:0] : _GEN_11135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12186 = 10'h6c == _T_29 ? _ram_T_311[287:0] : _GEN_11136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12187 = 10'h6d == _T_29 ? _ram_T_311[287:0] : _GEN_11137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12188 = 10'h6e == _T_29 ? _ram_T_311[287:0] : _GEN_11138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12189 = 10'h6f == _T_29 ? _ram_T_311[287:0] : _GEN_11139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12190 = 10'h70 == _T_29 ? _ram_T_311[287:0] : _GEN_11140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12191 = 10'h71 == _T_29 ? _ram_T_311[287:0] : _GEN_11141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12192 = 10'h72 == _T_29 ? _ram_T_311[287:0] : _GEN_11142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12193 = 10'h73 == _T_29 ? _ram_T_311[287:0] : _GEN_11143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12194 = 10'h74 == _T_29 ? _ram_T_311[287:0] : _GEN_11144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12195 = 10'h75 == _T_29 ? _ram_T_311[287:0] : _GEN_11145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12196 = 10'h76 == _T_29 ? _ram_T_311[287:0] : _GEN_11146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12197 = 10'h77 == _T_29 ? _ram_T_311[287:0] : _GEN_11147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12198 = 10'h78 == _T_29 ? _ram_T_311[287:0] : _GEN_11148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12199 = 10'h79 == _T_29 ? _ram_T_311[287:0] : _GEN_11149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12200 = 10'h7a == _T_29 ? _ram_T_311[287:0] : _GEN_11150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12201 = 10'h7b == _T_29 ? _ram_T_311[287:0] : _GEN_11151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12202 = 10'h7c == _T_29 ? _ram_T_311[287:0] : _GEN_11152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12203 = 10'h7d == _T_29 ? _ram_T_311[287:0] : _GEN_11153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12204 = 10'h7e == _T_29 ? _ram_T_311[287:0] : _GEN_11154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12205 = 10'h7f == _T_29 ? _ram_T_311[287:0] : _GEN_11155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12206 = 10'h80 == _T_29 ? _ram_T_311[287:0] : _GEN_11156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12207 = 10'h81 == _T_29 ? _ram_T_311[287:0] : _GEN_11157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12208 = 10'h82 == _T_29 ? _ram_T_311[287:0] : _GEN_11158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12209 = 10'h83 == _T_29 ? _ram_T_311[287:0] : _GEN_11159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12210 = 10'h84 == _T_29 ? _ram_T_311[287:0] : _GEN_11160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12211 = 10'h85 == _T_29 ? _ram_T_311[287:0] : _GEN_11161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12212 = 10'h86 == _T_29 ? _ram_T_311[287:0] : _GEN_11162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12213 = 10'h87 == _T_29 ? _ram_T_311[287:0] : _GEN_11163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12214 = 10'h88 == _T_29 ? _ram_T_311[287:0] : _GEN_11164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12215 = 10'h89 == _T_29 ? _ram_T_311[287:0] : _GEN_11165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12216 = 10'h8a == _T_29 ? _ram_T_311[287:0] : _GEN_11166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12217 = 10'h8b == _T_29 ? _ram_T_311[287:0] : _GEN_11167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12218 = 10'h8c == _T_29 ? _ram_T_311[287:0] : _GEN_11168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12219 = 10'h8d == _T_29 ? _ram_T_311[287:0] : _GEN_11169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12220 = 10'h8e == _T_29 ? _ram_T_311[287:0] : _GEN_11170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12221 = 10'h8f == _T_29 ? _ram_T_311[287:0] : _GEN_11171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12222 = 10'h90 == _T_29 ? _ram_T_311[287:0] : _GEN_11172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12223 = 10'h91 == _T_29 ? _ram_T_311[287:0] : _GEN_11173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12224 = 10'h92 == _T_29 ? _ram_T_311[287:0] : _GEN_11174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12225 = 10'h93 == _T_29 ? _ram_T_311[287:0] : _GEN_11175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12226 = 10'h94 == _T_29 ? _ram_T_311[287:0] : _GEN_11176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12227 = 10'h95 == _T_29 ? _ram_T_311[287:0] : _GEN_11177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12228 = 10'h96 == _T_29 ? _ram_T_311[287:0] : _GEN_11178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12229 = 10'h97 == _T_29 ? _ram_T_311[287:0] : _GEN_11179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12230 = 10'h98 == _T_29 ? _ram_T_311[287:0] : _GEN_11180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12231 = 10'h99 == _T_29 ? _ram_T_311[287:0] : _GEN_11181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12232 = 10'h9a == _T_29 ? _ram_T_311[287:0] : _GEN_11182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12233 = 10'h9b == _T_29 ? _ram_T_311[287:0] : _GEN_11183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12234 = 10'h9c == _T_29 ? _ram_T_311[287:0] : _GEN_11184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12235 = 10'h9d == _T_29 ? _ram_T_311[287:0] : _GEN_11185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12236 = 10'h9e == _T_29 ? _ram_T_311[287:0] : _GEN_11186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12237 = 10'h9f == _T_29 ? _ram_T_311[287:0] : _GEN_11187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12238 = 10'ha0 == _T_29 ? _ram_T_311[287:0] : _GEN_11188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12239 = 10'ha1 == _T_29 ? _ram_T_311[287:0] : _GEN_11189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12240 = 10'ha2 == _T_29 ? _ram_T_311[287:0] : _GEN_11190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12241 = 10'ha3 == _T_29 ? _ram_T_311[287:0] : _GEN_11191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12242 = 10'ha4 == _T_29 ? _ram_T_311[287:0] : _GEN_11192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12243 = 10'ha5 == _T_29 ? _ram_T_311[287:0] : _GEN_11193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12244 = 10'ha6 == _T_29 ? _ram_T_311[287:0] : _GEN_11194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12245 = 10'ha7 == _T_29 ? _ram_T_311[287:0] : _GEN_11195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12246 = 10'ha8 == _T_29 ? _ram_T_311[287:0] : _GEN_11196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12247 = 10'ha9 == _T_29 ? _ram_T_311[287:0] : _GEN_11197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12248 = 10'haa == _T_29 ? _ram_T_311[287:0] : _GEN_11198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12249 = 10'hab == _T_29 ? _ram_T_311[287:0] : _GEN_11199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12250 = 10'hac == _T_29 ? _ram_T_311[287:0] : _GEN_11200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12251 = 10'had == _T_29 ? _ram_T_311[287:0] : _GEN_11201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12252 = 10'hae == _T_29 ? _ram_T_311[287:0] : _GEN_11202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12253 = 10'haf == _T_29 ? _ram_T_311[287:0] : _GEN_11203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12254 = 10'hb0 == _T_29 ? _ram_T_311[287:0] : _GEN_11204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12255 = 10'hb1 == _T_29 ? _ram_T_311[287:0] : _GEN_11205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12256 = 10'hb2 == _T_29 ? _ram_T_311[287:0] : _GEN_11206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12257 = 10'hb3 == _T_29 ? _ram_T_311[287:0] : _GEN_11207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12258 = 10'hb4 == _T_29 ? _ram_T_311[287:0] : _GEN_11208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12259 = 10'hb5 == _T_29 ? _ram_T_311[287:0] : _GEN_11209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12260 = 10'hb6 == _T_29 ? _ram_T_311[287:0] : _GEN_11210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12261 = 10'hb7 == _T_29 ? _ram_T_311[287:0] : _GEN_11211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12262 = 10'hb8 == _T_29 ? _ram_T_311[287:0] : _GEN_11212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12263 = 10'hb9 == _T_29 ? _ram_T_311[287:0] : _GEN_11213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12264 = 10'hba == _T_29 ? _ram_T_311[287:0] : _GEN_11214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12265 = 10'hbb == _T_29 ? _ram_T_311[287:0] : _GEN_11215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12266 = 10'hbc == _T_29 ? _ram_T_311[287:0] : _GEN_11216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12267 = 10'hbd == _T_29 ? _ram_T_311[287:0] : _GEN_11217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12268 = 10'hbe == _T_29 ? _ram_T_311[287:0] : _GEN_11218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12269 = 10'hbf == _T_29 ? _ram_T_311[287:0] : _GEN_11219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12270 = 10'hc0 == _T_29 ? _ram_T_311[287:0] : _GEN_11220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12271 = 10'hc1 == _T_29 ? _ram_T_311[287:0] : _GEN_11221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12272 = 10'hc2 == _T_29 ? _ram_T_311[287:0] : _GEN_11222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12273 = 10'hc3 == _T_29 ? _ram_T_311[287:0] : _GEN_11223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12274 = 10'hc4 == _T_29 ? _ram_T_311[287:0] : _GEN_11224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12275 = 10'hc5 == _T_29 ? _ram_T_311[287:0] : _GEN_11225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12276 = 10'hc6 == _T_29 ? _ram_T_311[287:0] : _GEN_11226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12277 = 10'hc7 == _T_29 ? _ram_T_311[287:0] : _GEN_11227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12278 = 10'hc8 == _T_29 ? _ram_T_311[287:0] : _GEN_11228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12279 = 10'hc9 == _T_29 ? _ram_T_311[287:0] : _GEN_11229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12280 = 10'hca == _T_29 ? _ram_T_311[287:0] : _GEN_11230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12281 = 10'hcb == _T_29 ? _ram_T_311[287:0] : _GEN_11231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12282 = 10'hcc == _T_29 ? _ram_T_311[287:0] : _GEN_11232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12283 = 10'hcd == _T_29 ? _ram_T_311[287:0] : _GEN_11233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12284 = 10'hce == _T_29 ? _ram_T_311[287:0] : _GEN_11234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12285 = 10'hcf == _T_29 ? _ram_T_311[287:0] : _GEN_11235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12286 = 10'hd0 == _T_29 ? _ram_T_311[287:0] : _GEN_11236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12287 = 10'hd1 == _T_29 ? _ram_T_311[287:0] : _GEN_11237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12288 = 10'hd2 == _T_29 ? _ram_T_311[287:0] : _GEN_11238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12289 = 10'hd3 == _T_29 ? _ram_T_311[287:0] : _GEN_11239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12290 = 10'hd4 == _T_29 ? _ram_T_311[287:0] : _GEN_11240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12291 = 10'hd5 == _T_29 ? _ram_T_311[287:0] : _GEN_11241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12292 = 10'hd6 == _T_29 ? _ram_T_311[287:0] : _GEN_11242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12293 = 10'hd7 == _T_29 ? _ram_T_311[287:0] : _GEN_11243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12294 = 10'hd8 == _T_29 ? _ram_T_311[287:0] : _GEN_11244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12295 = 10'hd9 == _T_29 ? _ram_T_311[287:0] : _GEN_11245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12296 = 10'hda == _T_29 ? _ram_T_311[287:0] : _GEN_11246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12297 = 10'hdb == _T_29 ? _ram_T_311[287:0] : _GEN_11247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12298 = 10'hdc == _T_29 ? _ram_T_311[287:0] : _GEN_11248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12299 = 10'hdd == _T_29 ? _ram_T_311[287:0] : _GEN_11249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12300 = 10'hde == _T_29 ? _ram_T_311[287:0] : _GEN_11250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12301 = 10'hdf == _T_29 ? _ram_T_311[287:0] : _GEN_11251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12302 = 10'he0 == _T_29 ? _ram_T_311[287:0] : _GEN_11252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12303 = 10'he1 == _T_29 ? _ram_T_311[287:0] : _GEN_11253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12304 = 10'he2 == _T_29 ? _ram_T_311[287:0] : _GEN_11254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12305 = 10'he3 == _T_29 ? _ram_T_311[287:0] : _GEN_11255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12306 = 10'he4 == _T_29 ? _ram_T_311[287:0] : _GEN_11256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12307 = 10'he5 == _T_29 ? _ram_T_311[287:0] : _GEN_11257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12308 = 10'he6 == _T_29 ? _ram_T_311[287:0] : _GEN_11258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12309 = 10'he7 == _T_29 ? _ram_T_311[287:0] : _GEN_11259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12310 = 10'he8 == _T_29 ? _ram_T_311[287:0] : _GEN_11260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12311 = 10'he9 == _T_29 ? _ram_T_311[287:0] : _GEN_11261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12312 = 10'hea == _T_29 ? _ram_T_311[287:0] : _GEN_11262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12313 = 10'heb == _T_29 ? _ram_T_311[287:0] : _GEN_11263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12314 = 10'hec == _T_29 ? _ram_T_311[287:0] : _GEN_11264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12315 = 10'hed == _T_29 ? _ram_T_311[287:0] : _GEN_11265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12316 = 10'hee == _T_29 ? _ram_T_311[287:0] : _GEN_11266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12317 = 10'hef == _T_29 ? _ram_T_311[287:0] : _GEN_11267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12318 = 10'hf0 == _T_29 ? _ram_T_311[287:0] : _GEN_11268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12319 = 10'hf1 == _T_29 ? _ram_T_311[287:0] : _GEN_11269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12320 = 10'hf2 == _T_29 ? _ram_T_311[287:0] : _GEN_11270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12321 = 10'hf3 == _T_29 ? _ram_T_311[287:0] : _GEN_11271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12322 = 10'hf4 == _T_29 ? _ram_T_311[287:0] : _GEN_11272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12323 = 10'hf5 == _T_29 ? _ram_T_311[287:0] : _GEN_11273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12324 = 10'hf6 == _T_29 ? _ram_T_311[287:0] : _GEN_11274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12325 = 10'hf7 == _T_29 ? _ram_T_311[287:0] : _GEN_11275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12326 = 10'hf8 == _T_29 ? _ram_T_311[287:0] : _GEN_11276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12327 = 10'hf9 == _T_29 ? _ram_T_311[287:0] : _GEN_11277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12328 = 10'hfa == _T_29 ? _ram_T_311[287:0] : _GEN_11278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12329 = 10'hfb == _T_29 ? _ram_T_311[287:0] : _GEN_11279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12330 = 10'hfc == _T_29 ? _ram_T_311[287:0] : _GEN_11280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12331 = 10'hfd == _T_29 ? _ram_T_311[287:0] : _GEN_11281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12332 = 10'hfe == _T_29 ? _ram_T_311[287:0] : _GEN_11282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12333 = 10'hff == _T_29 ? _ram_T_311[287:0] : _GEN_11283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12334 = 10'h100 == _T_29 ? _ram_T_311[287:0] : _GEN_11284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12335 = 10'h101 == _T_29 ? _ram_T_311[287:0] : _GEN_11285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12336 = 10'h102 == _T_29 ? _ram_T_311[287:0] : _GEN_11286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12337 = 10'h103 == _T_29 ? _ram_T_311[287:0] : _GEN_11287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12338 = 10'h104 == _T_29 ? _ram_T_311[287:0] : _GEN_11288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12339 = 10'h105 == _T_29 ? _ram_T_311[287:0] : _GEN_11289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12340 = 10'h106 == _T_29 ? _ram_T_311[287:0] : _GEN_11290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12341 = 10'h107 == _T_29 ? _ram_T_311[287:0] : _GEN_11291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12342 = 10'h108 == _T_29 ? _ram_T_311[287:0] : _GEN_11292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12343 = 10'h109 == _T_29 ? _ram_T_311[287:0] : _GEN_11293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12344 = 10'h10a == _T_29 ? _ram_T_311[287:0] : _GEN_11294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12345 = 10'h10b == _T_29 ? _ram_T_311[287:0] : _GEN_11295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12346 = 10'h10c == _T_29 ? _ram_T_311[287:0] : _GEN_11296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12347 = 10'h10d == _T_29 ? _ram_T_311[287:0] : _GEN_11297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12348 = 10'h10e == _T_29 ? _ram_T_311[287:0] : _GEN_11298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12349 = 10'h10f == _T_29 ? _ram_T_311[287:0] : _GEN_11299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12350 = 10'h110 == _T_29 ? _ram_T_311[287:0] : _GEN_11300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12351 = 10'h111 == _T_29 ? _ram_T_311[287:0] : _GEN_11301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12352 = 10'h112 == _T_29 ? _ram_T_311[287:0] : _GEN_11302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12353 = 10'h113 == _T_29 ? _ram_T_311[287:0] : _GEN_11303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12354 = 10'h114 == _T_29 ? _ram_T_311[287:0] : _GEN_11304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12355 = 10'h115 == _T_29 ? _ram_T_311[287:0] : _GEN_11305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12356 = 10'h116 == _T_29 ? _ram_T_311[287:0] : _GEN_11306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12357 = 10'h117 == _T_29 ? _ram_T_311[287:0] : _GEN_11307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12358 = 10'h118 == _T_29 ? _ram_T_311[287:0] : _GEN_11308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12359 = 10'h119 == _T_29 ? _ram_T_311[287:0] : _GEN_11309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12360 = 10'h11a == _T_29 ? _ram_T_311[287:0] : _GEN_11310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12361 = 10'h11b == _T_29 ? _ram_T_311[287:0] : _GEN_11311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12362 = 10'h11c == _T_29 ? _ram_T_311[287:0] : _GEN_11312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12363 = 10'h11d == _T_29 ? _ram_T_311[287:0] : _GEN_11313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12364 = 10'h11e == _T_29 ? _ram_T_311[287:0] : _GEN_11314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12365 = 10'h11f == _T_29 ? _ram_T_311[287:0] : _GEN_11315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12366 = 10'h120 == _T_29 ? _ram_T_311[287:0] : _GEN_11316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12367 = 10'h121 == _T_29 ? _ram_T_311[287:0] : _GEN_11317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12368 = 10'h122 == _T_29 ? _ram_T_311[287:0] : _GEN_11318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12369 = 10'h123 == _T_29 ? _ram_T_311[287:0] : _GEN_11319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12370 = 10'h124 == _T_29 ? _ram_T_311[287:0] : _GEN_11320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12371 = 10'h125 == _T_29 ? _ram_T_311[287:0] : _GEN_11321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12372 = 10'h126 == _T_29 ? _ram_T_311[287:0] : _GEN_11322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12373 = 10'h127 == _T_29 ? _ram_T_311[287:0] : _GEN_11323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12374 = 10'h128 == _T_29 ? _ram_T_311[287:0] : _GEN_11324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12375 = 10'h129 == _T_29 ? _ram_T_311[287:0] : _GEN_11325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12376 = 10'h12a == _T_29 ? _ram_T_311[287:0] : _GEN_11326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12377 = 10'h12b == _T_29 ? _ram_T_311[287:0] : _GEN_11327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12378 = 10'h12c == _T_29 ? _ram_T_311[287:0] : _GEN_11328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12379 = 10'h12d == _T_29 ? _ram_T_311[287:0] : _GEN_11329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12380 = 10'h12e == _T_29 ? _ram_T_311[287:0] : _GEN_11330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12381 = 10'h12f == _T_29 ? _ram_T_311[287:0] : _GEN_11331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12382 = 10'h130 == _T_29 ? _ram_T_311[287:0] : _GEN_11332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12383 = 10'h131 == _T_29 ? _ram_T_311[287:0] : _GEN_11333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12384 = 10'h132 == _T_29 ? _ram_T_311[287:0] : _GEN_11334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12385 = 10'h133 == _T_29 ? _ram_T_311[287:0] : _GEN_11335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12386 = 10'h134 == _T_29 ? _ram_T_311[287:0] : _GEN_11336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12387 = 10'h135 == _T_29 ? _ram_T_311[287:0] : _GEN_11337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12388 = 10'h136 == _T_29 ? _ram_T_311[287:0] : _GEN_11338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12389 = 10'h137 == _T_29 ? _ram_T_311[287:0] : _GEN_11339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12390 = 10'h138 == _T_29 ? _ram_T_311[287:0] : _GEN_11340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12391 = 10'h139 == _T_29 ? _ram_T_311[287:0] : _GEN_11341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12392 = 10'h13a == _T_29 ? _ram_T_311[287:0] : _GEN_11342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12393 = 10'h13b == _T_29 ? _ram_T_311[287:0] : _GEN_11343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12394 = 10'h13c == _T_29 ? _ram_T_311[287:0] : _GEN_11344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12395 = 10'h13d == _T_29 ? _ram_T_311[287:0] : _GEN_11345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12396 = 10'h13e == _T_29 ? _ram_T_311[287:0] : _GEN_11346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12397 = 10'h13f == _T_29 ? _ram_T_311[287:0] : _GEN_11347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12398 = 10'h140 == _T_29 ? _ram_T_311[287:0] : _GEN_11348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12399 = 10'h141 == _T_29 ? _ram_T_311[287:0] : _GEN_11349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12400 = 10'h142 == _T_29 ? _ram_T_311[287:0] : _GEN_11350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12401 = 10'h143 == _T_29 ? _ram_T_311[287:0] : _GEN_11351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12402 = 10'h144 == _T_29 ? _ram_T_311[287:0] : _GEN_11352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12403 = 10'h145 == _T_29 ? _ram_T_311[287:0] : _GEN_11353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12404 = 10'h146 == _T_29 ? _ram_T_311[287:0] : _GEN_11354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12405 = 10'h147 == _T_29 ? _ram_T_311[287:0] : _GEN_11355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12406 = 10'h148 == _T_29 ? _ram_T_311[287:0] : _GEN_11356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12407 = 10'h149 == _T_29 ? _ram_T_311[287:0] : _GEN_11357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12408 = 10'h14a == _T_29 ? _ram_T_311[287:0] : _GEN_11358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12409 = 10'h14b == _T_29 ? _ram_T_311[287:0] : _GEN_11359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12410 = 10'h14c == _T_29 ? _ram_T_311[287:0] : _GEN_11360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12411 = 10'h14d == _T_29 ? _ram_T_311[287:0] : _GEN_11361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12412 = 10'h14e == _T_29 ? _ram_T_311[287:0] : _GEN_11362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12413 = 10'h14f == _T_29 ? _ram_T_311[287:0] : _GEN_11363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12414 = 10'h150 == _T_29 ? _ram_T_311[287:0] : _GEN_11364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12415 = 10'h151 == _T_29 ? _ram_T_311[287:0] : _GEN_11365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12416 = 10'h152 == _T_29 ? _ram_T_311[287:0] : _GEN_11366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12417 = 10'h153 == _T_29 ? _ram_T_311[287:0] : _GEN_11367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12418 = 10'h154 == _T_29 ? _ram_T_311[287:0] : _GEN_11368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12419 = 10'h155 == _T_29 ? _ram_T_311[287:0] : _GEN_11369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12420 = 10'h156 == _T_29 ? _ram_T_311[287:0] : _GEN_11370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12421 = 10'h157 == _T_29 ? _ram_T_311[287:0] : _GEN_11371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12422 = 10'h158 == _T_29 ? _ram_T_311[287:0] : _GEN_11372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12423 = 10'h159 == _T_29 ? _ram_T_311[287:0] : _GEN_11373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12424 = 10'h15a == _T_29 ? _ram_T_311[287:0] : _GEN_11374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12425 = 10'h15b == _T_29 ? _ram_T_311[287:0] : _GEN_11375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12426 = 10'h15c == _T_29 ? _ram_T_311[287:0] : _GEN_11376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12427 = 10'h15d == _T_29 ? _ram_T_311[287:0] : _GEN_11377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12428 = 10'h15e == _T_29 ? _ram_T_311[287:0] : _GEN_11378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12429 = 10'h15f == _T_29 ? _ram_T_311[287:0] : _GEN_11379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12430 = 10'h160 == _T_29 ? _ram_T_311[287:0] : _GEN_11380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12431 = 10'h161 == _T_29 ? _ram_T_311[287:0] : _GEN_11381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12432 = 10'h162 == _T_29 ? _ram_T_311[287:0] : _GEN_11382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12433 = 10'h163 == _T_29 ? _ram_T_311[287:0] : _GEN_11383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12434 = 10'h164 == _T_29 ? _ram_T_311[287:0] : _GEN_11384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12435 = 10'h165 == _T_29 ? _ram_T_311[287:0] : _GEN_11385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12436 = 10'h166 == _T_29 ? _ram_T_311[287:0] : _GEN_11386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12437 = 10'h167 == _T_29 ? _ram_T_311[287:0] : _GEN_11387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12438 = 10'h168 == _T_29 ? _ram_T_311[287:0] : _GEN_11388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12439 = 10'h169 == _T_29 ? _ram_T_311[287:0] : _GEN_11389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12440 = 10'h16a == _T_29 ? _ram_T_311[287:0] : _GEN_11390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12441 = 10'h16b == _T_29 ? _ram_T_311[287:0] : _GEN_11391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12442 = 10'h16c == _T_29 ? _ram_T_311[287:0] : _GEN_11392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12443 = 10'h16d == _T_29 ? _ram_T_311[287:0] : _GEN_11393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12444 = 10'h16e == _T_29 ? _ram_T_311[287:0] : _GEN_11394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12445 = 10'h16f == _T_29 ? _ram_T_311[287:0] : _GEN_11395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12446 = 10'h170 == _T_29 ? _ram_T_311[287:0] : _GEN_11396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12447 = 10'h171 == _T_29 ? _ram_T_311[287:0] : _GEN_11397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12448 = 10'h172 == _T_29 ? _ram_T_311[287:0] : _GEN_11398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12449 = 10'h173 == _T_29 ? _ram_T_311[287:0] : _GEN_11399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12450 = 10'h174 == _T_29 ? _ram_T_311[287:0] : _GEN_11400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12451 = 10'h175 == _T_29 ? _ram_T_311[287:0] : _GEN_11401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12452 = 10'h176 == _T_29 ? _ram_T_311[287:0] : _GEN_11402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12453 = 10'h177 == _T_29 ? _ram_T_311[287:0] : _GEN_11403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12454 = 10'h178 == _T_29 ? _ram_T_311[287:0] : _GEN_11404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12455 = 10'h179 == _T_29 ? _ram_T_311[287:0] : _GEN_11405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12456 = 10'h17a == _T_29 ? _ram_T_311[287:0] : _GEN_11406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12457 = 10'h17b == _T_29 ? _ram_T_311[287:0] : _GEN_11407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12458 = 10'h17c == _T_29 ? _ram_T_311[287:0] : _GEN_11408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12459 = 10'h17d == _T_29 ? _ram_T_311[287:0] : _GEN_11409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12460 = 10'h17e == _T_29 ? _ram_T_311[287:0] : _GEN_11410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12461 = 10'h17f == _T_29 ? _ram_T_311[287:0] : _GEN_11411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12462 = 10'h180 == _T_29 ? _ram_T_311[287:0] : _GEN_11412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12463 = 10'h181 == _T_29 ? _ram_T_311[287:0] : _GEN_11413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12464 = 10'h182 == _T_29 ? _ram_T_311[287:0] : _GEN_11414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12465 = 10'h183 == _T_29 ? _ram_T_311[287:0] : _GEN_11415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12466 = 10'h184 == _T_29 ? _ram_T_311[287:0] : _GEN_11416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12467 = 10'h185 == _T_29 ? _ram_T_311[287:0] : _GEN_11417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12468 = 10'h186 == _T_29 ? _ram_T_311[287:0] : _GEN_11418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12469 = 10'h187 == _T_29 ? _ram_T_311[287:0] : _GEN_11419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12470 = 10'h188 == _T_29 ? _ram_T_311[287:0] : _GEN_11420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12471 = 10'h189 == _T_29 ? _ram_T_311[287:0] : _GEN_11421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12472 = 10'h18a == _T_29 ? _ram_T_311[287:0] : _GEN_11422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12473 = 10'h18b == _T_29 ? _ram_T_311[287:0] : _GEN_11423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12474 = 10'h18c == _T_29 ? _ram_T_311[287:0] : _GEN_11424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12475 = 10'h18d == _T_29 ? _ram_T_311[287:0] : _GEN_11425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12476 = 10'h18e == _T_29 ? _ram_T_311[287:0] : _GEN_11426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12477 = 10'h18f == _T_29 ? _ram_T_311[287:0] : _GEN_11427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12478 = 10'h190 == _T_29 ? _ram_T_311[287:0] : _GEN_11428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12479 = 10'h191 == _T_29 ? _ram_T_311[287:0] : _GEN_11429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12480 = 10'h192 == _T_29 ? _ram_T_311[287:0] : _GEN_11430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12481 = 10'h193 == _T_29 ? _ram_T_311[287:0] : _GEN_11431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12482 = 10'h194 == _T_29 ? _ram_T_311[287:0] : _GEN_11432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12483 = 10'h195 == _T_29 ? _ram_T_311[287:0] : _GEN_11433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12484 = 10'h196 == _T_29 ? _ram_T_311[287:0] : _GEN_11434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12485 = 10'h197 == _T_29 ? _ram_T_311[287:0] : _GEN_11435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12486 = 10'h198 == _T_29 ? _ram_T_311[287:0] : _GEN_11436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12487 = 10'h199 == _T_29 ? _ram_T_311[287:0] : _GEN_11437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12488 = 10'h19a == _T_29 ? _ram_T_311[287:0] : _GEN_11438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12489 = 10'h19b == _T_29 ? _ram_T_311[287:0] : _GEN_11439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12490 = 10'h19c == _T_29 ? _ram_T_311[287:0] : _GEN_11440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12491 = 10'h19d == _T_29 ? _ram_T_311[287:0] : _GEN_11441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12492 = 10'h19e == _T_29 ? _ram_T_311[287:0] : _GEN_11442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12493 = 10'h19f == _T_29 ? _ram_T_311[287:0] : _GEN_11443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12494 = 10'h1a0 == _T_29 ? _ram_T_311[287:0] : _GEN_11444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12495 = 10'h1a1 == _T_29 ? _ram_T_311[287:0] : _GEN_11445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12496 = 10'h1a2 == _T_29 ? _ram_T_311[287:0] : _GEN_11446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12497 = 10'h1a3 == _T_29 ? _ram_T_311[287:0] : _GEN_11447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12498 = 10'h1a4 == _T_29 ? _ram_T_311[287:0] : _GEN_11448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12499 = 10'h1a5 == _T_29 ? _ram_T_311[287:0] : _GEN_11449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12500 = 10'h1a6 == _T_29 ? _ram_T_311[287:0] : _GEN_11450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12501 = 10'h1a7 == _T_29 ? _ram_T_311[287:0] : _GEN_11451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12502 = 10'h1a8 == _T_29 ? _ram_T_311[287:0] : _GEN_11452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12503 = 10'h1a9 == _T_29 ? _ram_T_311[287:0] : _GEN_11453; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12504 = 10'h1aa == _T_29 ? _ram_T_311[287:0] : _GEN_11454; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12505 = 10'h1ab == _T_29 ? _ram_T_311[287:0] : _GEN_11455; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12506 = 10'h1ac == _T_29 ? _ram_T_311[287:0] : _GEN_11456; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12507 = 10'h1ad == _T_29 ? _ram_T_311[287:0] : _GEN_11457; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12508 = 10'h1ae == _T_29 ? _ram_T_311[287:0] : _GEN_11458; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12509 = 10'h1af == _T_29 ? _ram_T_311[287:0] : _GEN_11459; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12510 = 10'h1b0 == _T_29 ? _ram_T_311[287:0] : _GEN_11460; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12511 = 10'h1b1 == _T_29 ? _ram_T_311[287:0] : _GEN_11461; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12512 = 10'h1b2 == _T_29 ? _ram_T_311[287:0] : _GEN_11462; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12513 = 10'h1b3 == _T_29 ? _ram_T_311[287:0] : _GEN_11463; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12514 = 10'h1b4 == _T_29 ? _ram_T_311[287:0] : _GEN_11464; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12515 = 10'h1b5 == _T_29 ? _ram_T_311[287:0] : _GEN_11465; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12516 = 10'h1b6 == _T_29 ? _ram_T_311[287:0] : _GEN_11466; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12517 = 10'h1b7 == _T_29 ? _ram_T_311[287:0] : _GEN_11467; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12518 = 10'h1b8 == _T_29 ? _ram_T_311[287:0] : _GEN_11468; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12519 = 10'h1b9 == _T_29 ? _ram_T_311[287:0] : _GEN_11469; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12520 = 10'h1ba == _T_29 ? _ram_T_311[287:0] : _GEN_11470; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12521 = 10'h1bb == _T_29 ? _ram_T_311[287:0] : _GEN_11471; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12522 = 10'h1bc == _T_29 ? _ram_T_311[287:0] : _GEN_11472; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12523 = 10'h1bd == _T_29 ? _ram_T_311[287:0] : _GEN_11473; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12524 = 10'h1be == _T_29 ? _ram_T_311[287:0] : _GEN_11474; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12525 = 10'h1bf == _T_29 ? _ram_T_311[287:0] : _GEN_11475; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12526 = 10'h1c0 == _T_29 ? _ram_T_311[287:0] : _GEN_11476; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12527 = 10'h1c1 == _T_29 ? _ram_T_311[287:0] : _GEN_11477; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12528 = 10'h1c2 == _T_29 ? _ram_T_311[287:0] : _GEN_11478; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12529 = 10'h1c3 == _T_29 ? _ram_T_311[287:0] : _GEN_11479; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12530 = 10'h1c4 == _T_29 ? _ram_T_311[287:0] : _GEN_11480; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12531 = 10'h1c5 == _T_29 ? _ram_T_311[287:0] : _GEN_11481; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12532 = 10'h1c6 == _T_29 ? _ram_T_311[287:0] : _GEN_11482; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12533 = 10'h1c7 == _T_29 ? _ram_T_311[287:0] : _GEN_11483; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12534 = 10'h1c8 == _T_29 ? _ram_T_311[287:0] : _GEN_11484; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12535 = 10'h1c9 == _T_29 ? _ram_T_311[287:0] : _GEN_11485; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12536 = 10'h1ca == _T_29 ? _ram_T_311[287:0] : _GEN_11486; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12537 = 10'h1cb == _T_29 ? _ram_T_311[287:0] : _GEN_11487; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12538 = 10'h1cc == _T_29 ? _ram_T_311[287:0] : _GEN_11488; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12539 = 10'h1cd == _T_29 ? _ram_T_311[287:0] : _GEN_11489; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12540 = 10'h1ce == _T_29 ? _ram_T_311[287:0] : _GEN_11490; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12541 = 10'h1cf == _T_29 ? _ram_T_311[287:0] : _GEN_11491; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12542 = 10'h1d0 == _T_29 ? _ram_T_311[287:0] : _GEN_11492; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12543 = 10'h1d1 == _T_29 ? _ram_T_311[287:0] : _GEN_11493; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12544 = 10'h1d2 == _T_29 ? _ram_T_311[287:0] : _GEN_11494; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12545 = 10'h1d3 == _T_29 ? _ram_T_311[287:0] : _GEN_11495; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12546 = 10'h1d4 == _T_29 ? _ram_T_311[287:0] : _GEN_11496; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12547 = 10'h1d5 == _T_29 ? _ram_T_311[287:0] : _GEN_11497; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12548 = 10'h1d6 == _T_29 ? _ram_T_311[287:0] : _GEN_11498; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12549 = 10'h1d7 == _T_29 ? _ram_T_311[287:0] : _GEN_11499; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12550 = 10'h1d8 == _T_29 ? _ram_T_311[287:0] : _GEN_11500; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12551 = 10'h1d9 == _T_29 ? _ram_T_311[287:0] : _GEN_11501; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12552 = 10'h1da == _T_29 ? _ram_T_311[287:0] : _GEN_11502; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12553 = 10'h1db == _T_29 ? _ram_T_311[287:0] : _GEN_11503; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12554 = 10'h1dc == _T_29 ? _ram_T_311[287:0] : _GEN_11504; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12555 = 10'h1dd == _T_29 ? _ram_T_311[287:0] : _GEN_11505; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12556 = 10'h1de == _T_29 ? _ram_T_311[287:0] : _GEN_11506; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12557 = 10'h1df == _T_29 ? _ram_T_311[287:0] : _GEN_11507; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12558 = 10'h1e0 == _T_29 ? _ram_T_311[287:0] : _GEN_11508; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12559 = 10'h1e1 == _T_29 ? _ram_T_311[287:0] : _GEN_11509; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12560 = 10'h1e2 == _T_29 ? _ram_T_311[287:0] : _GEN_11510; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12561 = 10'h1e3 == _T_29 ? _ram_T_311[287:0] : _GEN_11511; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12562 = 10'h1e4 == _T_29 ? _ram_T_311[287:0] : _GEN_11512; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12563 = 10'h1e5 == _T_29 ? _ram_T_311[287:0] : _GEN_11513; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12564 = 10'h1e6 == _T_29 ? _ram_T_311[287:0] : _GEN_11514; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12565 = 10'h1e7 == _T_29 ? _ram_T_311[287:0] : _GEN_11515; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12566 = 10'h1e8 == _T_29 ? _ram_T_311[287:0] : _GEN_11516; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12567 = 10'h1e9 == _T_29 ? _ram_T_311[287:0] : _GEN_11517; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12568 = 10'h1ea == _T_29 ? _ram_T_311[287:0] : _GEN_11518; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12569 = 10'h1eb == _T_29 ? _ram_T_311[287:0] : _GEN_11519; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12570 = 10'h1ec == _T_29 ? _ram_T_311[287:0] : _GEN_11520; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12571 = 10'h1ed == _T_29 ? _ram_T_311[287:0] : _GEN_11521; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12572 = 10'h1ee == _T_29 ? _ram_T_311[287:0] : _GEN_11522; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12573 = 10'h1ef == _T_29 ? _ram_T_311[287:0] : _GEN_11523; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12574 = 10'h1f0 == _T_29 ? _ram_T_311[287:0] : _GEN_11524; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12575 = 10'h1f1 == _T_29 ? _ram_T_311[287:0] : _GEN_11525; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12576 = 10'h1f2 == _T_29 ? _ram_T_311[287:0] : _GEN_11526; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12577 = 10'h1f3 == _T_29 ? _ram_T_311[287:0] : _GEN_11527; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12578 = 10'h1f4 == _T_29 ? _ram_T_311[287:0] : _GEN_11528; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12579 = 10'h1f5 == _T_29 ? _ram_T_311[287:0] : _GEN_11529; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12580 = 10'h1f6 == _T_29 ? _ram_T_311[287:0] : _GEN_11530; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12581 = 10'h1f7 == _T_29 ? _ram_T_311[287:0] : _GEN_11531; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12582 = 10'h1f8 == _T_29 ? _ram_T_311[287:0] : _GEN_11532; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12583 = 10'h1f9 == _T_29 ? _ram_T_311[287:0] : _GEN_11533; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12584 = 10'h1fa == _T_29 ? _ram_T_311[287:0] : _GEN_11534; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12585 = 10'h1fb == _T_29 ? _ram_T_311[287:0] : _GEN_11535; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12586 = 10'h1fc == _T_29 ? _ram_T_311[287:0] : _GEN_11536; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12587 = 10'h1fd == _T_29 ? _ram_T_311[287:0] : _GEN_11537; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12588 = 10'h1fe == _T_29 ? _ram_T_311[287:0] : _GEN_11538; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12589 = 10'h1ff == _T_29 ? _ram_T_311[287:0] : _GEN_11539; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12590 = 10'h200 == _T_29 ? _ram_T_311[287:0] : _GEN_11540; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12591 = 10'h201 == _T_29 ? _ram_T_311[287:0] : _GEN_11541; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12592 = 10'h202 == _T_29 ? _ram_T_311[287:0] : _GEN_11542; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12593 = 10'h203 == _T_29 ? _ram_T_311[287:0] : _GEN_11543; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12594 = 10'h204 == _T_29 ? _ram_T_311[287:0] : _GEN_11544; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12595 = 10'h205 == _T_29 ? _ram_T_311[287:0] : _GEN_11545; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12596 = 10'h206 == _T_29 ? _ram_T_311[287:0] : _GEN_11546; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12597 = 10'h207 == _T_29 ? _ram_T_311[287:0] : _GEN_11547; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12598 = 10'h208 == _T_29 ? _ram_T_311[287:0] : _GEN_11548; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12599 = 10'h209 == _T_29 ? _ram_T_311[287:0] : _GEN_11549; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12600 = 10'h20a == _T_29 ? _ram_T_311[287:0] : _GEN_11550; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12601 = 10'h20b == _T_29 ? _ram_T_311[287:0] : _GEN_11551; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_12602 = 10'h20c == _T_29 ? _ram_T_311[287:0] : _GEN_11552; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_31 = h + 10'hc; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_12 = vga_mem_ram_MPORT_108_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_12 = vga_mem_ram_MPORT_109_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_12 = vga_mem_ram_MPORT_110_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_12 = vga_mem_ram_MPORT_111_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_12 = vga_mem_ram_MPORT_112_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_12 = vga_mem_ram_MPORT_113_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_12 = vga_mem_ram_MPORT_114_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_12 = vga_mem_ram_MPORT_115_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_12 = vga_mem_ram_MPORT_116_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_332 = {278'h0,ram_hi_hi_hi_lo_12,ram_hi_hi_lo_12,ram_hi_lo_hi_12,ram_hi_lo_lo_12,
    ram_lo_hi_hi_hi_12,ram_lo_hi_hi_lo_12,ram_lo_hi_lo_12,ram_lo_lo_hi_12,ram_lo_lo_lo_12}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19084 = {{8191'd0}, _ram_T_332}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_336 = _GEN_19084 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_12604 = 10'h1 == _T_31 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12605 = 10'h2 == _T_31 ? ram_2 : _GEN_12604; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12606 = 10'h3 == _T_31 ? ram_3 : _GEN_12605; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12607 = 10'h4 == _T_31 ? ram_4 : _GEN_12606; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12608 = 10'h5 == _T_31 ? ram_5 : _GEN_12607; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12609 = 10'h6 == _T_31 ? ram_6 : _GEN_12608; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12610 = 10'h7 == _T_31 ? ram_7 : _GEN_12609; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12611 = 10'h8 == _T_31 ? ram_8 : _GEN_12610; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12612 = 10'h9 == _T_31 ? ram_9 : _GEN_12611; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12613 = 10'ha == _T_31 ? ram_10 : _GEN_12612; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12614 = 10'hb == _T_31 ? ram_11 : _GEN_12613; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12615 = 10'hc == _T_31 ? ram_12 : _GEN_12614; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12616 = 10'hd == _T_31 ? ram_13 : _GEN_12615; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12617 = 10'he == _T_31 ? ram_14 : _GEN_12616; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12618 = 10'hf == _T_31 ? ram_15 : _GEN_12617; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12619 = 10'h10 == _T_31 ? ram_16 : _GEN_12618; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12620 = 10'h11 == _T_31 ? ram_17 : _GEN_12619; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12621 = 10'h12 == _T_31 ? ram_18 : _GEN_12620; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12622 = 10'h13 == _T_31 ? ram_19 : _GEN_12621; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12623 = 10'h14 == _T_31 ? ram_20 : _GEN_12622; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12624 = 10'h15 == _T_31 ? ram_21 : _GEN_12623; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12625 = 10'h16 == _T_31 ? ram_22 : _GEN_12624; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12626 = 10'h17 == _T_31 ? ram_23 : _GEN_12625; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12627 = 10'h18 == _T_31 ? ram_24 : _GEN_12626; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12628 = 10'h19 == _T_31 ? ram_25 : _GEN_12627; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12629 = 10'h1a == _T_31 ? ram_26 : _GEN_12628; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12630 = 10'h1b == _T_31 ? ram_27 : _GEN_12629; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12631 = 10'h1c == _T_31 ? ram_28 : _GEN_12630; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12632 = 10'h1d == _T_31 ? ram_29 : _GEN_12631; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12633 = 10'h1e == _T_31 ? ram_30 : _GEN_12632; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12634 = 10'h1f == _T_31 ? ram_31 : _GEN_12633; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12635 = 10'h20 == _T_31 ? ram_32 : _GEN_12634; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12636 = 10'h21 == _T_31 ? ram_33 : _GEN_12635; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12637 = 10'h22 == _T_31 ? ram_34 : _GEN_12636; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12638 = 10'h23 == _T_31 ? ram_35 : _GEN_12637; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12639 = 10'h24 == _T_31 ? ram_36 : _GEN_12638; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12640 = 10'h25 == _T_31 ? ram_37 : _GEN_12639; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12641 = 10'h26 == _T_31 ? ram_38 : _GEN_12640; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12642 = 10'h27 == _T_31 ? ram_39 : _GEN_12641; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12643 = 10'h28 == _T_31 ? ram_40 : _GEN_12642; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12644 = 10'h29 == _T_31 ? ram_41 : _GEN_12643; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12645 = 10'h2a == _T_31 ? ram_42 : _GEN_12644; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12646 = 10'h2b == _T_31 ? ram_43 : _GEN_12645; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12647 = 10'h2c == _T_31 ? ram_44 : _GEN_12646; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12648 = 10'h2d == _T_31 ? ram_45 : _GEN_12647; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12649 = 10'h2e == _T_31 ? ram_46 : _GEN_12648; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12650 = 10'h2f == _T_31 ? ram_47 : _GEN_12649; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12651 = 10'h30 == _T_31 ? ram_48 : _GEN_12650; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12652 = 10'h31 == _T_31 ? ram_49 : _GEN_12651; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12653 = 10'h32 == _T_31 ? ram_50 : _GEN_12652; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12654 = 10'h33 == _T_31 ? ram_51 : _GEN_12653; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12655 = 10'h34 == _T_31 ? ram_52 : _GEN_12654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12656 = 10'h35 == _T_31 ? ram_53 : _GEN_12655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12657 = 10'h36 == _T_31 ? ram_54 : _GEN_12656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12658 = 10'h37 == _T_31 ? ram_55 : _GEN_12657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12659 = 10'h38 == _T_31 ? ram_56 : _GEN_12658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12660 = 10'h39 == _T_31 ? ram_57 : _GEN_12659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12661 = 10'h3a == _T_31 ? ram_58 : _GEN_12660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12662 = 10'h3b == _T_31 ? ram_59 : _GEN_12661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12663 = 10'h3c == _T_31 ? ram_60 : _GEN_12662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12664 = 10'h3d == _T_31 ? ram_61 : _GEN_12663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12665 = 10'h3e == _T_31 ? ram_62 : _GEN_12664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12666 = 10'h3f == _T_31 ? ram_63 : _GEN_12665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12667 = 10'h40 == _T_31 ? ram_64 : _GEN_12666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12668 = 10'h41 == _T_31 ? ram_65 : _GEN_12667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12669 = 10'h42 == _T_31 ? ram_66 : _GEN_12668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12670 = 10'h43 == _T_31 ? ram_67 : _GEN_12669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12671 = 10'h44 == _T_31 ? ram_68 : _GEN_12670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12672 = 10'h45 == _T_31 ? ram_69 : _GEN_12671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12673 = 10'h46 == _T_31 ? ram_70 : _GEN_12672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12674 = 10'h47 == _T_31 ? ram_71 : _GEN_12673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12675 = 10'h48 == _T_31 ? ram_72 : _GEN_12674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12676 = 10'h49 == _T_31 ? ram_73 : _GEN_12675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12677 = 10'h4a == _T_31 ? ram_74 : _GEN_12676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12678 = 10'h4b == _T_31 ? ram_75 : _GEN_12677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12679 = 10'h4c == _T_31 ? ram_76 : _GEN_12678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12680 = 10'h4d == _T_31 ? ram_77 : _GEN_12679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12681 = 10'h4e == _T_31 ? ram_78 : _GEN_12680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12682 = 10'h4f == _T_31 ? ram_79 : _GEN_12681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12683 = 10'h50 == _T_31 ? ram_80 : _GEN_12682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12684 = 10'h51 == _T_31 ? ram_81 : _GEN_12683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12685 = 10'h52 == _T_31 ? ram_82 : _GEN_12684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12686 = 10'h53 == _T_31 ? ram_83 : _GEN_12685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12687 = 10'h54 == _T_31 ? ram_84 : _GEN_12686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12688 = 10'h55 == _T_31 ? ram_85 : _GEN_12687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12689 = 10'h56 == _T_31 ? ram_86 : _GEN_12688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12690 = 10'h57 == _T_31 ? ram_87 : _GEN_12689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12691 = 10'h58 == _T_31 ? ram_88 : _GEN_12690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12692 = 10'h59 == _T_31 ? ram_89 : _GEN_12691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12693 = 10'h5a == _T_31 ? ram_90 : _GEN_12692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12694 = 10'h5b == _T_31 ? ram_91 : _GEN_12693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12695 = 10'h5c == _T_31 ? ram_92 : _GEN_12694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12696 = 10'h5d == _T_31 ? ram_93 : _GEN_12695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12697 = 10'h5e == _T_31 ? ram_94 : _GEN_12696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12698 = 10'h5f == _T_31 ? ram_95 : _GEN_12697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12699 = 10'h60 == _T_31 ? ram_96 : _GEN_12698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12700 = 10'h61 == _T_31 ? ram_97 : _GEN_12699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12701 = 10'h62 == _T_31 ? ram_98 : _GEN_12700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12702 = 10'h63 == _T_31 ? ram_99 : _GEN_12701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12703 = 10'h64 == _T_31 ? ram_100 : _GEN_12702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12704 = 10'h65 == _T_31 ? ram_101 : _GEN_12703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12705 = 10'h66 == _T_31 ? ram_102 : _GEN_12704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12706 = 10'h67 == _T_31 ? ram_103 : _GEN_12705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12707 = 10'h68 == _T_31 ? ram_104 : _GEN_12706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12708 = 10'h69 == _T_31 ? ram_105 : _GEN_12707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12709 = 10'h6a == _T_31 ? ram_106 : _GEN_12708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12710 = 10'h6b == _T_31 ? ram_107 : _GEN_12709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12711 = 10'h6c == _T_31 ? ram_108 : _GEN_12710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12712 = 10'h6d == _T_31 ? ram_109 : _GEN_12711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12713 = 10'h6e == _T_31 ? ram_110 : _GEN_12712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12714 = 10'h6f == _T_31 ? ram_111 : _GEN_12713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12715 = 10'h70 == _T_31 ? ram_112 : _GEN_12714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12716 = 10'h71 == _T_31 ? ram_113 : _GEN_12715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12717 = 10'h72 == _T_31 ? ram_114 : _GEN_12716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12718 = 10'h73 == _T_31 ? ram_115 : _GEN_12717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12719 = 10'h74 == _T_31 ? ram_116 : _GEN_12718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12720 = 10'h75 == _T_31 ? ram_117 : _GEN_12719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12721 = 10'h76 == _T_31 ? ram_118 : _GEN_12720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12722 = 10'h77 == _T_31 ? ram_119 : _GEN_12721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12723 = 10'h78 == _T_31 ? ram_120 : _GEN_12722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12724 = 10'h79 == _T_31 ? ram_121 : _GEN_12723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12725 = 10'h7a == _T_31 ? ram_122 : _GEN_12724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12726 = 10'h7b == _T_31 ? ram_123 : _GEN_12725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12727 = 10'h7c == _T_31 ? ram_124 : _GEN_12726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12728 = 10'h7d == _T_31 ? ram_125 : _GEN_12727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12729 = 10'h7e == _T_31 ? ram_126 : _GEN_12728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12730 = 10'h7f == _T_31 ? ram_127 : _GEN_12729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12731 = 10'h80 == _T_31 ? ram_128 : _GEN_12730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12732 = 10'h81 == _T_31 ? ram_129 : _GEN_12731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12733 = 10'h82 == _T_31 ? ram_130 : _GEN_12732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12734 = 10'h83 == _T_31 ? ram_131 : _GEN_12733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12735 = 10'h84 == _T_31 ? ram_132 : _GEN_12734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12736 = 10'h85 == _T_31 ? ram_133 : _GEN_12735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12737 = 10'h86 == _T_31 ? ram_134 : _GEN_12736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12738 = 10'h87 == _T_31 ? ram_135 : _GEN_12737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12739 = 10'h88 == _T_31 ? ram_136 : _GEN_12738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12740 = 10'h89 == _T_31 ? ram_137 : _GEN_12739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12741 = 10'h8a == _T_31 ? ram_138 : _GEN_12740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12742 = 10'h8b == _T_31 ? ram_139 : _GEN_12741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12743 = 10'h8c == _T_31 ? ram_140 : _GEN_12742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12744 = 10'h8d == _T_31 ? ram_141 : _GEN_12743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12745 = 10'h8e == _T_31 ? ram_142 : _GEN_12744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12746 = 10'h8f == _T_31 ? ram_143 : _GEN_12745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12747 = 10'h90 == _T_31 ? ram_144 : _GEN_12746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12748 = 10'h91 == _T_31 ? ram_145 : _GEN_12747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12749 = 10'h92 == _T_31 ? ram_146 : _GEN_12748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12750 = 10'h93 == _T_31 ? ram_147 : _GEN_12749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12751 = 10'h94 == _T_31 ? ram_148 : _GEN_12750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12752 = 10'h95 == _T_31 ? ram_149 : _GEN_12751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12753 = 10'h96 == _T_31 ? ram_150 : _GEN_12752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12754 = 10'h97 == _T_31 ? ram_151 : _GEN_12753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12755 = 10'h98 == _T_31 ? ram_152 : _GEN_12754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12756 = 10'h99 == _T_31 ? ram_153 : _GEN_12755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12757 = 10'h9a == _T_31 ? ram_154 : _GEN_12756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12758 = 10'h9b == _T_31 ? ram_155 : _GEN_12757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12759 = 10'h9c == _T_31 ? ram_156 : _GEN_12758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12760 = 10'h9d == _T_31 ? ram_157 : _GEN_12759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12761 = 10'h9e == _T_31 ? ram_158 : _GEN_12760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12762 = 10'h9f == _T_31 ? ram_159 : _GEN_12761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12763 = 10'ha0 == _T_31 ? ram_160 : _GEN_12762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12764 = 10'ha1 == _T_31 ? ram_161 : _GEN_12763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12765 = 10'ha2 == _T_31 ? ram_162 : _GEN_12764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12766 = 10'ha3 == _T_31 ? ram_163 : _GEN_12765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12767 = 10'ha4 == _T_31 ? ram_164 : _GEN_12766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12768 = 10'ha5 == _T_31 ? ram_165 : _GEN_12767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12769 = 10'ha6 == _T_31 ? ram_166 : _GEN_12768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12770 = 10'ha7 == _T_31 ? ram_167 : _GEN_12769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12771 = 10'ha8 == _T_31 ? ram_168 : _GEN_12770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12772 = 10'ha9 == _T_31 ? ram_169 : _GEN_12771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12773 = 10'haa == _T_31 ? ram_170 : _GEN_12772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12774 = 10'hab == _T_31 ? ram_171 : _GEN_12773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12775 = 10'hac == _T_31 ? ram_172 : _GEN_12774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12776 = 10'had == _T_31 ? ram_173 : _GEN_12775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12777 = 10'hae == _T_31 ? ram_174 : _GEN_12776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12778 = 10'haf == _T_31 ? ram_175 : _GEN_12777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12779 = 10'hb0 == _T_31 ? ram_176 : _GEN_12778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12780 = 10'hb1 == _T_31 ? ram_177 : _GEN_12779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12781 = 10'hb2 == _T_31 ? ram_178 : _GEN_12780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12782 = 10'hb3 == _T_31 ? ram_179 : _GEN_12781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12783 = 10'hb4 == _T_31 ? ram_180 : _GEN_12782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12784 = 10'hb5 == _T_31 ? ram_181 : _GEN_12783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12785 = 10'hb6 == _T_31 ? ram_182 : _GEN_12784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12786 = 10'hb7 == _T_31 ? ram_183 : _GEN_12785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12787 = 10'hb8 == _T_31 ? ram_184 : _GEN_12786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12788 = 10'hb9 == _T_31 ? ram_185 : _GEN_12787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12789 = 10'hba == _T_31 ? ram_186 : _GEN_12788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12790 = 10'hbb == _T_31 ? ram_187 : _GEN_12789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12791 = 10'hbc == _T_31 ? ram_188 : _GEN_12790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12792 = 10'hbd == _T_31 ? ram_189 : _GEN_12791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12793 = 10'hbe == _T_31 ? ram_190 : _GEN_12792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12794 = 10'hbf == _T_31 ? ram_191 : _GEN_12793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12795 = 10'hc0 == _T_31 ? ram_192 : _GEN_12794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12796 = 10'hc1 == _T_31 ? ram_193 : _GEN_12795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12797 = 10'hc2 == _T_31 ? ram_194 : _GEN_12796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12798 = 10'hc3 == _T_31 ? ram_195 : _GEN_12797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12799 = 10'hc4 == _T_31 ? ram_196 : _GEN_12798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12800 = 10'hc5 == _T_31 ? ram_197 : _GEN_12799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12801 = 10'hc6 == _T_31 ? ram_198 : _GEN_12800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12802 = 10'hc7 == _T_31 ? ram_199 : _GEN_12801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12803 = 10'hc8 == _T_31 ? ram_200 : _GEN_12802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12804 = 10'hc9 == _T_31 ? ram_201 : _GEN_12803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12805 = 10'hca == _T_31 ? ram_202 : _GEN_12804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12806 = 10'hcb == _T_31 ? ram_203 : _GEN_12805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12807 = 10'hcc == _T_31 ? ram_204 : _GEN_12806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12808 = 10'hcd == _T_31 ? ram_205 : _GEN_12807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12809 = 10'hce == _T_31 ? ram_206 : _GEN_12808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12810 = 10'hcf == _T_31 ? ram_207 : _GEN_12809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12811 = 10'hd0 == _T_31 ? ram_208 : _GEN_12810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12812 = 10'hd1 == _T_31 ? ram_209 : _GEN_12811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12813 = 10'hd2 == _T_31 ? ram_210 : _GEN_12812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12814 = 10'hd3 == _T_31 ? ram_211 : _GEN_12813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12815 = 10'hd4 == _T_31 ? ram_212 : _GEN_12814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12816 = 10'hd5 == _T_31 ? ram_213 : _GEN_12815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12817 = 10'hd6 == _T_31 ? ram_214 : _GEN_12816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12818 = 10'hd7 == _T_31 ? ram_215 : _GEN_12817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12819 = 10'hd8 == _T_31 ? ram_216 : _GEN_12818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12820 = 10'hd9 == _T_31 ? ram_217 : _GEN_12819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12821 = 10'hda == _T_31 ? ram_218 : _GEN_12820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12822 = 10'hdb == _T_31 ? ram_219 : _GEN_12821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12823 = 10'hdc == _T_31 ? ram_220 : _GEN_12822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12824 = 10'hdd == _T_31 ? ram_221 : _GEN_12823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12825 = 10'hde == _T_31 ? ram_222 : _GEN_12824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12826 = 10'hdf == _T_31 ? ram_223 : _GEN_12825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12827 = 10'he0 == _T_31 ? ram_224 : _GEN_12826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12828 = 10'he1 == _T_31 ? ram_225 : _GEN_12827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12829 = 10'he2 == _T_31 ? ram_226 : _GEN_12828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12830 = 10'he3 == _T_31 ? ram_227 : _GEN_12829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12831 = 10'he4 == _T_31 ? ram_228 : _GEN_12830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12832 = 10'he5 == _T_31 ? ram_229 : _GEN_12831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12833 = 10'he6 == _T_31 ? ram_230 : _GEN_12832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12834 = 10'he7 == _T_31 ? ram_231 : _GEN_12833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12835 = 10'he8 == _T_31 ? ram_232 : _GEN_12834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12836 = 10'he9 == _T_31 ? ram_233 : _GEN_12835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12837 = 10'hea == _T_31 ? ram_234 : _GEN_12836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12838 = 10'heb == _T_31 ? ram_235 : _GEN_12837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12839 = 10'hec == _T_31 ? ram_236 : _GEN_12838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12840 = 10'hed == _T_31 ? ram_237 : _GEN_12839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12841 = 10'hee == _T_31 ? ram_238 : _GEN_12840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12842 = 10'hef == _T_31 ? ram_239 : _GEN_12841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12843 = 10'hf0 == _T_31 ? ram_240 : _GEN_12842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12844 = 10'hf1 == _T_31 ? ram_241 : _GEN_12843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12845 = 10'hf2 == _T_31 ? ram_242 : _GEN_12844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12846 = 10'hf3 == _T_31 ? ram_243 : _GEN_12845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12847 = 10'hf4 == _T_31 ? ram_244 : _GEN_12846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12848 = 10'hf5 == _T_31 ? ram_245 : _GEN_12847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12849 = 10'hf6 == _T_31 ? ram_246 : _GEN_12848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12850 = 10'hf7 == _T_31 ? ram_247 : _GEN_12849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12851 = 10'hf8 == _T_31 ? ram_248 : _GEN_12850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12852 = 10'hf9 == _T_31 ? ram_249 : _GEN_12851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12853 = 10'hfa == _T_31 ? ram_250 : _GEN_12852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12854 = 10'hfb == _T_31 ? ram_251 : _GEN_12853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12855 = 10'hfc == _T_31 ? ram_252 : _GEN_12854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12856 = 10'hfd == _T_31 ? ram_253 : _GEN_12855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12857 = 10'hfe == _T_31 ? ram_254 : _GEN_12856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12858 = 10'hff == _T_31 ? ram_255 : _GEN_12857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12859 = 10'h100 == _T_31 ? ram_256 : _GEN_12858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12860 = 10'h101 == _T_31 ? ram_257 : _GEN_12859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12861 = 10'h102 == _T_31 ? ram_258 : _GEN_12860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12862 = 10'h103 == _T_31 ? ram_259 : _GEN_12861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12863 = 10'h104 == _T_31 ? ram_260 : _GEN_12862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12864 = 10'h105 == _T_31 ? ram_261 : _GEN_12863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12865 = 10'h106 == _T_31 ? ram_262 : _GEN_12864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12866 = 10'h107 == _T_31 ? ram_263 : _GEN_12865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12867 = 10'h108 == _T_31 ? ram_264 : _GEN_12866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12868 = 10'h109 == _T_31 ? ram_265 : _GEN_12867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12869 = 10'h10a == _T_31 ? ram_266 : _GEN_12868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12870 = 10'h10b == _T_31 ? ram_267 : _GEN_12869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12871 = 10'h10c == _T_31 ? ram_268 : _GEN_12870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12872 = 10'h10d == _T_31 ? ram_269 : _GEN_12871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12873 = 10'h10e == _T_31 ? ram_270 : _GEN_12872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12874 = 10'h10f == _T_31 ? ram_271 : _GEN_12873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12875 = 10'h110 == _T_31 ? ram_272 : _GEN_12874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12876 = 10'h111 == _T_31 ? ram_273 : _GEN_12875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12877 = 10'h112 == _T_31 ? ram_274 : _GEN_12876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12878 = 10'h113 == _T_31 ? ram_275 : _GEN_12877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12879 = 10'h114 == _T_31 ? ram_276 : _GEN_12878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12880 = 10'h115 == _T_31 ? ram_277 : _GEN_12879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12881 = 10'h116 == _T_31 ? ram_278 : _GEN_12880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12882 = 10'h117 == _T_31 ? ram_279 : _GEN_12881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12883 = 10'h118 == _T_31 ? ram_280 : _GEN_12882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12884 = 10'h119 == _T_31 ? ram_281 : _GEN_12883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12885 = 10'h11a == _T_31 ? ram_282 : _GEN_12884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12886 = 10'h11b == _T_31 ? ram_283 : _GEN_12885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12887 = 10'h11c == _T_31 ? ram_284 : _GEN_12886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12888 = 10'h11d == _T_31 ? ram_285 : _GEN_12887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12889 = 10'h11e == _T_31 ? ram_286 : _GEN_12888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12890 = 10'h11f == _T_31 ? ram_287 : _GEN_12889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12891 = 10'h120 == _T_31 ? ram_288 : _GEN_12890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12892 = 10'h121 == _T_31 ? ram_289 : _GEN_12891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12893 = 10'h122 == _T_31 ? ram_290 : _GEN_12892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12894 = 10'h123 == _T_31 ? ram_291 : _GEN_12893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12895 = 10'h124 == _T_31 ? ram_292 : _GEN_12894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12896 = 10'h125 == _T_31 ? ram_293 : _GEN_12895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12897 = 10'h126 == _T_31 ? ram_294 : _GEN_12896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12898 = 10'h127 == _T_31 ? ram_295 : _GEN_12897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12899 = 10'h128 == _T_31 ? ram_296 : _GEN_12898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12900 = 10'h129 == _T_31 ? ram_297 : _GEN_12899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12901 = 10'h12a == _T_31 ? ram_298 : _GEN_12900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12902 = 10'h12b == _T_31 ? ram_299 : _GEN_12901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12903 = 10'h12c == _T_31 ? ram_300 : _GEN_12902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12904 = 10'h12d == _T_31 ? ram_301 : _GEN_12903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12905 = 10'h12e == _T_31 ? ram_302 : _GEN_12904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12906 = 10'h12f == _T_31 ? ram_303 : _GEN_12905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12907 = 10'h130 == _T_31 ? ram_304 : _GEN_12906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12908 = 10'h131 == _T_31 ? ram_305 : _GEN_12907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12909 = 10'h132 == _T_31 ? ram_306 : _GEN_12908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12910 = 10'h133 == _T_31 ? ram_307 : _GEN_12909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12911 = 10'h134 == _T_31 ? ram_308 : _GEN_12910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12912 = 10'h135 == _T_31 ? ram_309 : _GEN_12911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12913 = 10'h136 == _T_31 ? ram_310 : _GEN_12912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12914 = 10'h137 == _T_31 ? ram_311 : _GEN_12913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12915 = 10'h138 == _T_31 ? ram_312 : _GEN_12914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12916 = 10'h139 == _T_31 ? ram_313 : _GEN_12915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12917 = 10'h13a == _T_31 ? ram_314 : _GEN_12916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12918 = 10'h13b == _T_31 ? ram_315 : _GEN_12917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12919 = 10'h13c == _T_31 ? ram_316 : _GEN_12918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12920 = 10'h13d == _T_31 ? ram_317 : _GEN_12919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12921 = 10'h13e == _T_31 ? ram_318 : _GEN_12920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12922 = 10'h13f == _T_31 ? ram_319 : _GEN_12921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12923 = 10'h140 == _T_31 ? ram_320 : _GEN_12922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12924 = 10'h141 == _T_31 ? ram_321 : _GEN_12923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12925 = 10'h142 == _T_31 ? ram_322 : _GEN_12924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12926 = 10'h143 == _T_31 ? ram_323 : _GEN_12925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12927 = 10'h144 == _T_31 ? ram_324 : _GEN_12926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12928 = 10'h145 == _T_31 ? ram_325 : _GEN_12927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12929 = 10'h146 == _T_31 ? ram_326 : _GEN_12928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12930 = 10'h147 == _T_31 ? ram_327 : _GEN_12929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12931 = 10'h148 == _T_31 ? ram_328 : _GEN_12930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12932 = 10'h149 == _T_31 ? ram_329 : _GEN_12931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12933 = 10'h14a == _T_31 ? ram_330 : _GEN_12932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12934 = 10'h14b == _T_31 ? ram_331 : _GEN_12933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12935 = 10'h14c == _T_31 ? ram_332 : _GEN_12934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12936 = 10'h14d == _T_31 ? ram_333 : _GEN_12935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12937 = 10'h14e == _T_31 ? ram_334 : _GEN_12936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12938 = 10'h14f == _T_31 ? ram_335 : _GEN_12937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12939 = 10'h150 == _T_31 ? ram_336 : _GEN_12938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12940 = 10'h151 == _T_31 ? ram_337 : _GEN_12939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12941 = 10'h152 == _T_31 ? ram_338 : _GEN_12940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12942 = 10'h153 == _T_31 ? ram_339 : _GEN_12941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12943 = 10'h154 == _T_31 ? ram_340 : _GEN_12942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12944 = 10'h155 == _T_31 ? ram_341 : _GEN_12943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12945 = 10'h156 == _T_31 ? ram_342 : _GEN_12944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12946 = 10'h157 == _T_31 ? ram_343 : _GEN_12945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12947 = 10'h158 == _T_31 ? ram_344 : _GEN_12946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12948 = 10'h159 == _T_31 ? ram_345 : _GEN_12947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12949 = 10'h15a == _T_31 ? ram_346 : _GEN_12948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12950 = 10'h15b == _T_31 ? ram_347 : _GEN_12949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12951 = 10'h15c == _T_31 ? ram_348 : _GEN_12950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12952 = 10'h15d == _T_31 ? ram_349 : _GEN_12951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12953 = 10'h15e == _T_31 ? ram_350 : _GEN_12952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12954 = 10'h15f == _T_31 ? ram_351 : _GEN_12953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12955 = 10'h160 == _T_31 ? ram_352 : _GEN_12954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12956 = 10'h161 == _T_31 ? ram_353 : _GEN_12955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12957 = 10'h162 == _T_31 ? ram_354 : _GEN_12956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12958 = 10'h163 == _T_31 ? ram_355 : _GEN_12957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12959 = 10'h164 == _T_31 ? ram_356 : _GEN_12958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12960 = 10'h165 == _T_31 ? ram_357 : _GEN_12959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12961 = 10'h166 == _T_31 ? ram_358 : _GEN_12960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12962 = 10'h167 == _T_31 ? ram_359 : _GEN_12961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12963 = 10'h168 == _T_31 ? ram_360 : _GEN_12962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12964 = 10'h169 == _T_31 ? ram_361 : _GEN_12963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12965 = 10'h16a == _T_31 ? ram_362 : _GEN_12964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12966 = 10'h16b == _T_31 ? ram_363 : _GEN_12965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12967 = 10'h16c == _T_31 ? ram_364 : _GEN_12966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12968 = 10'h16d == _T_31 ? ram_365 : _GEN_12967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12969 = 10'h16e == _T_31 ? ram_366 : _GEN_12968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12970 = 10'h16f == _T_31 ? ram_367 : _GEN_12969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12971 = 10'h170 == _T_31 ? ram_368 : _GEN_12970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12972 = 10'h171 == _T_31 ? ram_369 : _GEN_12971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12973 = 10'h172 == _T_31 ? ram_370 : _GEN_12972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12974 = 10'h173 == _T_31 ? ram_371 : _GEN_12973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12975 = 10'h174 == _T_31 ? ram_372 : _GEN_12974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12976 = 10'h175 == _T_31 ? ram_373 : _GEN_12975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12977 = 10'h176 == _T_31 ? ram_374 : _GEN_12976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12978 = 10'h177 == _T_31 ? ram_375 : _GEN_12977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12979 = 10'h178 == _T_31 ? ram_376 : _GEN_12978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12980 = 10'h179 == _T_31 ? ram_377 : _GEN_12979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12981 = 10'h17a == _T_31 ? ram_378 : _GEN_12980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12982 = 10'h17b == _T_31 ? ram_379 : _GEN_12981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12983 = 10'h17c == _T_31 ? ram_380 : _GEN_12982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12984 = 10'h17d == _T_31 ? ram_381 : _GEN_12983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12985 = 10'h17e == _T_31 ? ram_382 : _GEN_12984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12986 = 10'h17f == _T_31 ? ram_383 : _GEN_12985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12987 = 10'h180 == _T_31 ? ram_384 : _GEN_12986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12988 = 10'h181 == _T_31 ? ram_385 : _GEN_12987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12989 = 10'h182 == _T_31 ? ram_386 : _GEN_12988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12990 = 10'h183 == _T_31 ? ram_387 : _GEN_12989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12991 = 10'h184 == _T_31 ? ram_388 : _GEN_12990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12992 = 10'h185 == _T_31 ? ram_389 : _GEN_12991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12993 = 10'h186 == _T_31 ? ram_390 : _GEN_12992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12994 = 10'h187 == _T_31 ? ram_391 : _GEN_12993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12995 = 10'h188 == _T_31 ? ram_392 : _GEN_12994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12996 = 10'h189 == _T_31 ? ram_393 : _GEN_12995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12997 = 10'h18a == _T_31 ? ram_394 : _GEN_12996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12998 = 10'h18b == _T_31 ? ram_395 : _GEN_12997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_12999 = 10'h18c == _T_31 ? ram_396 : _GEN_12998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13000 = 10'h18d == _T_31 ? ram_397 : _GEN_12999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13001 = 10'h18e == _T_31 ? ram_398 : _GEN_13000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13002 = 10'h18f == _T_31 ? ram_399 : _GEN_13001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13003 = 10'h190 == _T_31 ? ram_400 : _GEN_13002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13004 = 10'h191 == _T_31 ? ram_401 : _GEN_13003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13005 = 10'h192 == _T_31 ? ram_402 : _GEN_13004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13006 = 10'h193 == _T_31 ? ram_403 : _GEN_13005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13007 = 10'h194 == _T_31 ? ram_404 : _GEN_13006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13008 = 10'h195 == _T_31 ? ram_405 : _GEN_13007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13009 = 10'h196 == _T_31 ? ram_406 : _GEN_13008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13010 = 10'h197 == _T_31 ? ram_407 : _GEN_13009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13011 = 10'h198 == _T_31 ? ram_408 : _GEN_13010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13012 = 10'h199 == _T_31 ? ram_409 : _GEN_13011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13013 = 10'h19a == _T_31 ? ram_410 : _GEN_13012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13014 = 10'h19b == _T_31 ? ram_411 : _GEN_13013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13015 = 10'h19c == _T_31 ? ram_412 : _GEN_13014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13016 = 10'h19d == _T_31 ? ram_413 : _GEN_13015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13017 = 10'h19e == _T_31 ? ram_414 : _GEN_13016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13018 = 10'h19f == _T_31 ? ram_415 : _GEN_13017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13019 = 10'h1a0 == _T_31 ? ram_416 : _GEN_13018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13020 = 10'h1a1 == _T_31 ? ram_417 : _GEN_13019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13021 = 10'h1a2 == _T_31 ? ram_418 : _GEN_13020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13022 = 10'h1a3 == _T_31 ? ram_419 : _GEN_13021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13023 = 10'h1a4 == _T_31 ? ram_420 : _GEN_13022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13024 = 10'h1a5 == _T_31 ? ram_421 : _GEN_13023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13025 = 10'h1a6 == _T_31 ? ram_422 : _GEN_13024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13026 = 10'h1a7 == _T_31 ? ram_423 : _GEN_13025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13027 = 10'h1a8 == _T_31 ? ram_424 : _GEN_13026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13028 = 10'h1a9 == _T_31 ? ram_425 : _GEN_13027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13029 = 10'h1aa == _T_31 ? ram_426 : _GEN_13028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13030 = 10'h1ab == _T_31 ? ram_427 : _GEN_13029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13031 = 10'h1ac == _T_31 ? ram_428 : _GEN_13030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13032 = 10'h1ad == _T_31 ? ram_429 : _GEN_13031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13033 = 10'h1ae == _T_31 ? ram_430 : _GEN_13032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13034 = 10'h1af == _T_31 ? ram_431 : _GEN_13033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13035 = 10'h1b0 == _T_31 ? ram_432 : _GEN_13034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13036 = 10'h1b1 == _T_31 ? ram_433 : _GEN_13035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13037 = 10'h1b2 == _T_31 ? ram_434 : _GEN_13036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13038 = 10'h1b3 == _T_31 ? ram_435 : _GEN_13037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13039 = 10'h1b4 == _T_31 ? ram_436 : _GEN_13038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13040 = 10'h1b5 == _T_31 ? ram_437 : _GEN_13039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13041 = 10'h1b6 == _T_31 ? ram_438 : _GEN_13040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13042 = 10'h1b7 == _T_31 ? ram_439 : _GEN_13041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13043 = 10'h1b8 == _T_31 ? ram_440 : _GEN_13042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13044 = 10'h1b9 == _T_31 ? ram_441 : _GEN_13043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13045 = 10'h1ba == _T_31 ? ram_442 : _GEN_13044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13046 = 10'h1bb == _T_31 ? ram_443 : _GEN_13045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13047 = 10'h1bc == _T_31 ? ram_444 : _GEN_13046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13048 = 10'h1bd == _T_31 ? ram_445 : _GEN_13047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13049 = 10'h1be == _T_31 ? ram_446 : _GEN_13048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13050 = 10'h1bf == _T_31 ? ram_447 : _GEN_13049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13051 = 10'h1c0 == _T_31 ? ram_448 : _GEN_13050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13052 = 10'h1c1 == _T_31 ? ram_449 : _GEN_13051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13053 = 10'h1c2 == _T_31 ? ram_450 : _GEN_13052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13054 = 10'h1c3 == _T_31 ? ram_451 : _GEN_13053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13055 = 10'h1c4 == _T_31 ? ram_452 : _GEN_13054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13056 = 10'h1c5 == _T_31 ? ram_453 : _GEN_13055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13057 = 10'h1c6 == _T_31 ? ram_454 : _GEN_13056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13058 = 10'h1c7 == _T_31 ? ram_455 : _GEN_13057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13059 = 10'h1c8 == _T_31 ? ram_456 : _GEN_13058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13060 = 10'h1c9 == _T_31 ? ram_457 : _GEN_13059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13061 = 10'h1ca == _T_31 ? ram_458 : _GEN_13060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13062 = 10'h1cb == _T_31 ? ram_459 : _GEN_13061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13063 = 10'h1cc == _T_31 ? ram_460 : _GEN_13062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13064 = 10'h1cd == _T_31 ? ram_461 : _GEN_13063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13065 = 10'h1ce == _T_31 ? ram_462 : _GEN_13064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13066 = 10'h1cf == _T_31 ? ram_463 : _GEN_13065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13067 = 10'h1d0 == _T_31 ? ram_464 : _GEN_13066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13068 = 10'h1d1 == _T_31 ? ram_465 : _GEN_13067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13069 = 10'h1d2 == _T_31 ? ram_466 : _GEN_13068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13070 = 10'h1d3 == _T_31 ? ram_467 : _GEN_13069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13071 = 10'h1d4 == _T_31 ? ram_468 : _GEN_13070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13072 = 10'h1d5 == _T_31 ? ram_469 : _GEN_13071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13073 = 10'h1d6 == _T_31 ? ram_470 : _GEN_13072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13074 = 10'h1d7 == _T_31 ? ram_471 : _GEN_13073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13075 = 10'h1d8 == _T_31 ? ram_472 : _GEN_13074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13076 = 10'h1d9 == _T_31 ? ram_473 : _GEN_13075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13077 = 10'h1da == _T_31 ? ram_474 : _GEN_13076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13078 = 10'h1db == _T_31 ? ram_475 : _GEN_13077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13079 = 10'h1dc == _T_31 ? ram_476 : _GEN_13078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13080 = 10'h1dd == _T_31 ? ram_477 : _GEN_13079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13081 = 10'h1de == _T_31 ? ram_478 : _GEN_13080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13082 = 10'h1df == _T_31 ? ram_479 : _GEN_13081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13083 = 10'h1e0 == _T_31 ? ram_480 : _GEN_13082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13084 = 10'h1e1 == _T_31 ? ram_481 : _GEN_13083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13085 = 10'h1e2 == _T_31 ? ram_482 : _GEN_13084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13086 = 10'h1e3 == _T_31 ? ram_483 : _GEN_13085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13087 = 10'h1e4 == _T_31 ? ram_484 : _GEN_13086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13088 = 10'h1e5 == _T_31 ? ram_485 : _GEN_13087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13089 = 10'h1e6 == _T_31 ? ram_486 : _GEN_13088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13090 = 10'h1e7 == _T_31 ? ram_487 : _GEN_13089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13091 = 10'h1e8 == _T_31 ? ram_488 : _GEN_13090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13092 = 10'h1e9 == _T_31 ? ram_489 : _GEN_13091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13093 = 10'h1ea == _T_31 ? ram_490 : _GEN_13092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13094 = 10'h1eb == _T_31 ? ram_491 : _GEN_13093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13095 = 10'h1ec == _T_31 ? ram_492 : _GEN_13094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13096 = 10'h1ed == _T_31 ? ram_493 : _GEN_13095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13097 = 10'h1ee == _T_31 ? ram_494 : _GEN_13096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13098 = 10'h1ef == _T_31 ? ram_495 : _GEN_13097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13099 = 10'h1f0 == _T_31 ? ram_496 : _GEN_13098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13100 = 10'h1f1 == _T_31 ? ram_497 : _GEN_13099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13101 = 10'h1f2 == _T_31 ? ram_498 : _GEN_13100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13102 = 10'h1f3 == _T_31 ? ram_499 : _GEN_13101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13103 = 10'h1f4 == _T_31 ? ram_500 : _GEN_13102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13104 = 10'h1f5 == _T_31 ? ram_501 : _GEN_13103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13105 = 10'h1f6 == _T_31 ? ram_502 : _GEN_13104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13106 = 10'h1f7 == _T_31 ? ram_503 : _GEN_13105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13107 = 10'h1f8 == _T_31 ? ram_504 : _GEN_13106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13108 = 10'h1f9 == _T_31 ? ram_505 : _GEN_13107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13109 = 10'h1fa == _T_31 ? ram_506 : _GEN_13108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13110 = 10'h1fb == _T_31 ? ram_507 : _GEN_13109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13111 = 10'h1fc == _T_31 ? ram_508 : _GEN_13110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13112 = 10'h1fd == _T_31 ? ram_509 : _GEN_13111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13113 = 10'h1fe == _T_31 ? ram_510 : _GEN_13112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13114 = 10'h1ff == _T_31 ? ram_511 : _GEN_13113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13115 = 10'h200 == _T_31 ? ram_512 : _GEN_13114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13116 = 10'h201 == _T_31 ? ram_513 : _GEN_13115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13117 = 10'h202 == _T_31 ? ram_514 : _GEN_13116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13118 = 10'h203 == _T_31 ? ram_515 : _GEN_13117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13119 = 10'h204 == _T_31 ? ram_516 : _GEN_13118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13120 = 10'h205 == _T_31 ? ram_517 : _GEN_13119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13121 = 10'h206 == _T_31 ? ram_518 : _GEN_13120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13122 = 10'h207 == _T_31 ? ram_519 : _GEN_13121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13123 = 10'h208 == _T_31 ? ram_520 : _GEN_13122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13124 = 10'h209 == _T_31 ? ram_521 : _GEN_13123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13125 = 10'h20a == _T_31 ? ram_522 : _GEN_13124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13126 = 10'h20b == _T_31 ? ram_523 : _GEN_13125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13127 = 10'h20c == _T_31 ? ram_524 : _GEN_13126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19085 = {{8190'd0}, _GEN_13127}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_337 = _GEN_19085 ^ _ram_T_336; // @[vga.scala 64:41]
  wire [287:0] _GEN_13128 = 10'h0 == _T_31 ? _ram_T_337[287:0] : _GEN_12078; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13129 = 10'h1 == _T_31 ? _ram_T_337[287:0] : _GEN_12079; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13130 = 10'h2 == _T_31 ? _ram_T_337[287:0] : _GEN_12080; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13131 = 10'h3 == _T_31 ? _ram_T_337[287:0] : _GEN_12081; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13132 = 10'h4 == _T_31 ? _ram_T_337[287:0] : _GEN_12082; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13133 = 10'h5 == _T_31 ? _ram_T_337[287:0] : _GEN_12083; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13134 = 10'h6 == _T_31 ? _ram_T_337[287:0] : _GEN_12084; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13135 = 10'h7 == _T_31 ? _ram_T_337[287:0] : _GEN_12085; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13136 = 10'h8 == _T_31 ? _ram_T_337[287:0] : _GEN_12086; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13137 = 10'h9 == _T_31 ? _ram_T_337[287:0] : _GEN_12087; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13138 = 10'ha == _T_31 ? _ram_T_337[287:0] : _GEN_12088; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13139 = 10'hb == _T_31 ? _ram_T_337[287:0] : _GEN_12089; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13140 = 10'hc == _T_31 ? _ram_T_337[287:0] : _GEN_12090; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13141 = 10'hd == _T_31 ? _ram_T_337[287:0] : _GEN_12091; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13142 = 10'he == _T_31 ? _ram_T_337[287:0] : _GEN_12092; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13143 = 10'hf == _T_31 ? _ram_T_337[287:0] : _GEN_12093; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13144 = 10'h10 == _T_31 ? _ram_T_337[287:0] : _GEN_12094; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13145 = 10'h11 == _T_31 ? _ram_T_337[287:0] : _GEN_12095; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13146 = 10'h12 == _T_31 ? _ram_T_337[287:0] : _GEN_12096; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13147 = 10'h13 == _T_31 ? _ram_T_337[287:0] : _GEN_12097; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13148 = 10'h14 == _T_31 ? _ram_T_337[287:0] : _GEN_12098; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13149 = 10'h15 == _T_31 ? _ram_T_337[287:0] : _GEN_12099; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13150 = 10'h16 == _T_31 ? _ram_T_337[287:0] : _GEN_12100; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13151 = 10'h17 == _T_31 ? _ram_T_337[287:0] : _GEN_12101; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13152 = 10'h18 == _T_31 ? _ram_T_337[287:0] : _GEN_12102; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13153 = 10'h19 == _T_31 ? _ram_T_337[287:0] : _GEN_12103; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13154 = 10'h1a == _T_31 ? _ram_T_337[287:0] : _GEN_12104; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13155 = 10'h1b == _T_31 ? _ram_T_337[287:0] : _GEN_12105; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13156 = 10'h1c == _T_31 ? _ram_T_337[287:0] : _GEN_12106; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13157 = 10'h1d == _T_31 ? _ram_T_337[287:0] : _GEN_12107; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13158 = 10'h1e == _T_31 ? _ram_T_337[287:0] : _GEN_12108; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13159 = 10'h1f == _T_31 ? _ram_T_337[287:0] : _GEN_12109; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13160 = 10'h20 == _T_31 ? _ram_T_337[287:0] : _GEN_12110; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13161 = 10'h21 == _T_31 ? _ram_T_337[287:0] : _GEN_12111; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13162 = 10'h22 == _T_31 ? _ram_T_337[287:0] : _GEN_12112; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13163 = 10'h23 == _T_31 ? _ram_T_337[287:0] : _GEN_12113; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13164 = 10'h24 == _T_31 ? _ram_T_337[287:0] : _GEN_12114; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13165 = 10'h25 == _T_31 ? _ram_T_337[287:0] : _GEN_12115; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13166 = 10'h26 == _T_31 ? _ram_T_337[287:0] : _GEN_12116; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13167 = 10'h27 == _T_31 ? _ram_T_337[287:0] : _GEN_12117; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13168 = 10'h28 == _T_31 ? _ram_T_337[287:0] : _GEN_12118; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13169 = 10'h29 == _T_31 ? _ram_T_337[287:0] : _GEN_12119; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13170 = 10'h2a == _T_31 ? _ram_T_337[287:0] : _GEN_12120; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13171 = 10'h2b == _T_31 ? _ram_T_337[287:0] : _GEN_12121; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13172 = 10'h2c == _T_31 ? _ram_T_337[287:0] : _GEN_12122; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13173 = 10'h2d == _T_31 ? _ram_T_337[287:0] : _GEN_12123; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13174 = 10'h2e == _T_31 ? _ram_T_337[287:0] : _GEN_12124; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13175 = 10'h2f == _T_31 ? _ram_T_337[287:0] : _GEN_12125; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13176 = 10'h30 == _T_31 ? _ram_T_337[287:0] : _GEN_12126; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13177 = 10'h31 == _T_31 ? _ram_T_337[287:0] : _GEN_12127; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13178 = 10'h32 == _T_31 ? _ram_T_337[287:0] : _GEN_12128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13179 = 10'h33 == _T_31 ? _ram_T_337[287:0] : _GEN_12129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13180 = 10'h34 == _T_31 ? _ram_T_337[287:0] : _GEN_12130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13181 = 10'h35 == _T_31 ? _ram_T_337[287:0] : _GEN_12131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13182 = 10'h36 == _T_31 ? _ram_T_337[287:0] : _GEN_12132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13183 = 10'h37 == _T_31 ? _ram_T_337[287:0] : _GEN_12133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13184 = 10'h38 == _T_31 ? _ram_T_337[287:0] : _GEN_12134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13185 = 10'h39 == _T_31 ? _ram_T_337[287:0] : _GEN_12135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13186 = 10'h3a == _T_31 ? _ram_T_337[287:0] : _GEN_12136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13187 = 10'h3b == _T_31 ? _ram_T_337[287:0] : _GEN_12137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13188 = 10'h3c == _T_31 ? _ram_T_337[287:0] : _GEN_12138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13189 = 10'h3d == _T_31 ? _ram_T_337[287:0] : _GEN_12139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13190 = 10'h3e == _T_31 ? _ram_T_337[287:0] : _GEN_12140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13191 = 10'h3f == _T_31 ? _ram_T_337[287:0] : _GEN_12141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13192 = 10'h40 == _T_31 ? _ram_T_337[287:0] : _GEN_12142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13193 = 10'h41 == _T_31 ? _ram_T_337[287:0] : _GEN_12143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13194 = 10'h42 == _T_31 ? _ram_T_337[287:0] : _GEN_12144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13195 = 10'h43 == _T_31 ? _ram_T_337[287:0] : _GEN_12145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13196 = 10'h44 == _T_31 ? _ram_T_337[287:0] : _GEN_12146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13197 = 10'h45 == _T_31 ? _ram_T_337[287:0] : _GEN_12147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13198 = 10'h46 == _T_31 ? _ram_T_337[287:0] : _GEN_12148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13199 = 10'h47 == _T_31 ? _ram_T_337[287:0] : _GEN_12149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13200 = 10'h48 == _T_31 ? _ram_T_337[287:0] : _GEN_12150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13201 = 10'h49 == _T_31 ? _ram_T_337[287:0] : _GEN_12151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13202 = 10'h4a == _T_31 ? _ram_T_337[287:0] : _GEN_12152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13203 = 10'h4b == _T_31 ? _ram_T_337[287:0] : _GEN_12153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13204 = 10'h4c == _T_31 ? _ram_T_337[287:0] : _GEN_12154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13205 = 10'h4d == _T_31 ? _ram_T_337[287:0] : _GEN_12155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13206 = 10'h4e == _T_31 ? _ram_T_337[287:0] : _GEN_12156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13207 = 10'h4f == _T_31 ? _ram_T_337[287:0] : _GEN_12157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13208 = 10'h50 == _T_31 ? _ram_T_337[287:0] : _GEN_12158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13209 = 10'h51 == _T_31 ? _ram_T_337[287:0] : _GEN_12159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13210 = 10'h52 == _T_31 ? _ram_T_337[287:0] : _GEN_12160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13211 = 10'h53 == _T_31 ? _ram_T_337[287:0] : _GEN_12161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13212 = 10'h54 == _T_31 ? _ram_T_337[287:0] : _GEN_12162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13213 = 10'h55 == _T_31 ? _ram_T_337[287:0] : _GEN_12163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13214 = 10'h56 == _T_31 ? _ram_T_337[287:0] : _GEN_12164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13215 = 10'h57 == _T_31 ? _ram_T_337[287:0] : _GEN_12165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13216 = 10'h58 == _T_31 ? _ram_T_337[287:0] : _GEN_12166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13217 = 10'h59 == _T_31 ? _ram_T_337[287:0] : _GEN_12167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13218 = 10'h5a == _T_31 ? _ram_T_337[287:0] : _GEN_12168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13219 = 10'h5b == _T_31 ? _ram_T_337[287:0] : _GEN_12169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13220 = 10'h5c == _T_31 ? _ram_T_337[287:0] : _GEN_12170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13221 = 10'h5d == _T_31 ? _ram_T_337[287:0] : _GEN_12171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13222 = 10'h5e == _T_31 ? _ram_T_337[287:0] : _GEN_12172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13223 = 10'h5f == _T_31 ? _ram_T_337[287:0] : _GEN_12173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13224 = 10'h60 == _T_31 ? _ram_T_337[287:0] : _GEN_12174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13225 = 10'h61 == _T_31 ? _ram_T_337[287:0] : _GEN_12175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13226 = 10'h62 == _T_31 ? _ram_T_337[287:0] : _GEN_12176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13227 = 10'h63 == _T_31 ? _ram_T_337[287:0] : _GEN_12177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13228 = 10'h64 == _T_31 ? _ram_T_337[287:0] : _GEN_12178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13229 = 10'h65 == _T_31 ? _ram_T_337[287:0] : _GEN_12179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13230 = 10'h66 == _T_31 ? _ram_T_337[287:0] : _GEN_12180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13231 = 10'h67 == _T_31 ? _ram_T_337[287:0] : _GEN_12181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13232 = 10'h68 == _T_31 ? _ram_T_337[287:0] : _GEN_12182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13233 = 10'h69 == _T_31 ? _ram_T_337[287:0] : _GEN_12183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13234 = 10'h6a == _T_31 ? _ram_T_337[287:0] : _GEN_12184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13235 = 10'h6b == _T_31 ? _ram_T_337[287:0] : _GEN_12185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13236 = 10'h6c == _T_31 ? _ram_T_337[287:0] : _GEN_12186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13237 = 10'h6d == _T_31 ? _ram_T_337[287:0] : _GEN_12187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13238 = 10'h6e == _T_31 ? _ram_T_337[287:0] : _GEN_12188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13239 = 10'h6f == _T_31 ? _ram_T_337[287:0] : _GEN_12189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13240 = 10'h70 == _T_31 ? _ram_T_337[287:0] : _GEN_12190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13241 = 10'h71 == _T_31 ? _ram_T_337[287:0] : _GEN_12191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13242 = 10'h72 == _T_31 ? _ram_T_337[287:0] : _GEN_12192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13243 = 10'h73 == _T_31 ? _ram_T_337[287:0] : _GEN_12193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13244 = 10'h74 == _T_31 ? _ram_T_337[287:0] : _GEN_12194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13245 = 10'h75 == _T_31 ? _ram_T_337[287:0] : _GEN_12195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13246 = 10'h76 == _T_31 ? _ram_T_337[287:0] : _GEN_12196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13247 = 10'h77 == _T_31 ? _ram_T_337[287:0] : _GEN_12197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13248 = 10'h78 == _T_31 ? _ram_T_337[287:0] : _GEN_12198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13249 = 10'h79 == _T_31 ? _ram_T_337[287:0] : _GEN_12199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13250 = 10'h7a == _T_31 ? _ram_T_337[287:0] : _GEN_12200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13251 = 10'h7b == _T_31 ? _ram_T_337[287:0] : _GEN_12201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13252 = 10'h7c == _T_31 ? _ram_T_337[287:0] : _GEN_12202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13253 = 10'h7d == _T_31 ? _ram_T_337[287:0] : _GEN_12203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13254 = 10'h7e == _T_31 ? _ram_T_337[287:0] : _GEN_12204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13255 = 10'h7f == _T_31 ? _ram_T_337[287:0] : _GEN_12205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13256 = 10'h80 == _T_31 ? _ram_T_337[287:0] : _GEN_12206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13257 = 10'h81 == _T_31 ? _ram_T_337[287:0] : _GEN_12207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13258 = 10'h82 == _T_31 ? _ram_T_337[287:0] : _GEN_12208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13259 = 10'h83 == _T_31 ? _ram_T_337[287:0] : _GEN_12209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13260 = 10'h84 == _T_31 ? _ram_T_337[287:0] : _GEN_12210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13261 = 10'h85 == _T_31 ? _ram_T_337[287:0] : _GEN_12211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13262 = 10'h86 == _T_31 ? _ram_T_337[287:0] : _GEN_12212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13263 = 10'h87 == _T_31 ? _ram_T_337[287:0] : _GEN_12213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13264 = 10'h88 == _T_31 ? _ram_T_337[287:0] : _GEN_12214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13265 = 10'h89 == _T_31 ? _ram_T_337[287:0] : _GEN_12215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13266 = 10'h8a == _T_31 ? _ram_T_337[287:0] : _GEN_12216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13267 = 10'h8b == _T_31 ? _ram_T_337[287:0] : _GEN_12217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13268 = 10'h8c == _T_31 ? _ram_T_337[287:0] : _GEN_12218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13269 = 10'h8d == _T_31 ? _ram_T_337[287:0] : _GEN_12219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13270 = 10'h8e == _T_31 ? _ram_T_337[287:0] : _GEN_12220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13271 = 10'h8f == _T_31 ? _ram_T_337[287:0] : _GEN_12221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13272 = 10'h90 == _T_31 ? _ram_T_337[287:0] : _GEN_12222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13273 = 10'h91 == _T_31 ? _ram_T_337[287:0] : _GEN_12223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13274 = 10'h92 == _T_31 ? _ram_T_337[287:0] : _GEN_12224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13275 = 10'h93 == _T_31 ? _ram_T_337[287:0] : _GEN_12225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13276 = 10'h94 == _T_31 ? _ram_T_337[287:0] : _GEN_12226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13277 = 10'h95 == _T_31 ? _ram_T_337[287:0] : _GEN_12227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13278 = 10'h96 == _T_31 ? _ram_T_337[287:0] : _GEN_12228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13279 = 10'h97 == _T_31 ? _ram_T_337[287:0] : _GEN_12229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13280 = 10'h98 == _T_31 ? _ram_T_337[287:0] : _GEN_12230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13281 = 10'h99 == _T_31 ? _ram_T_337[287:0] : _GEN_12231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13282 = 10'h9a == _T_31 ? _ram_T_337[287:0] : _GEN_12232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13283 = 10'h9b == _T_31 ? _ram_T_337[287:0] : _GEN_12233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13284 = 10'h9c == _T_31 ? _ram_T_337[287:0] : _GEN_12234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13285 = 10'h9d == _T_31 ? _ram_T_337[287:0] : _GEN_12235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13286 = 10'h9e == _T_31 ? _ram_T_337[287:0] : _GEN_12236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13287 = 10'h9f == _T_31 ? _ram_T_337[287:0] : _GEN_12237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13288 = 10'ha0 == _T_31 ? _ram_T_337[287:0] : _GEN_12238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13289 = 10'ha1 == _T_31 ? _ram_T_337[287:0] : _GEN_12239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13290 = 10'ha2 == _T_31 ? _ram_T_337[287:0] : _GEN_12240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13291 = 10'ha3 == _T_31 ? _ram_T_337[287:0] : _GEN_12241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13292 = 10'ha4 == _T_31 ? _ram_T_337[287:0] : _GEN_12242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13293 = 10'ha5 == _T_31 ? _ram_T_337[287:0] : _GEN_12243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13294 = 10'ha6 == _T_31 ? _ram_T_337[287:0] : _GEN_12244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13295 = 10'ha7 == _T_31 ? _ram_T_337[287:0] : _GEN_12245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13296 = 10'ha8 == _T_31 ? _ram_T_337[287:0] : _GEN_12246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13297 = 10'ha9 == _T_31 ? _ram_T_337[287:0] : _GEN_12247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13298 = 10'haa == _T_31 ? _ram_T_337[287:0] : _GEN_12248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13299 = 10'hab == _T_31 ? _ram_T_337[287:0] : _GEN_12249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13300 = 10'hac == _T_31 ? _ram_T_337[287:0] : _GEN_12250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13301 = 10'had == _T_31 ? _ram_T_337[287:0] : _GEN_12251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13302 = 10'hae == _T_31 ? _ram_T_337[287:0] : _GEN_12252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13303 = 10'haf == _T_31 ? _ram_T_337[287:0] : _GEN_12253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13304 = 10'hb0 == _T_31 ? _ram_T_337[287:0] : _GEN_12254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13305 = 10'hb1 == _T_31 ? _ram_T_337[287:0] : _GEN_12255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13306 = 10'hb2 == _T_31 ? _ram_T_337[287:0] : _GEN_12256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13307 = 10'hb3 == _T_31 ? _ram_T_337[287:0] : _GEN_12257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13308 = 10'hb4 == _T_31 ? _ram_T_337[287:0] : _GEN_12258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13309 = 10'hb5 == _T_31 ? _ram_T_337[287:0] : _GEN_12259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13310 = 10'hb6 == _T_31 ? _ram_T_337[287:0] : _GEN_12260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13311 = 10'hb7 == _T_31 ? _ram_T_337[287:0] : _GEN_12261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13312 = 10'hb8 == _T_31 ? _ram_T_337[287:0] : _GEN_12262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13313 = 10'hb9 == _T_31 ? _ram_T_337[287:0] : _GEN_12263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13314 = 10'hba == _T_31 ? _ram_T_337[287:0] : _GEN_12264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13315 = 10'hbb == _T_31 ? _ram_T_337[287:0] : _GEN_12265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13316 = 10'hbc == _T_31 ? _ram_T_337[287:0] : _GEN_12266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13317 = 10'hbd == _T_31 ? _ram_T_337[287:0] : _GEN_12267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13318 = 10'hbe == _T_31 ? _ram_T_337[287:0] : _GEN_12268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13319 = 10'hbf == _T_31 ? _ram_T_337[287:0] : _GEN_12269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13320 = 10'hc0 == _T_31 ? _ram_T_337[287:0] : _GEN_12270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13321 = 10'hc1 == _T_31 ? _ram_T_337[287:0] : _GEN_12271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13322 = 10'hc2 == _T_31 ? _ram_T_337[287:0] : _GEN_12272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13323 = 10'hc3 == _T_31 ? _ram_T_337[287:0] : _GEN_12273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13324 = 10'hc4 == _T_31 ? _ram_T_337[287:0] : _GEN_12274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13325 = 10'hc5 == _T_31 ? _ram_T_337[287:0] : _GEN_12275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13326 = 10'hc6 == _T_31 ? _ram_T_337[287:0] : _GEN_12276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13327 = 10'hc7 == _T_31 ? _ram_T_337[287:0] : _GEN_12277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13328 = 10'hc8 == _T_31 ? _ram_T_337[287:0] : _GEN_12278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13329 = 10'hc9 == _T_31 ? _ram_T_337[287:0] : _GEN_12279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13330 = 10'hca == _T_31 ? _ram_T_337[287:0] : _GEN_12280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13331 = 10'hcb == _T_31 ? _ram_T_337[287:0] : _GEN_12281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13332 = 10'hcc == _T_31 ? _ram_T_337[287:0] : _GEN_12282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13333 = 10'hcd == _T_31 ? _ram_T_337[287:0] : _GEN_12283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13334 = 10'hce == _T_31 ? _ram_T_337[287:0] : _GEN_12284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13335 = 10'hcf == _T_31 ? _ram_T_337[287:0] : _GEN_12285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13336 = 10'hd0 == _T_31 ? _ram_T_337[287:0] : _GEN_12286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13337 = 10'hd1 == _T_31 ? _ram_T_337[287:0] : _GEN_12287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13338 = 10'hd2 == _T_31 ? _ram_T_337[287:0] : _GEN_12288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13339 = 10'hd3 == _T_31 ? _ram_T_337[287:0] : _GEN_12289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13340 = 10'hd4 == _T_31 ? _ram_T_337[287:0] : _GEN_12290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13341 = 10'hd5 == _T_31 ? _ram_T_337[287:0] : _GEN_12291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13342 = 10'hd6 == _T_31 ? _ram_T_337[287:0] : _GEN_12292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13343 = 10'hd7 == _T_31 ? _ram_T_337[287:0] : _GEN_12293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13344 = 10'hd8 == _T_31 ? _ram_T_337[287:0] : _GEN_12294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13345 = 10'hd9 == _T_31 ? _ram_T_337[287:0] : _GEN_12295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13346 = 10'hda == _T_31 ? _ram_T_337[287:0] : _GEN_12296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13347 = 10'hdb == _T_31 ? _ram_T_337[287:0] : _GEN_12297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13348 = 10'hdc == _T_31 ? _ram_T_337[287:0] : _GEN_12298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13349 = 10'hdd == _T_31 ? _ram_T_337[287:0] : _GEN_12299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13350 = 10'hde == _T_31 ? _ram_T_337[287:0] : _GEN_12300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13351 = 10'hdf == _T_31 ? _ram_T_337[287:0] : _GEN_12301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13352 = 10'he0 == _T_31 ? _ram_T_337[287:0] : _GEN_12302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13353 = 10'he1 == _T_31 ? _ram_T_337[287:0] : _GEN_12303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13354 = 10'he2 == _T_31 ? _ram_T_337[287:0] : _GEN_12304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13355 = 10'he3 == _T_31 ? _ram_T_337[287:0] : _GEN_12305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13356 = 10'he4 == _T_31 ? _ram_T_337[287:0] : _GEN_12306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13357 = 10'he5 == _T_31 ? _ram_T_337[287:0] : _GEN_12307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13358 = 10'he6 == _T_31 ? _ram_T_337[287:0] : _GEN_12308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13359 = 10'he7 == _T_31 ? _ram_T_337[287:0] : _GEN_12309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13360 = 10'he8 == _T_31 ? _ram_T_337[287:0] : _GEN_12310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13361 = 10'he9 == _T_31 ? _ram_T_337[287:0] : _GEN_12311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13362 = 10'hea == _T_31 ? _ram_T_337[287:0] : _GEN_12312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13363 = 10'heb == _T_31 ? _ram_T_337[287:0] : _GEN_12313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13364 = 10'hec == _T_31 ? _ram_T_337[287:0] : _GEN_12314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13365 = 10'hed == _T_31 ? _ram_T_337[287:0] : _GEN_12315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13366 = 10'hee == _T_31 ? _ram_T_337[287:0] : _GEN_12316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13367 = 10'hef == _T_31 ? _ram_T_337[287:0] : _GEN_12317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13368 = 10'hf0 == _T_31 ? _ram_T_337[287:0] : _GEN_12318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13369 = 10'hf1 == _T_31 ? _ram_T_337[287:0] : _GEN_12319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13370 = 10'hf2 == _T_31 ? _ram_T_337[287:0] : _GEN_12320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13371 = 10'hf3 == _T_31 ? _ram_T_337[287:0] : _GEN_12321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13372 = 10'hf4 == _T_31 ? _ram_T_337[287:0] : _GEN_12322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13373 = 10'hf5 == _T_31 ? _ram_T_337[287:0] : _GEN_12323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13374 = 10'hf6 == _T_31 ? _ram_T_337[287:0] : _GEN_12324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13375 = 10'hf7 == _T_31 ? _ram_T_337[287:0] : _GEN_12325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13376 = 10'hf8 == _T_31 ? _ram_T_337[287:0] : _GEN_12326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13377 = 10'hf9 == _T_31 ? _ram_T_337[287:0] : _GEN_12327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13378 = 10'hfa == _T_31 ? _ram_T_337[287:0] : _GEN_12328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13379 = 10'hfb == _T_31 ? _ram_T_337[287:0] : _GEN_12329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13380 = 10'hfc == _T_31 ? _ram_T_337[287:0] : _GEN_12330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13381 = 10'hfd == _T_31 ? _ram_T_337[287:0] : _GEN_12331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13382 = 10'hfe == _T_31 ? _ram_T_337[287:0] : _GEN_12332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13383 = 10'hff == _T_31 ? _ram_T_337[287:0] : _GEN_12333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13384 = 10'h100 == _T_31 ? _ram_T_337[287:0] : _GEN_12334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13385 = 10'h101 == _T_31 ? _ram_T_337[287:0] : _GEN_12335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13386 = 10'h102 == _T_31 ? _ram_T_337[287:0] : _GEN_12336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13387 = 10'h103 == _T_31 ? _ram_T_337[287:0] : _GEN_12337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13388 = 10'h104 == _T_31 ? _ram_T_337[287:0] : _GEN_12338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13389 = 10'h105 == _T_31 ? _ram_T_337[287:0] : _GEN_12339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13390 = 10'h106 == _T_31 ? _ram_T_337[287:0] : _GEN_12340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13391 = 10'h107 == _T_31 ? _ram_T_337[287:0] : _GEN_12341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13392 = 10'h108 == _T_31 ? _ram_T_337[287:0] : _GEN_12342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13393 = 10'h109 == _T_31 ? _ram_T_337[287:0] : _GEN_12343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13394 = 10'h10a == _T_31 ? _ram_T_337[287:0] : _GEN_12344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13395 = 10'h10b == _T_31 ? _ram_T_337[287:0] : _GEN_12345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13396 = 10'h10c == _T_31 ? _ram_T_337[287:0] : _GEN_12346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13397 = 10'h10d == _T_31 ? _ram_T_337[287:0] : _GEN_12347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13398 = 10'h10e == _T_31 ? _ram_T_337[287:0] : _GEN_12348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13399 = 10'h10f == _T_31 ? _ram_T_337[287:0] : _GEN_12349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13400 = 10'h110 == _T_31 ? _ram_T_337[287:0] : _GEN_12350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13401 = 10'h111 == _T_31 ? _ram_T_337[287:0] : _GEN_12351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13402 = 10'h112 == _T_31 ? _ram_T_337[287:0] : _GEN_12352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13403 = 10'h113 == _T_31 ? _ram_T_337[287:0] : _GEN_12353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13404 = 10'h114 == _T_31 ? _ram_T_337[287:0] : _GEN_12354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13405 = 10'h115 == _T_31 ? _ram_T_337[287:0] : _GEN_12355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13406 = 10'h116 == _T_31 ? _ram_T_337[287:0] : _GEN_12356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13407 = 10'h117 == _T_31 ? _ram_T_337[287:0] : _GEN_12357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13408 = 10'h118 == _T_31 ? _ram_T_337[287:0] : _GEN_12358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13409 = 10'h119 == _T_31 ? _ram_T_337[287:0] : _GEN_12359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13410 = 10'h11a == _T_31 ? _ram_T_337[287:0] : _GEN_12360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13411 = 10'h11b == _T_31 ? _ram_T_337[287:0] : _GEN_12361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13412 = 10'h11c == _T_31 ? _ram_T_337[287:0] : _GEN_12362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13413 = 10'h11d == _T_31 ? _ram_T_337[287:0] : _GEN_12363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13414 = 10'h11e == _T_31 ? _ram_T_337[287:0] : _GEN_12364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13415 = 10'h11f == _T_31 ? _ram_T_337[287:0] : _GEN_12365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13416 = 10'h120 == _T_31 ? _ram_T_337[287:0] : _GEN_12366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13417 = 10'h121 == _T_31 ? _ram_T_337[287:0] : _GEN_12367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13418 = 10'h122 == _T_31 ? _ram_T_337[287:0] : _GEN_12368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13419 = 10'h123 == _T_31 ? _ram_T_337[287:0] : _GEN_12369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13420 = 10'h124 == _T_31 ? _ram_T_337[287:0] : _GEN_12370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13421 = 10'h125 == _T_31 ? _ram_T_337[287:0] : _GEN_12371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13422 = 10'h126 == _T_31 ? _ram_T_337[287:0] : _GEN_12372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13423 = 10'h127 == _T_31 ? _ram_T_337[287:0] : _GEN_12373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13424 = 10'h128 == _T_31 ? _ram_T_337[287:0] : _GEN_12374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13425 = 10'h129 == _T_31 ? _ram_T_337[287:0] : _GEN_12375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13426 = 10'h12a == _T_31 ? _ram_T_337[287:0] : _GEN_12376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13427 = 10'h12b == _T_31 ? _ram_T_337[287:0] : _GEN_12377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13428 = 10'h12c == _T_31 ? _ram_T_337[287:0] : _GEN_12378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13429 = 10'h12d == _T_31 ? _ram_T_337[287:0] : _GEN_12379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13430 = 10'h12e == _T_31 ? _ram_T_337[287:0] : _GEN_12380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13431 = 10'h12f == _T_31 ? _ram_T_337[287:0] : _GEN_12381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13432 = 10'h130 == _T_31 ? _ram_T_337[287:0] : _GEN_12382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13433 = 10'h131 == _T_31 ? _ram_T_337[287:0] : _GEN_12383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13434 = 10'h132 == _T_31 ? _ram_T_337[287:0] : _GEN_12384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13435 = 10'h133 == _T_31 ? _ram_T_337[287:0] : _GEN_12385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13436 = 10'h134 == _T_31 ? _ram_T_337[287:0] : _GEN_12386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13437 = 10'h135 == _T_31 ? _ram_T_337[287:0] : _GEN_12387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13438 = 10'h136 == _T_31 ? _ram_T_337[287:0] : _GEN_12388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13439 = 10'h137 == _T_31 ? _ram_T_337[287:0] : _GEN_12389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13440 = 10'h138 == _T_31 ? _ram_T_337[287:0] : _GEN_12390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13441 = 10'h139 == _T_31 ? _ram_T_337[287:0] : _GEN_12391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13442 = 10'h13a == _T_31 ? _ram_T_337[287:0] : _GEN_12392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13443 = 10'h13b == _T_31 ? _ram_T_337[287:0] : _GEN_12393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13444 = 10'h13c == _T_31 ? _ram_T_337[287:0] : _GEN_12394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13445 = 10'h13d == _T_31 ? _ram_T_337[287:0] : _GEN_12395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13446 = 10'h13e == _T_31 ? _ram_T_337[287:0] : _GEN_12396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13447 = 10'h13f == _T_31 ? _ram_T_337[287:0] : _GEN_12397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13448 = 10'h140 == _T_31 ? _ram_T_337[287:0] : _GEN_12398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13449 = 10'h141 == _T_31 ? _ram_T_337[287:0] : _GEN_12399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13450 = 10'h142 == _T_31 ? _ram_T_337[287:0] : _GEN_12400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13451 = 10'h143 == _T_31 ? _ram_T_337[287:0] : _GEN_12401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13452 = 10'h144 == _T_31 ? _ram_T_337[287:0] : _GEN_12402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13453 = 10'h145 == _T_31 ? _ram_T_337[287:0] : _GEN_12403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13454 = 10'h146 == _T_31 ? _ram_T_337[287:0] : _GEN_12404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13455 = 10'h147 == _T_31 ? _ram_T_337[287:0] : _GEN_12405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13456 = 10'h148 == _T_31 ? _ram_T_337[287:0] : _GEN_12406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13457 = 10'h149 == _T_31 ? _ram_T_337[287:0] : _GEN_12407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13458 = 10'h14a == _T_31 ? _ram_T_337[287:0] : _GEN_12408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13459 = 10'h14b == _T_31 ? _ram_T_337[287:0] : _GEN_12409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13460 = 10'h14c == _T_31 ? _ram_T_337[287:0] : _GEN_12410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13461 = 10'h14d == _T_31 ? _ram_T_337[287:0] : _GEN_12411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13462 = 10'h14e == _T_31 ? _ram_T_337[287:0] : _GEN_12412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13463 = 10'h14f == _T_31 ? _ram_T_337[287:0] : _GEN_12413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13464 = 10'h150 == _T_31 ? _ram_T_337[287:0] : _GEN_12414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13465 = 10'h151 == _T_31 ? _ram_T_337[287:0] : _GEN_12415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13466 = 10'h152 == _T_31 ? _ram_T_337[287:0] : _GEN_12416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13467 = 10'h153 == _T_31 ? _ram_T_337[287:0] : _GEN_12417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13468 = 10'h154 == _T_31 ? _ram_T_337[287:0] : _GEN_12418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13469 = 10'h155 == _T_31 ? _ram_T_337[287:0] : _GEN_12419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13470 = 10'h156 == _T_31 ? _ram_T_337[287:0] : _GEN_12420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13471 = 10'h157 == _T_31 ? _ram_T_337[287:0] : _GEN_12421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13472 = 10'h158 == _T_31 ? _ram_T_337[287:0] : _GEN_12422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13473 = 10'h159 == _T_31 ? _ram_T_337[287:0] : _GEN_12423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13474 = 10'h15a == _T_31 ? _ram_T_337[287:0] : _GEN_12424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13475 = 10'h15b == _T_31 ? _ram_T_337[287:0] : _GEN_12425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13476 = 10'h15c == _T_31 ? _ram_T_337[287:0] : _GEN_12426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13477 = 10'h15d == _T_31 ? _ram_T_337[287:0] : _GEN_12427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13478 = 10'h15e == _T_31 ? _ram_T_337[287:0] : _GEN_12428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13479 = 10'h15f == _T_31 ? _ram_T_337[287:0] : _GEN_12429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13480 = 10'h160 == _T_31 ? _ram_T_337[287:0] : _GEN_12430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13481 = 10'h161 == _T_31 ? _ram_T_337[287:0] : _GEN_12431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13482 = 10'h162 == _T_31 ? _ram_T_337[287:0] : _GEN_12432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13483 = 10'h163 == _T_31 ? _ram_T_337[287:0] : _GEN_12433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13484 = 10'h164 == _T_31 ? _ram_T_337[287:0] : _GEN_12434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13485 = 10'h165 == _T_31 ? _ram_T_337[287:0] : _GEN_12435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13486 = 10'h166 == _T_31 ? _ram_T_337[287:0] : _GEN_12436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13487 = 10'h167 == _T_31 ? _ram_T_337[287:0] : _GEN_12437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13488 = 10'h168 == _T_31 ? _ram_T_337[287:0] : _GEN_12438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13489 = 10'h169 == _T_31 ? _ram_T_337[287:0] : _GEN_12439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13490 = 10'h16a == _T_31 ? _ram_T_337[287:0] : _GEN_12440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13491 = 10'h16b == _T_31 ? _ram_T_337[287:0] : _GEN_12441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13492 = 10'h16c == _T_31 ? _ram_T_337[287:0] : _GEN_12442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13493 = 10'h16d == _T_31 ? _ram_T_337[287:0] : _GEN_12443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13494 = 10'h16e == _T_31 ? _ram_T_337[287:0] : _GEN_12444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13495 = 10'h16f == _T_31 ? _ram_T_337[287:0] : _GEN_12445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13496 = 10'h170 == _T_31 ? _ram_T_337[287:0] : _GEN_12446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13497 = 10'h171 == _T_31 ? _ram_T_337[287:0] : _GEN_12447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13498 = 10'h172 == _T_31 ? _ram_T_337[287:0] : _GEN_12448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13499 = 10'h173 == _T_31 ? _ram_T_337[287:0] : _GEN_12449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13500 = 10'h174 == _T_31 ? _ram_T_337[287:0] : _GEN_12450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13501 = 10'h175 == _T_31 ? _ram_T_337[287:0] : _GEN_12451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13502 = 10'h176 == _T_31 ? _ram_T_337[287:0] : _GEN_12452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13503 = 10'h177 == _T_31 ? _ram_T_337[287:0] : _GEN_12453; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13504 = 10'h178 == _T_31 ? _ram_T_337[287:0] : _GEN_12454; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13505 = 10'h179 == _T_31 ? _ram_T_337[287:0] : _GEN_12455; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13506 = 10'h17a == _T_31 ? _ram_T_337[287:0] : _GEN_12456; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13507 = 10'h17b == _T_31 ? _ram_T_337[287:0] : _GEN_12457; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13508 = 10'h17c == _T_31 ? _ram_T_337[287:0] : _GEN_12458; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13509 = 10'h17d == _T_31 ? _ram_T_337[287:0] : _GEN_12459; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13510 = 10'h17e == _T_31 ? _ram_T_337[287:0] : _GEN_12460; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13511 = 10'h17f == _T_31 ? _ram_T_337[287:0] : _GEN_12461; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13512 = 10'h180 == _T_31 ? _ram_T_337[287:0] : _GEN_12462; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13513 = 10'h181 == _T_31 ? _ram_T_337[287:0] : _GEN_12463; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13514 = 10'h182 == _T_31 ? _ram_T_337[287:0] : _GEN_12464; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13515 = 10'h183 == _T_31 ? _ram_T_337[287:0] : _GEN_12465; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13516 = 10'h184 == _T_31 ? _ram_T_337[287:0] : _GEN_12466; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13517 = 10'h185 == _T_31 ? _ram_T_337[287:0] : _GEN_12467; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13518 = 10'h186 == _T_31 ? _ram_T_337[287:0] : _GEN_12468; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13519 = 10'h187 == _T_31 ? _ram_T_337[287:0] : _GEN_12469; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13520 = 10'h188 == _T_31 ? _ram_T_337[287:0] : _GEN_12470; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13521 = 10'h189 == _T_31 ? _ram_T_337[287:0] : _GEN_12471; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13522 = 10'h18a == _T_31 ? _ram_T_337[287:0] : _GEN_12472; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13523 = 10'h18b == _T_31 ? _ram_T_337[287:0] : _GEN_12473; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13524 = 10'h18c == _T_31 ? _ram_T_337[287:0] : _GEN_12474; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13525 = 10'h18d == _T_31 ? _ram_T_337[287:0] : _GEN_12475; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13526 = 10'h18e == _T_31 ? _ram_T_337[287:0] : _GEN_12476; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13527 = 10'h18f == _T_31 ? _ram_T_337[287:0] : _GEN_12477; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13528 = 10'h190 == _T_31 ? _ram_T_337[287:0] : _GEN_12478; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13529 = 10'h191 == _T_31 ? _ram_T_337[287:0] : _GEN_12479; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13530 = 10'h192 == _T_31 ? _ram_T_337[287:0] : _GEN_12480; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13531 = 10'h193 == _T_31 ? _ram_T_337[287:0] : _GEN_12481; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13532 = 10'h194 == _T_31 ? _ram_T_337[287:0] : _GEN_12482; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13533 = 10'h195 == _T_31 ? _ram_T_337[287:0] : _GEN_12483; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13534 = 10'h196 == _T_31 ? _ram_T_337[287:0] : _GEN_12484; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13535 = 10'h197 == _T_31 ? _ram_T_337[287:0] : _GEN_12485; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13536 = 10'h198 == _T_31 ? _ram_T_337[287:0] : _GEN_12486; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13537 = 10'h199 == _T_31 ? _ram_T_337[287:0] : _GEN_12487; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13538 = 10'h19a == _T_31 ? _ram_T_337[287:0] : _GEN_12488; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13539 = 10'h19b == _T_31 ? _ram_T_337[287:0] : _GEN_12489; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13540 = 10'h19c == _T_31 ? _ram_T_337[287:0] : _GEN_12490; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13541 = 10'h19d == _T_31 ? _ram_T_337[287:0] : _GEN_12491; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13542 = 10'h19e == _T_31 ? _ram_T_337[287:0] : _GEN_12492; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13543 = 10'h19f == _T_31 ? _ram_T_337[287:0] : _GEN_12493; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13544 = 10'h1a0 == _T_31 ? _ram_T_337[287:0] : _GEN_12494; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13545 = 10'h1a1 == _T_31 ? _ram_T_337[287:0] : _GEN_12495; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13546 = 10'h1a2 == _T_31 ? _ram_T_337[287:0] : _GEN_12496; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13547 = 10'h1a3 == _T_31 ? _ram_T_337[287:0] : _GEN_12497; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13548 = 10'h1a4 == _T_31 ? _ram_T_337[287:0] : _GEN_12498; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13549 = 10'h1a5 == _T_31 ? _ram_T_337[287:0] : _GEN_12499; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13550 = 10'h1a6 == _T_31 ? _ram_T_337[287:0] : _GEN_12500; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13551 = 10'h1a7 == _T_31 ? _ram_T_337[287:0] : _GEN_12501; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13552 = 10'h1a8 == _T_31 ? _ram_T_337[287:0] : _GEN_12502; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13553 = 10'h1a9 == _T_31 ? _ram_T_337[287:0] : _GEN_12503; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13554 = 10'h1aa == _T_31 ? _ram_T_337[287:0] : _GEN_12504; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13555 = 10'h1ab == _T_31 ? _ram_T_337[287:0] : _GEN_12505; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13556 = 10'h1ac == _T_31 ? _ram_T_337[287:0] : _GEN_12506; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13557 = 10'h1ad == _T_31 ? _ram_T_337[287:0] : _GEN_12507; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13558 = 10'h1ae == _T_31 ? _ram_T_337[287:0] : _GEN_12508; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13559 = 10'h1af == _T_31 ? _ram_T_337[287:0] : _GEN_12509; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13560 = 10'h1b0 == _T_31 ? _ram_T_337[287:0] : _GEN_12510; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13561 = 10'h1b1 == _T_31 ? _ram_T_337[287:0] : _GEN_12511; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13562 = 10'h1b2 == _T_31 ? _ram_T_337[287:0] : _GEN_12512; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13563 = 10'h1b3 == _T_31 ? _ram_T_337[287:0] : _GEN_12513; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13564 = 10'h1b4 == _T_31 ? _ram_T_337[287:0] : _GEN_12514; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13565 = 10'h1b5 == _T_31 ? _ram_T_337[287:0] : _GEN_12515; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13566 = 10'h1b6 == _T_31 ? _ram_T_337[287:0] : _GEN_12516; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13567 = 10'h1b7 == _T_31 ? _ram_T_337[287:0] : _GEN_12517; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13568 = 10'h1b8 == _T_31 ? _ram_T_337[287:0] : _GEN_12518; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13569 = 10'h1b9 == _T_31 ? _ram_T_337[287:0] : _GEN_12519; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13570 = 10'h1ba == _T_31 ? _ram_T_337[287:0] : _GEN_12520; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13571 = 10'h1bb == _T_31 ? _ram_T_337[287:0] : _GEN_12521; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13572 = 10'h1bc == _T_31 ? _ram_T_337[287:0] : _GEN_12522; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13573 = 10'h1bd == _T_31 ? _ram_T_337[287:0] : _GEN_12523; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13574 = 10'h1be == _T_31 ? _ram_T_337[287:0] : _GEN_12524; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13575 = 10'h1bf == _T_31 ? _ram_T_337[287:0] : _GEN_12525; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13576 = 10'h1c0 == _T_31 ? _ram_T_337[287:0] : _GEN_12526; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13577 = 10'h1c1 == _T_31 ? _ram_T_337[287:0] : _GEN_12527; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13578 = 10'h1c2 == _T_31 ? _ram_T_337[287:0] : _GEN_12528; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13579 = 10'h1c3 == _T_31 ? _ram_T_337[287:0] : _GEN_12529; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13580 = 10'h1c4 == _T_31 ? _ram_T_337[287:0] : _GEN_12530; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13581 = 10'h1c5 == _T_31 ? _ram_T_337[287:0] : _GEN_12531; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13582 = 10'h1c6 == _T_31 ? _ram_T_337[287:0] : _GEN_12532; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13583 = 10'h1c7 == _T_31 ? _ram_T_337[287:0] : _GEN_12533; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13584 = 10'h1c8 == _T_31 ? _ram_T_337[287:0] : _GEN_12534; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13585 = 10'h1c9 == _T_31 ? _ram_T_337[287:0] : _GEN_12535; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13586 = 10'h1ca == _T_31 ? _ram_T_337[287:0] : _GEN_12536; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13587 = 10'h1cb == _T_31 ? _ram_T_337[287:0] : _GEN_12537; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13588 = 10'h1cc == _T_31 ? _ram_T_337[287:0] : _GEN_12538; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13589 = 10'h1cd == _T_31 ? _ram_T_337[287:0] : _GEN_12539; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13590 = 10'h1ce == _T_31 ? _ram_T_337[287:0] : _GEN_12540; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13591 = 10'h1cf == _T_31 ? _ram_T_337[287:0] : _GEN_12541; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13592 = 10'h1d0 == _T_31 ? _ram_T_337[287:0] : _GEN_12542; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13593 = 10'h1d1 == _T_31 ? _ram_T_337[287:0] : _GEN_12543; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13594 = 10'h1d2 == _T_31 ? _ram_T_337[287:0] : _GEN_12544; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13595 = 10'h1d3 == _T_31 ? _ram_T_337[287:0] : _GEN_12545; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13596 = 10'h1d4 == _T_31 ? _ram_T_337[287:0] : _GEN_12546; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13597 = 10'h1d5 == _T_31 ? _ram_T_337[287:0] : _GEN_12547; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13598 = 10'h1d6 == _T_31 ? _ram_T_337[287:0] : _GEN_12548; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13599 = 10'h1d7 == _T_31 ? _ram_T_337[287:0] : _GEN_12549; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13600 = 10'h1d8 == _T_31 ? _ram_T_337[287:0] : _GEN_12550; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13601 = 10'h1d9 == _T_31 ? _ram_T_337[287:0] : _GEN_12551; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13602 = 10'h1da == _T_31 ? _ram_T_337[287:0] : _GEN_12552; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13603 = 10'h1db == _T_31 ? _ram_T_337[287:0] : _GEN_12553; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13604 = 10'h1dc == _T_31 ? _ram_T_337[287:0] : _GEN_12554; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13605 = 10'h1dd == _T_31 ? _ram_T_337[287:0] : _GEN_12555; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13606 = 10'h1de == _T_31 ? _ram_T_337[287:0] : _GEN_12556; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13607 = 10'h1df == _T_31 ? _ram_T_337[287:0] : _GEN_12557; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13608 = 10'h1e0 == _T_31 ? _ram_T_337[287:0] : _GEN_12558; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13609 = 10'h1e1 == _T_31 ? _ram_T_337[287:0] : _GEN_12559; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13610 = 10'h1e2 == _T_31 ? _ram_T_337[287:0] : _GEN_12560; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13611 = 10'h1e3 == _T_31 ? _ram_T_337[287:0] : _GEN_12561; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13612 = 10'h1e4 == _T_31 ? _ram_T_337[287:0] : _GEN_12562; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13613 = 10'h1e5 == _T_31 ? _ram_T_337[287:0] : _GEN_12563; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13614 = 10'h1e6 == _T_31 ? _ram_T_337[287:0] : _GEN_12564; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13615 = 10'h1e7 == _T_31 ? _ram_T_337[287:0] : _GEN_12565; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13616 = 10'h1e8 == _T_31 ? _ram_T_337[287:0] : _GEN_12566; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13617 = 10'h1e9 == _T_31 ? _ram_T_337[287:0] : _GEN_12567; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13618 = 10'h1ea == _T_31 ? _ram_T_337[287:0] : _GEN_12568; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13619 = 10'h1eb == _T_31 ? _ram_T_337[287:0] : _GEN_12569; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13620 = 10'h1ec == _T_31 ? _ram_T_337[287:0] : _GEN_12570; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13621 = 10'h1ed == _T_31 ? _ram_T_337[287:0] : _GEN_12571; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13622 = 10'h1ee == _T_31 ? _ram_T_337[287:0] : _GEN_12572; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13623 = 10'h1ef == _T_31 ? _ram_T_337[287:0] : _GEN_12573; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13624 = 10'h1f0 == _T_31 ? _ram_T_337[287:0] : _GEN_12574; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13625 = 10'h1f1 == _T_31 ? _ram_T_337[287:0] : _GEN_12575; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13626 = 10'h1f2 == _T_31 ? _ram_T_337[287:0] : _GEN_12576; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13627 = 10'h1f3 == _T_31 ? _ram_T_337[287:0] : _GEN_12577; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13628 = 10'h1f4 == _T_31 ? _ram_T_337[287:0] : _GEN_12578; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13629 = 10'h1f5 == _T_31 ? _ram_T_337[287:0] : _GEN_12579; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13630 = 10'h1f6 == _T_31 ? _ram_T_337[287:0] : _GEN_12580; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13631 = 10'h1f7 == _T_31 ? _ram_T_337[287:0] : _GEN_12581; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13632 = 10'h1f8 == _T_31 ? _ram_T_337[287:0] : _GEN_12582; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13633 = 10'h1f9 == _T_31 ? _ram_T_337[287:0] : _GEN_12583; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13634 = 10'h1fa == _T_31 ? _ram_T_337[287:0] : _GEN_12584; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13635 = 10'h1fb == _T_31 ? _ram_T_337[287:0] : _GEN_12585; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13636 = 10'h1fc == _T_31 ? _ram_T_337[287:0] : _GEN_12586; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13637 = 10'h1fd == _T_31 ? _ram_T_337[287:0] : _GEN_12587; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13638 = 10'h1fe == _T_31 ? _ram_T_337[287:0] : _GEN_12588; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13639 = 10'h1ff == _T_31 ? _ram_T_337[287:0] : _GEN_12589; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13640 = 10'h200 == _T_31 ? _ram_T_337[287:0] : _GEN_12590; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13641 = 10'h201 == _T_31 ? _ram_T_337[287:0] : _GEN_12591; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13642 = 10'h202 == _T_31 ? _ram_T_337[287:0] : _GEN_12592; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13643 = 10'h203 == _T_31 ? _ram_T_337[287:0] : _GEN_12593; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13644 = 10'h204 == _T_31 ? _ram_T_337[287:0] : _GEN_12594; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13645 = 10'h205 == _T_31 ? _ram_T_337[287:0] : _GEN_12595; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13646 = 10'h206 == _T_31 ? _ram_T_337[287:0] : _GEN_12596; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13647 = 10'h207 == _T_31 ? _ram_T_337[287:0] : _GEN_12597; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13648 = 10'h208 == _T_31 ? _ram_T_337[287:0] : _GEN_12598; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13649 = 10'h209 == _T_31 ? _ram_T_337[287:0] : _GEN_12599; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13650 = 10'h20a == _T_31 ? _ram_T_337[287:0] : _GEN_12600; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13651 = 10'h20b == _T_31 ? _ram_T_337[287:0] : _GEN_12601; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_13652 = 10'h20c == _T_31 ? _ram_T_337[287:0] : _GEN_12602; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_33 = h + 10'hd; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_13 = vga_mem_ram_MPORT_117_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_13 = vga_mem_ram_MPORT_118_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_13 = vga_mem_ram_MPORT_119_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_13 = vga_mem_ram_MPORT_120_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_13 = vga_mem_ram_MPORT_121_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_13 = vga_mem_ram_MPORT_122_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_13 = vga_mem_ram_MPORT_123_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_13 = vga_mem_ram_MPORT_124_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_13 = vga_mem_ram_MPORT_125_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_358 = {278'h0,ram_hi_hi_hi_lo_13,ram_hi_hi_lo_13,ram_hi_lo_hi_13,ram_hi_lo_lo_13,
    ram_lo_hi_hi_hi_13,ram_lo_hi_hi_lo_13,ram_lo_hi_lo_13,ram_lo_lo_hi_13,ram_lo_lo_lo_13}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19086 = {{8191'd0}, _ram_T_358}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_362 = _GEN_19086 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_13654 = 10'h1 == _T_33 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13655 = 10'h2 == _T_33 ? ram_2 : _GEN_13654; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13656 = 10'h3 == _T_33 ? ram_3 : _GEN_13655; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13657 = 10'h4 == _T_33 ? ram_4 : _GEN_13656; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13658 = 10'h5 == _T_33 ? ram_5 : _GEN_13657; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13659 = 10'h6 == _T_33 ? ram_6 : _GEN_13658; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13660 = 10'h7 == _T_33 ? ram_7 : _GEN_13659; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13661 = 10'h8 == _T_33 ? ram_8 : _GEN_13660; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13662 = 10'h9 == _T_33 ? ram_9 : _GEN_13661; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13663 = 10'ha == _T_33 ? ram_10 : _GEN_13662; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13664 = 10'hb == _T_33 ? ram_11 : _GEN_13663; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13665 = 10'hc == _T_33 ? ram_12 : _GEN_13664; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13666 = 10'hd == _T_33 ? ram_13 : _GEN_13665; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13667 = 10'he == _T_33 ? ram_14 : _GEN_13666; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13668 = 10'hf == _T_33 ? ram_15 : _GEN_13667; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13669 = 10'h10 == _T_33 ? ram_16 : _GEN_13668; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13670 = 10'h11 == _T_33 ? ram_17 : _GEN_13669; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13671 = 10'h12 == _T_33 ? ram_18 : _GEN_13670; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13672 = 10'h13 == _T_33 ? ram_19 : _GEN_13671; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13673 = 10'h14 == _T_33 ? ram_20 : _GEN_13672; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13674 = 10'h15 == _T_33 ? ram_21 : _GEN_13673; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13675 = 10'h16 == _T_33 ? ram_22 : _GEN_13674; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13676 = 10'h17 == _T_33 ? ram_23 : _GEN_13675; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13677 = 10'h18 == _T_33 ? ram_24 : _GEN_13676; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13678 = 10'h19 == _T_33 ? ram_25 : _GEN_13677; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13679 = 10'h1a == _T_33 ? ram_26 : _GEN_13678; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13680 = 10'h1b == _T_33 ? ram_27 : _GEN_13679; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13681 = 10'h1c == _T_33 ? ram_28 : _GEN_13680; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13682 = 10'h1d == _T_33 ? ram_29 : _GEN_13681; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13683 = 10'h1e == _T_33 ? ram_30 : _GEN_13682; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13684 = 10'h1f == _T_33 ? ram_31 : _GEN_13683; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13685 = 10'h20 == _T_33 ? ram_32 : _GEN_13684; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13686 = 10'h21 == _T_33 ? ram_33 : _GEN_13685; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13687 = 10'h22 == _T_33 ? ram_34 : _GEN_13686; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13688 = 10'h23 == _T_33 ? ram_35 : _GEN_13687; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13689 = 10'h24 == _T_33 ? ram_36 : _GEN_13688; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13690 = 10'h25 == _T_33 ? ram_37 : _GEN_13689; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13691 = 10'h26 == _T_33 ? ram_38 : _GEN_13690; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13692 = 10'h27 == _T_33 ? ram_39 : _GEN_13691; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13693 = 10'h28 == _T_33 ? ram_40 : _GEN_13692; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13694 = 10'h29 == _T_33 ? ram_41 : _GEN_13693; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13695 = 10'h2a == _T_33 ? ram_42 : _GEN_13694; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13696 = 10'h2b == _T_33 ? ram_43 : _GEN_13695; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13697 = 10'h2c == _T_33 ? ram_44 : _GEN_13696; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13698 = 10'h2d == _T_33 ? ram_45 : _GEN_13697; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13699 = 10'h2e == _T_33 ? ram_46 : _GEN_13698; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13700 = 10'h2f == _T_33 ? ram_47 : _GEN_13699; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13701 = 10'h30 == _T_33 ? ram_48 : _GEN_13700; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13702 = 10'h31 == _T_33 ? ram_49 : _GEN_13701; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13703 = 10'h32 == _T_33 ? ram_50 : _GEN_13702; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13704 = 10'h33 == _T_33 ? ram_51 : _GEN_13703; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13705 = 10'h34 == _T_33 ? ram_52 : _GEN_13704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13706 = 10'h35 == _T_33 ? ram_53 : _GEN_13705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13707 = 10'h36 == _T_33 ? ram_54 : _GEN_13706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13708 = 10'h37 == _T_33 ? ram_55 : _GEN_13707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13709 = 10'h38 == _T_33 ? ram_56 : _GEN_13708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13710 = 10'h39 == _T_33 ? ram_57 : _GEN_13709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13711 = 10'h3a == _T_33 ? ram_58 : _GEN_13710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13712 = 10'h3b == _T_33 ? ram_59 : _GEN_13711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13713 = 10'h3c == _T_33 ? ram_60 : _GEN_13712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13714 = 10'h3d == _T_33 ? ram_61 : _GEN_13713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13715 = 10'h3e == _T_33 ? ram_62 : _GEN_13714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13716 = 10'h3f == _T_33 ? ram_63 : _GEN_13715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13717 = 10'h40 == _T_33 ? ram_64 : _GEN_13716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13718 = 10'h41 == _T_33 ? ram_65 : _GEN_13717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13719 = 10'h42 == _T_33 ? ram_66 : _GEN_13718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13720 = 10'h43 == _T_33 ? ram_67 : _GEN_13719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13721 = 10'h44 == _T_33 ? ram_68 : _GEN_13720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13722 = 10'h45 == _T_33 ? ram_69 : _GEN_13721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13723 = 10'h46 == _T_33 ? ram_70 : _GEN_13722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13724 = 10'h47 == _T_33 ? ram_71 : _GEN_13723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13725 = 10'h48 == _T_33 ? ram_72 : _GEN_13724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13726 = 10'h49 == _T_33 ? ram_73 : _GEN_13725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13727 = 10'h4a == _T_33 ? ram_74 : _GEN_13726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13728 = 10'h4b == _T_33 ? ram_75 : _GEN_13727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13729 = 10'h4c == _T_33 ? ram_76 : _GEN_13728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13730 = 10'h4d == _T_33 ? ram_77 : _GEN_13729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13731 = 10'h4e == _T_33 ? ram_78 : _GEN_13730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13732 = 10'h4f == _T_33 ? ram_79 : _GEN_13731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13733 = 10'h50 == _T_33 ? ram_80 : _GEN_13732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13734 = 10'h51 == _T_33 ? ram_81 : _GEN_13733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13735 = 10'h52 == _T_33 ? ram_82 : _GEN_13734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13736 = 10'h53 == _T_33 ? ram_83 : _GEN_13735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13737 = 10'h54 == _T_33 ? ram_84 : _GEN_13736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13738 = 10'h55 == _T_33 ? ram_85 : _GEN_13737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13739 = 10'h56 == _T_33 ? ram_86 : _GEN_13738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13740 = 10'h57 == _T_33 ? ram_87 : _GEN_13739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13741 = 10'h58 == _T_33 ? ram_88 : _GEN_13740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13742 = 10'h59 == _T_33 ? ram_89 : _GEN_13741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13743 = 10'h5a == _T_33 ? ram_90 : _GEN_13742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13744 = 10'h5b == _T_33 ? ram_91 : _GEN_13743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13745 = 10'h5c == _T_33 ? ram_92 : _GEN_13744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13746 = 10'h5d == _T_33 ? ram_93 : _GEN_13745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13747 = 10'h5e == _T_33 ? ram_94 : _GEN_13746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13748 = 10'h5f == _T_33 ? ram_95 : _GEN_13747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13749 = 10'h60 == _T_33 ? ram_96 : _GEN_13748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13750 = 10'h61 == _T_33 ? ram_97 : _GEN_13749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13751 = 10'h62 == _T_33 ? ram_98 : _GEN_13750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13752 = 10'h63 == _T_33 ? ram_99 : _GEN_13751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13753 = 10'h64 == _T_33 ? ram_100 : _GEN_13752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13754 = 10'h65 == _T_33 ? ram_101 : _GEN_13753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13755 = 10'h66 == _T_33 ? ram_102 : _GEN_13754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13756 = 10'h67 == _T_33 ? ram_103 : _GEN_13755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13757 = 10'h68 == _T_33 ? ram_104 : _GEN_13756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13758 = 10'h69 == _T_33 ? ram_105 : _GEN_13757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13759 = 10'h6a == _T_33 ? ram_106 : _GEN_13758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13760 = 10'h6b == _T_33 ? ram_107 : _GEN_13759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13761 = 10'h6c == _T_33 ? ram_108 : _GEN_13760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13762 = 10'h6d == _T_33 ? ram_109 : _GEN_13761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13763 = 10'h6e == _T_33 ? ram_110 : _GEN_13762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13764 = 10'h6f == _T_33 ? ram_111 : _GEN_13763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13765 = 10'h70 == _T_33 ? ram_112 : _GEN_13764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13766 = 10'h71 == _T_33 ? ram_113 : _GEN_13765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13767 = 10'h72 == _T_33 ? ram_114 : _GEN_13766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13768 = 10'h73 == _T_33 ? ram_115 : _GEN_13767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13769 = 10'h74 == _T_33 ? ram_116 : _GEN_13768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13770 = 10'h75 == _T_33 ? ram_117 : _GEN_13769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13771 = 10'h76 == _T_33 ? ram_118 : _GEN_13770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13772 = 10'h77 == _T_33 ? ram_119 : _GEN_13771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13773 = 10'h78 == _T_33 ? ram_120 : _GEN_13772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13774 = 10'h79 == _T_33 ? ram_121 : _GEN_13773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13775 = 10'h7a == _T_33 ? ram_122 : _GEN_13774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13776 = 10'h7b == _T_33 ? ram_123 : _GEN_13775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13777 = 10'h7c == _T_33 ? ram_124 : _GEN_13776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13778 = 10'h7d == _T_33 ? ram_125 : _GEN_13777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13779 = 10'h7e == _T_33 ? ram_126 : _GEN_13778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13780 = 10'h7f == _T_33 ? ram_127 : _GEN_13779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13781 = 10'h80 == _T_33 ? ram_128 : _GEN_13780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13782 = 10'h81 == _T_33 ? ram_129 : _GEN_13781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13783 = 10'h82 == _T_33 ? ram_130 : _GEN_13782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13784 = 10'h83 == _T_33 ? ram_131 : _GEN_13783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13785 = 10'h84 == _T_33 ? ram_132 : _GEN_13784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13786 = 10'h85 == _T_33 ? ram_133 : _GEN_13785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13787 = 10'h86 == _T_33 ? ram_134 : _GEN_13786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13788 = 10'h87 == _T_33 ? ram_135 : _GEN_13787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13789 = 10'h88 == _T_33 ? ram_136 : _GEN_13788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13790 = 10'h89 == _T_33 ? ram_137 : _GEN_13789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13791 = 10'h8a == _T_33 ? ram_138 : _GEN_13790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13792 = 10'h8b == _T_33 ? ram_139 : _GEN_13791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13793 = 10'h8c == _T_33 ? ram_140 : _GEN_13792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13794 = 10'h8d == _T_33 ? ram_141 : _GEN_13793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13795 = 10'h8e == _T_33 ? ram_142 : _GEN_13794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13796 = 10'h8f == _T_33 ? ram_143 : _GEN_13795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13797 = 10'h90 == _T_33 ? ram_144 : _GEN_13796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13798 = 10'h91 == _T_33 ? ram_145 : _GEN_13797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13799 = 10'h92 == _T_33 ? ram_146 : _GEN_13798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13800 = 10'h93 == _T_33 ? ram_147 : _GEN_13799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13801 = 10'h94 == _T_33 ? ram_148 : _GEN_13800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13802 = 10'h95 == _T_33 ? ram_149 : _GEN_13801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13803 = 10'h96 == _T_33 ? ram_150 : _GEN_13802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13804 = 10'h97 == _T_33 ? ram_151 : _GEN_13803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13805 = 10'h98 == _T_33 ? ram_152 : _GEN_13804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13806 = 10'h99 == _T_33 ? ram_153 : _GEN_13805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13807 = 10'h9a == _T_33 ? ram_154 : _GEN_13806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13808 = 10'h9b == _T_33 ? ram_155 : _GEN_13807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13809 = 10'h9c == _T_33 ? ram_156 : _GEN_13808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13810 = 10'h9d == _T_33 ? ram_157 : _GEN_13809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13811 = 10'h9e == _T_33 ? ram_158 : _GEN_13810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13812 = 10'h9f == _T_33 ? ram_159 : _GEN_13811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13813 = 10'ha0 == _T_33 ? ram_160 : _GEN_13812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13814 = 10'ha1 == _T_33 ? ram_161 : _GEN_13813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13815 = 10'ha2 == _T_33 ? ram_162 : _GEN_13814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13816 = 10'ha3 == _T_33 ? ram_163 : _GEN_13815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13817 = 10'ha4 == _T_33 ? ram_164 : _GEN_13816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13818 = 10'ha5 == _T_33 ? ram_165 : _GEN_13817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13819 = 10'ha6 == _T_33 ? ram_166 : _GEN_13818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13820 = 10'ha7 == _T_33 ? ram_167 : _GEN_13819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13821 = 10'ha8 == _T_33 ? ram_168 : _GEN_13820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13822 = 10'ha9 == _T_33 ? ram_169 : _GEN_13821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13823 = 10'haa == _T_33 ? ram_170 : _GEN_13822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13824 = 10'hab == _T_33 ? ram_171 : _GEN_13823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13825 = 10'hac == _T_33 ? ram_172 : _GEN_13824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13826 = 10'had == _T_33 ? ram_173 : _GEN_13825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13827 = 10'hae == _T_33 ? ram_174 : _GEN_13826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13828 = 10'haf == _T_33 ? ram_175 : _GEN_13827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13829 = 10'hb0 == _T_33 ? ram_176 : _GEN_13828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13830 = 10'hb1 == _T_33 ? ram_177 : _GEN_13829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13831 = 10'hb2 == _T_33 ? ram_178 : _GEN_13830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13832 = 10'hb3 == _T_33 ? ram_179 : _GEN_13831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13833 = 10'hb4 == _T_33 ? ram_180 : _GEN_13832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13834 = 10'hb5 == _T_33 ? ram_181 : _GEN_13833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13835 = 10'hb6 == _T_33 ? ram_182 : _GEN_13834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13836 = 10'hb7 == _T_33 ? ram_183 : _GEN_13835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13837 = 10'hb8 == _T_33 ? ram_184 : _GEN_13836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13838 = 10'hb9 == _T_33 ? ram_185 : _GEN_13837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13839 = 10'hba == _T_33 ? ram_186 : _GEN_13838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13840 = 10'hbb == _T_33 ? ram_187 : _GEN_13839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13841 = 10'hbc == _T_33 ? ram_188 : _GEN_13840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13842 = 10'hbd == _T_33 ? ram_189 : _GEN_13841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13843 = 10'hbe == _T_33 ? ram_190 : _GEN_13842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13844 = 10'hbf == _T_33 ? ram_191 : _GEN_13843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13845 = 10'hc0 == _T_33 ? ram_192 : _GEN_13844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13846 = 10'hc1 == _T_33 ? ram_193 : _GEN_13845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13847 = 10'hc2 == _T_33 ? ram_194 : _GEN_13846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13848 = 10'hc3 == _T_33 ? ram_195 : _GEN_13847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13849 = 10'hc4 == _T_33 ? ram_196 : _GEN_13848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13850 = 10'hc5 == _T_33 ? ram_197 : _GEN_13849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13851 = 10'hc6 == _T_33 ? ram_198 : _GEN_13850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13852 = 10'hc7 == _T_33 ? ram_199 : _GEN_13851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13853 = 10'hc8 == _T_33 ? ram_200 : _GEN_13852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13854 = 10'hc9 == _T_33 ? ram_201 : _GEN_13853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13855 = 10'hca == _T_33 ? ram_202 : _GEN_13854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13856 = 10'hcb == _T_33 ? ram_203 : _GEN_13855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13857 = 10'hcc == _T_33 ? ram_204 : _GEN_13856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13858 = 10'hcd == _T_33 ? ram_205 : _GEN_13857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13859 = 10'hce == _T_33 ? ram_206 : _GEN_13858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13860 = 10'hcf == _T_33 ? ram_207 : _GEN_13859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13861 = 10'hd0 == _T_33 ? ram_208 : _GEN_13860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13862 = 10'hd1 == _T_33 ? ram_209 : _GEN_13861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13863 = 10'hd2 == _T_33 ? ram_210 : _GEN_13862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13864 = 10'hd3 == _T_33 ? ram_211 : _GEN_13863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13865 = 10'hd4 == _T_33 ? ram_212 : _GEN_13864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13866 = 10'hd5 == _T_33 ? ram_213 : _GEN_13865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13867 = 10'hd6 == _T_33 ? ram_214 : _GEN_13866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13868 = 10'hd7 == _T_33 ? ram_215 : _GEN_13867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13869 = 10'hd8 == _T_33 ? ram_216 : _GEN_13868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13870 = 10'hd9 == _T_33 ? ram_217 : _GEN_13869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13871 = 10'hda == _T_33 ? ram_218 : _GEN_13870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13872 = 10'hdb == _T_33 ? ram_219 : _GEN_13871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13873 = 10'hdc == _T_33 ? ram_220 : _GEN_13872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13874 = 10'hdd == _T_33 ? ram_221 : _GEN_13873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13875 = 10'hde == _T_33 ? ram_222 : _GEN_13874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13876 = 10'hdf == _T_33 ? ram_223 : _GEN_13875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13877 = 10'he0 == _T_33 ? ram_224 : _GEN_13876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13878 = 10'he1 == _T_33 ? ram_225 : _GEN_13877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13879 = 10'he2 == _T_33 ? ram_226 : _GEN_13878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13880 = 10'he3 == _T_33 ? ram_227 : _GEN_13879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13881 = 10'he4 == _T_33 ? ram_228 : _GEN_13880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13882 = 10'he5 == _T_33 ? ram_229 : _GEN_13881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13883 = 10'he6 == _T_33 ? ram_230 : _GEN_13882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13884 = 10'he7 == _T_33 ? ram_231 : _GEN_13883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13885 = 10'he8 == _T_33 ? ram_232 : _GEN_13884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13886 = 10'he9 == _T_33 ? ram_233 : _GEN_13885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13887 = 10'hea == _T_33 ? ram_234 : _GEN_13886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13888 = 10'heb == _T_33 ? ram_235 : _GEN_13887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13889 = 10'hec == _T_33 ? ram_236 : _GEN_13888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13890 = 10'hed == _T_33 ? ram_237 : _GEN_13889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13891 = 10'hee == _T_33 ? ram_238 : _GEN_13890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13892 = 10'hef == _T_33 ? ram_239 : _GEN_13891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13893 = 10'hf0 == _T_33 ? ram_240 : _GEN_13892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13894 = 10'hf1 == _T_33 ? ram_241 : _GEN_13893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13895 = 10'hf2 == _T_33 ? ram_242 : _GEN_13894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13896 = 10'hf3 == _T_33 ? ram_243 : _GEN_13895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13897 = 10'hf4 == _T_33 ? ram_244 : _GEN_13896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13898 = 10'hf5 == _T_33 ? ram_245 : _GEN_13897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13899 = 10'hf6 == _T_33 ? ram_246 : _GEN_13898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13900 = 10'hf7 == _T_33 ? ram_247 : _GEN_13899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13901 = 10'hf8 == _T_33 ? ram_248 : _GEN_13900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13902 = 10'hf9 == _T_33 ? ram_249 : _GEN_13901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13903 = 10'hfa == _T_33 ? ram_250 : _GEN_13902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13904 = 10'hfb == _T_33 ? ram_251 : _GEN_13903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13905 = 10'hfc == _T_33 ? ram_252 : _GEN_13904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13906 = 10'hfd == _T_33 ? ram_253 : _GEN_13905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13907 = 10'hfe == _T_33 ? ram_254 : _GEN_13906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13908 = 10'hff == _T_33 ? ram_255 : _GEN_13907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13909 = 10'h100 == _T_33 ? ram_256 : _GEN_13908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13910 = 10'h101 == _T_33 ? ram_257 : _GEN_13909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13911 = 10'h102 == _T_33 ? ram_258 : _GEN_13910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13912 = 10'h103 == _T_33 ? ram_259 : _GEN_13911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13913 = 10'h104 == _T_33 ? ram_260 : _GEN_13912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13914 = 10'h105 == _T_33 ? ram_261 : _GEN_13913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13915 = 10'h106 == _T_33 ? ram_262 : _GEN_13914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13916 = 10'h107 == _T_33 ? ram_263 : _GEN_13915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13917 = 10'h108 == _T_33 ? ram_264 : _GEN_13916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13918 = 10'h109 == _T_33 ? ram_265 : _GEN_13917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13919 = 10'h10a == _T_33 ? ram_266 : _GEN_13918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13920 = 10'h10b == _T_33 ? ram_267 : _GEN_13919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13921 = 10'h10c == _T_33 ? ram_268 : _GEN_13920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13922 = 10'h10d == _T_33 ? ram_269 : _GEN_13921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13923 = 10'h10e == _T_33 ? ram_270 : _GEN_13922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13924 = 10'h10f == _T_33 ? ram_271 : _GEN_13923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13925 = 10'h110 == _T_33 ? ram_272 : _GEN_13924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13926 = 10'h111 == _T_33 ? ram_273 : _GEN_13925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13927 = 10'h112 == _T_33 ? ram_274 : _GEN_13926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13928 = 10'h113 == _T_33 ? ram_275 : _GEN_13927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13929 = 10'h114 == _T_33 ? ram_276 : _GEN_13928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13930 = 10'h115 == _T_33 ? ram_277 : _GEN_13929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13931 = 10'h116 == _T_33 ? ram_278 : _GEN_13930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13932 = 10'h117 == _T_33 ? ram_279 : _GEN_13931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13933 = 10'h118 == _T_33 ? ram_280 : _GEN_13932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13934 = 10'h119 == _T_33 ? ram_281 : _GEN_13933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13935 = 10'h11a == _T_33 ? ram_282 : _GEN_13934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13936 = 10'h11b == _T_33 ? ram_283 : _GEN_13935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13937 = 10'h11c == _T_33 ? ram_284 : _GEN_13936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13938 = 10'h11d == _T_33 ? ram_285 : _GEN_13937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13939 = 10'h11e == _T_33 ? ram_286 : _GEN_13938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13940 = 10'h11f == _T_33 ? ram_287 : _GEN_13939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13941 = 10'h120 == _T_33 ? ram_288 : _GEN_13940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13942 = 10'h121 == _T_33 ? ram_289 : _GEN_13941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13943 = 10'h122 == _T_33 ? ram_290 : _GEN_13942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13944 = 10'h123 == _T_33 ? ram_291 : _GEN_13943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13945 = 10'h124 == _T_33 ? ram_292 : _GEN_13944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13946 = 10'h125 == _T_33 ? ram_293 : _GEN_13945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13947 = 10'h126 == _T_33 ? ram_294 : _GEN_13946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13948 = 10'h127 == _T_33 ? ram_295 : _GEN_13947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13949 = 10'h128 == _T_33 ? ram_296 : _GEN_13948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13950 = 10'h129 == _T_33 ? ram_297 : _GEN_13949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13951 = 10'h12a == _T_33 ? ram_298 : _GEN_13950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13952 = 10'h12b == _T_33 ? ram_299 : _GEN_13951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13953 = 10'h12c == _T_33 ? ram_300 : _GEN_13952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13954 = 10'h12d == _T_33 ? ram_301 : _GEN_13953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13955 = 10'h12e == _T_33 ? ram_302 : _GEN_13954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13956 = 10'h12f == _T_33 ? ram_303 : _GEN_13955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13957 = 10'h130 == _T_33 ? ram_304 : _GEN_13956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13958 = 10'h131 == _T_33 ? ram_305 : _GEN_13957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13959 = 10'h132 == _T_33 ? ram_306 : _GEN_13958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13960 = 10'h133 == _T_33 ? ram_307 : _GEN_13959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13961 = 10'h134 == _T_33 ? ram_308 : _GEN_13960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13962 = 10'h135 == _T_33 ? ram_309 : _GEN_13961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13963 = 10'h136 == _T_33 ? ram_310 : _GEN_13962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13964 = 10'h137 == _T_33 ? ram_311 : _GEN_13963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13965 = 10'h138 == _T_33 ? ram_312 : _GEN_13964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13966 = 10'h139 == _T_33 ? ram_313 : _GEN_13965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13967 = 10'h13a == _T_33 ? ram_314 : _GEN_13966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13968 = 10'h13b == _T_33 ? ram_315 : _GEN_13967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13969 = 10'h13c == _T_33 ? ram_316 : _GEN_13968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13970 = 10'h13d == _T_33 ? ram_317 : _GEN_13969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13971 = 10'h13e == _T_33 ? ram_318 : _GEN_13970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13972 = 10'h13f == _T_33 ? ram_319 : _GEN_13971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13973 = 10'h140 == _T_33 ? ram_320 : _GEN_13972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13974 = 10'h141 == _T_33 ? ram_321 : _GEN_13973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13975 = 10'h142 == _T_33 ? ram_322 : _GEN_13974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13976 = 10'h143 == _T_33 ? ram_323 : _GEN_13975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13977 = 10'h144 == _T_33 ? ram_324 : _GEN_13976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13978 = 10'h145 == _T_33 ? ram_325 : _GEN_13977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13979 = 10'h146 == _T_33 ? ram_326 : _GEN_13978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13980 = 10'h147 == _T_33 ? ram_327 : _GEN_13979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13981 = 10'h148 == _T_33 ? ram_328 : _GEN_13980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13982 = 10'h149 == _T_33 ? ram_329 : _GEN_13981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13983 = 10'h14a == _T_33 ? ram_330 : _GEN_13982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13984 = 10'h14b == _T_33 ? ram_331 : _GEN_13983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13985 = 10'h14c == _T_33 ? ram_332 : _GEN_13984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13986 = 10'h14d == _T_33 ? ram_333 : _GEN_13985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13987 = 10'h14e == _T_33 ? ram_334 : _GEN_13986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13988 = 10'h14f == _T_33 ? ram_335 : _GEN_13987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13989 = 10'h150 == _T_33 ? ram_336 : _GEN_13988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13990 = 10'h151 == _T_33 ? ram_337 : _GEN_13989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13991 = 10'h152 == _T_33 ? ram_338 : _GEN_13990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13992 = 10'h153 == _T_33 ? ram_339 : _GEN_13991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13993 = 10'h154 == _T_33 ? ram_340 : _GEN_13992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13994 = 10'h155 == _T_33 ? ram_341 : _GEN_13993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13995 = 10'h156 == _T_33 ? ram_342 : _GEN_13994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13996 = 10'h157 == _T_33 ? ram_343 : _GEN_13995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13997 = 10'h158 == _T_33 ? ram_344 : _GEN_13996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13998 = 10'h159 == _T_33 ? ram_345 : _GEN_13997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_13999 = 10'h15a == _T_33 ? ram_346 : _GEN_13998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14000 = 10'h15b == _T_33 ? ram_347 : _GEN_13999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14001 = 10'h15c == _T_33 ? ram_348 : _GEN_14000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14002 = 10'h15d == _T_33 ? ram_349 : _GEN_14001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14003 = 10'h15e == _T_33 ? ram_350 : _GEN_14002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14004 = 10'h15f == _T_33 ? ram_351 : _GEN_14003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14005 = 10'h160 == _T_33 ? ram_352 : _GEN_14004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14006 = 10'h161 == _T_33 ? ram_353 : _GEN_14005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14007 = 10'h162 == _T_33 ? ram_354 : _GEN_14006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14008 = 10'h163 == _T_33 ? ram_355 : _GEN_14007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14009 = 10'h164 == _T_33 ? ram_356 : _GEN_14008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14010 = 10'h165 == _T_33 ? ram_357 : _GEN_14009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14011 = 10'h166 == _T_33 ? ram_358 : _GEN_14010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14012 = 10'h167 == _T_33 ? ram_359 : _GEN_14011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14013 = 10'h168 == _T_33 ? ram_360 : _GEN_14012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14014 = 10'h169 == _T_33 ? ram_361 : _GEN_14013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14015 = 10'h16a == _T_33 ? ram_362 : _GEN_14014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14016 = 10'h16b == _T_33 ? ram_363 : _GEN_14015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14017 = 10'h16c == _T_33 ? ram_364 : _GEN_14016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14018 = 10'h16d == _T_33 ? ram_365 : _GEN_14017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14019 = 10'h16e == _T_33 ? ram_366 : _GEN_14018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14020 = 10'h16f == _T_33 ? ram_367 : _GEN_14019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14021 = 10'h170 == _T_33 ? ram_368 : _GEN_14020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14022 = 10'h171 == _T_33 ? ram_369 : _GEN_14021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14023 = 10'h172 == _T_33 ? ram_370 : _GEN_14022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14024 = 10'h173 == _T_33 ? ram_371 : _GEN_14023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14025 = 10'h174 == _T_33 ? ram_372 : _GEN_14024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14026 = 10'h175 == _T_33 ? ram_373 : _GEN_14025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14027 = 10'h176 == _T_33 ? ram_374 : _GEN_14026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14028 = 10'h177 == _T_33 ? ram_375 : _GEN_14027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14029 = 10'h178 == _T_33 ? ram_376 : _GEN_14028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14030 = 10'h179 == _T_33 ? ram_377 : _GEN_14029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14031 = 10'h17a == _T_33 ? ram_378 : _GEN_14030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14032 = 10'h17b == _T_33 ? ram_379 : _GEN_14031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14033 = 10'h17c == _T_33 ? ram_380 : _GEN_14032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14034 = 10'h17d == _T_33 ? ram_381 : _GEN_14033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14035 = 10'h17e == _T_33 ? ram_382 : _GEN_14034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14036 = 10'h17f == _T_33 ? ram_383 : _GEN_14035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14037 = 10'h180 == _T_33 ? ram_384 : _GEN_14036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14038 = 10'h181 == _T_33 ? ram_385 : _GEN_14037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14039 = 10'h182 == _T_33 ? ram_386 : _GEN_14038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14040 = 10'h183 == _T_33 ? ram_387 : _GEN_14039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14041 = 10'h184 == _T_33 ? ram_388 : _GEN_14040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14042 = 10'h185 == _T_33 ? ram_389 : _GEN_14041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14043 = 10'h186 == _T_33 ? ram_390 : _GEN_14042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14044 = 10'h187 == _T_33 ? ram_391 : _GEN_14043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14045 = 10'h188 == _T_33 ? ram_392 : _GEN_14044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14046 = 10'h189 == _T_33 ? ram_393 : _GEN_14045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14047 = 10'h18a == _T_33 ? ram_394 : _GEN_14046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14048 = 10'h18b == _T_33 ? ram_395 : _GEN_14047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14049 = 10'h18c == _T_33 ? ram_396 : _GEN_14048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14050 = 10'h18d == _T_33 ? ram_397 : _GEN_14049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14051 = 10'h18e == _T_33 ? ram_398 : _GEN_14050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14052 = 10'h18f == _T_33 ? ram_399 : _GEN_14051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14053 = 10'h190 == _T_33 ? ram_400 : _GEN_14052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14054 = 10'h191 == _T_33 ? ram_401 : _GEN_14053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14055 = 10'h192 == _T_33 ? ram_402 : _GEN_14054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14056 = 10'h193 == _T_33 ? ram_403 : _GEN_14055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14057 = 10'h194 == _T_33 ? ram_404 : _GEN_14056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14058 = 10'h195 == _T_33 ? ram_405 : _GEN_14057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14059 = 10'h196 == _T_33 ? ram_406 : _GEN_14058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14060 = 10'h197 == _T_33 ? ram_407 : _GEN_14059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14061 = 10'h198 == _T_33 ? ram_408 : _GEN_14060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14062 = 10'h199 == _T_33 ? ram_409 : _GEN_14061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14063 = 10'h19a == _T_33 ? ram_410 : _GEN_14062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14064 = 10'h19b == _T_33 ? ram_411 : _GEN_14063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14065 = 10'h19c == _T_33 ? ram_412 : _GEN_14064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14066 = 10'h19d == _T_33 ? ram_413 : _GEN_14065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14067 = 10'h19e == _T_33 ? ram_414 : _GEN_14066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14068 = 10'h19f == _T_33 ? ram_415 : _GEN_14067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14069 = 10'h1a0 == _T_33 ? ram_416 : _GEN_14068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14070 = 10'h1a1 == _T_33 ? ram_417 : _GEN_14069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14071 = 10'h1a2 == _T_33 ? ram_418 : _GEN_14070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14072 = 10'h1a3 == _T_33 ? ram_419 : _GEN_14071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14073 = 10'h1a4 == _T_33 ? ram_420 : _GEN_14072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14074 = 10'h1a5 == _T_33 ? ram_421 : _GEN_14073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14075 = 10'h1a6 == _T_33 ? ram_422 : _GEN_14074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14076 = 10'h1a7 == _T_33 ? ram_423 : _GEN_14075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14077 = 10'h1a8 == _T_33 ? ram_424 : _GEN_14076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14078 = 10'h1a9 == _T_33 ? ram_425 : _GEN_14077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14079 = 10'h1aa == _T_33 ? ram_426 : _GEN_14078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14080 = 10'h1ab == _T_33 ? ram_427 : _GEN_14079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14081 = 10'h1ac == _T_33 ? ram_428 : _GEN_14080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14082 = 10'h1ad == _T_33 ? ram_429 : _GEN_14081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14083 = 10'h1ae == _T_33 ? ram_430 : _GEN_14082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14084 = 10'h1af == _T_33 ? ram_431 : _GEN_14083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14085 = 10'h1b0 == _T_33 ? ram_432 : _GEN_14084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14086 = 10'h1b1 == _T_33 ? ram_433 : _GEN_14085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14087 = 10'h1b2 == _T_33 ? ram_434 : _GEN_14086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14088 = 10'h1b3 == _T_33 ? ram_435 : _GEN_14087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14089 = 10'h1b4 == _T_33 ? ram_436 : _GEN_14088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14090 = 10'h1b5 == _T_33 ? ram_437 : _GEN_14089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14091 = 10'h1b6 == _T_33 ? ram_438 : _GEN_14090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14092 = 10'h1b7 == _T_33 ? ram_439 : _GEN_14091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14093 = 10'h1b8 == _T_33 ? ram_440 : _GEN_14092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14094 = 10'h1b9 == _T_33 ? ram_441 : _GEN_14093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14095 = 10'h1ba == _T_33 ? ram_442 : _GEN_14094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14096 = 10'h1bb == _T_33 ? ram_443 : _GEN_14095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14097 = 10'h1bc == _T_33 ? ram_444 : _GEN_14096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14098 = 10'h1bd == _T_33 ? ram_445 : _GEN_14097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14099 = 10'h1be == _T_33 ? ram_446 : _GEN_14098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14100 = 10'h1bf == _T_33 ? ram_447 : _GEN_14099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14101 = 10'h1c0 == _T_33 ? ram_448 : _GEN_14100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14102 = 10'h1c1 == _T_33 ? ram_449 : _GEN_14101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14103 = 10'h1c2 == _T_33 ? ram_450 : _GEN_14102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14104 = 10'h1c3 == _T_33 ? ram_451 : _GEN_14103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14105 = 10'h1c4 == _T_33 ? ram_452 : _GEN_14104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14106 = 10'h1c5 == _T_33 ? ram_453 : _GEN_14105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14107 = 10'h1c6 == _T_33 ? ram_454 : _GEN_14106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14108 = 10'h1c7 == _T_33 ? ram_455 : _GEN_14107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14109 = 10'h1c8 == _T_33 ? ram_456 : _GEN_14108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14110 = 10'h1c9 == _T_33 ? ram_457 : _GEN_14109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14111 = 10'h1ca == _T_33 ? ram_458 : _GEN_14110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14112 = 10'h1cb == _T_33 ? ram_459 : _GEN_14111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14113 = 10'h1cc == _T_33 ? ram_460 : _GEN_14112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14114 = 10'h1cd == _T_33 ? ram_461 : _GEN_14113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14115 = 10'h1ce == _T_33 ? ram_462 : _GEN_14114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14116 = 10'h1cf == _T_33 ? ram_463 : _GEN_14115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14117 = 10'h1d0 == _T_33 ? ram_464 : _GEN_14116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14118 = 10'h1d1 == _T_33 ? ram_465 : _GEN_14117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14119 = 10'h1d2 == _T_33 ? ram_466 : _GEN_14118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14120 = 10'h1d3 == _T_33 ? ram_467 : _GEN_14119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14121 = 10'h1d4 == _T_33 ? ram_468 : _GEN_14120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14122 = 10'h1d5 == _T_33 ? ram_469 : _GEN_14121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14123 = 10'h1d6 == _T_33 ? ram_470 : _GEN_14122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14124 = 10'h1d7 == _T_33 ? ram_471 : _GEN_14123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14125 = 10'h1d8 == _T_33 ? ram_472 : _GEN_14124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14126 = 10'h1d9 == _T_33 ? ram_473 : _GEN_14125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14127 = 10'h1da == _T_33 ? ram_474 : _GEN_14126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14128 = 10'h1db == _T_33 ? ram_475 : _GEN_14127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14129 = 10'h1dc == _T_33 ? ram_476 : _GEN_14128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14130 = 10'h1dd == _T_33 ? ram_477 : _GEN_14129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14131 = 10'h1de == _T_33 ? ram_478 : _GEN_14130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14132 = 10'h1df == _T_33 ? ram_479 : _GEN_14131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14133 = 10'h1e0 == _T_33 ? ram_480 : _GEN_14132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14134 = 10'h1e1 == _T_33 ? ram_481 : _GEN_14133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14135 = 10'h1e2 == _T_33 ? ram_482 : _GEN_14134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14136 = 10'h1e3 == _T_33 ? ram_483 : _GEN_14135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14137 = 10'h1e4 == _T_33 ? ram_484 : _GEN_14136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14138 = 10'h1e5 == _T_33 ? ram_485 : _GEN_14137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14139 = 10'h1e6 == _T_33 ? ram_486 : _GEN_14138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14140 = 10'h1e7 == _T_33 ? ram_487 : _GEN_14139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14141 = 10'h1e8 == _T_33 ? ram_488 : _GEN_14140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14142 = 10'h1e9 == _T_33 ? ram_489 : _GEN_14141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14143 = 10'h1ea == _T_33 ? ram_490 : _GEN_14142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14144 = 10'h1eb == _T_33 ? ram_491 : _GEN_14143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14145 = 10'h1ec == _T_33 ? ram_492 : _GEN_14144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14146 = 10'h1ed == _T_33 ? ram_493 : _GEN_14145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14147 = 10'h1ee == _T_33 ? ram_494 : _GEN_14146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14148 = 10'h1ef == _T_33 ? ram_495 : _GEN_14147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14149 = 10'h1f0 == _T_33 ? ram_496 : _GEN_14148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14150 = 10'h1f1 == _T_33 ? ram_497 : _GEN_14149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14151 = 10'h1f2 == _T_33 ? ram_498 : _GEN_14150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14152 = 10'h1f3 == _T_33 ? ram_499 : _GEN_14151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14153 = 10'h1f4 == _T_33 ? ram_500 : _GEN_14152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14154 = 10'h1f5 == _T_33 ? ram_501 : _GEN_14153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14155 = 10'h1f6 == _T_33 ? ram_502 : _GEN_14154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14156 = 10'h1f7 == _T_33 ? ram_503 : _GEN_14155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14157 = 10'h1f8 == _T_33 ? ram_504 : _GEN_14156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14158 = 10'h1f9 == _T_33 ? ram_505 : _GEN_14157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14159 = 10'h1fa == _T_33 ? ram_506 : _GEN_14158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14160 = 10'h1fb == _T_33 ? ram_507 : _GEN_14159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14161 = 10'h1fc == _T_33 ? ram_508 : _GEN_14160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14162 = 10'h1fd == _T_33 ? ram_509 : _GEN_14161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14163 = 10'h1fe == _T_33 ? ram_510 : _GEN_14162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14164 = 10'h1ff == _T_33 ? ram_511 : _GEN_14163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14165 = 10'h200 == _T_33 ? ram_512 : _GEN_14164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14166 = 10'h201 == _T_33 ? ram_513 : _GEN_14165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14167 = 10'h202 == _T_33 ? ram_514 : _GEN_14166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14168 = 10'h203 == _T_33 ? ram_515 : _GEN_14167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14169 = 10'h204 == _T_33 ? ram_516 : _GEN_14168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14170 = 10'h205 == _T_33 ? ram_517 : _GEN_14169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14171 = 10'h206 == _T_33 ? ram_518 : _GEN_14170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14172 = 10'h207 == _T_33 ? ram_519 : _GEN_14171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14173 = 10'h208 == _T_33 ? ram_520 : _GEN_14172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14174 = 10'h209 == _T_33 ? ram_521 : _GEN_14173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14175 = 10'h20a == _T_33 ? ram_522 : _GEN_14174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14176 = 10'h20b == _T_33 ? ram_523 : _GEN_14175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14177 = 10'h20c == _T_33 ? ram_524 : _GEN_14176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19087 = {{8190'd0}, _GEN_14177}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_363 = _GEN_19087 ^ _ram_T_362; // @[vga.scala 64:41]
  wire [287:0] _GEN_14178 = 10'h0 == _T_33 ? _ram_T_363[287:0] : _GEN_13128; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14179 = 10'h1 == _T_33 ? _ram_T_363[287:0] : _GEN_13129; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14180 = 10'h2 == _T_33 ? _ram_T_363[287:0] : _GEN_13130; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14181 = 10'h3 == _T_33 ? _ram_T_363[287:0] : _GEN_13131; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14182 = 10'h4 == _T_33 ? _ram_T_363[287:0] : _GEN_13132; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14183 = 10'h5 == _T_33 ? _ram_T_363[287:0] : _GEN_13133; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14184 = 10'h6 == _T_33 ? _ram_T_363[287:0] : _GEN_13134; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14185 = 10'h7 == _T_33 ? _ram_T_363[287:0] : _GEN_13135; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14186 = 10'h8 == _T_33 ? _ram_T_363[287:0] : _GEN_13136; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14187 = 10'h9 == _T_33 ? _ram_T_363[287:0] : _GEN_13137; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14188 = 10'ha == _T_33 ? _ram_T_363[287:0] : _GEN_13138; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14189 = 10'hb == _T_33 ? _ram_T_363[287:0] : _GEN_13139; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14190 = 10'hc == _T_33 ? _ram_T_363[287:0] : _GEN_13140; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14191 = 10'hd == _T_33 ? _ram_T_363[287:0] : _GEN_13141; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14192 = 10'he == _T_33 ? _ram_T_363[287:0] : _GEN_13142; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14193 = 10'hf == _T_33 ? _ram_T_363[287:0] : _GEN_13143; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14194 = 10'h10 == _T_33 ? _ram_T_363[287:0] : _GEN_13144; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14195 = 10'h11 == _T_33 ? _ram_T_363[287:0] : _GEN_13145; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14196 = 10'h12 == _T_33 ? _ram_T_363[287:0] : _GEN_13146; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14197 = 10'h13 == _T_33 ? _ram_T_363[287:0] : _GEN_13147; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14198 = 10'h14 == _T_33 ? _ram_T_363[287:0] : _GEN_13148; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14199 = 10'h15 == _T_33 ? _ram_T_363[287:0] : _GEN_13149; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14200 = 10'h16 == _T_33 ? _ram_T_363[287:0] : _GEN_13150; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14201 = 10'h17 == _T_33 ? _ram_T_363[287:0] : _GEN_13151; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14202 = 10'h18 == _T_33 ? _ram_T_363[287:0] : _GEN_13152; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14203 = 10'h19 == _T_33 ? _ram_T_363[287:0] : _GEN_13153; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14204 = 10'h1a == _T_33 ? _ram_T_363[287:0] : _GEN_13154; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14205 = 10'h1b == _T_33 ? _ram_T_363[287:0] : _GEN_13155; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14206 = 10'h1c == _T_33 ? _ram_T_363[287:0] : _GEN_13156; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14207 = 10'h1d == _T_33 ? _ram_T_363[287:0] : _GEN_13157; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14208 = 10'h1e == _T_33 ? _ram_T_363[287:0] : _GEN_13158; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14209 = 10'h1f == _T_33 ? _ram_T_363[287:0] : _GEN_13159; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14210 = 10'h20 == _T_33 ? _ram_T_363[287:0] : _GEN_13160; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14211 = 10'h21 == _T_33 ? _ram_T_363[287:0] : _GEN_13161; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14212 = 10'h22 == _T_33 ? _ram_T_363[287:0] : _GEN_13162; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14213 = 10'h23 == _T_33 ? _ram_T_363[287:0] : _GEN_13163; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14214 = 10'h24 == _T_33 ? _ram_T_363[287:0] : _GEN_13164; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14215 = 10'h25 == _T_33 ? _ram_T_363[287:0] : _GEN_13165; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14216 = 10'h26 == _T_33 ? _ram_T_363[287:0] : _GEN_13166; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14217 = 10'h27 == _T_33 ? _ram_T_363[287:0] : _GEN_13167; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14218 = 10'h28 == _T_33 ? _ram_T_363[287:0] : _GEN_13168; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14219 = 10'h29 == _T_33 ? _ram_T_363[287:0] : _GEN_13169; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14220 = 10'h2a == _T_33 ? _ram_T_363[287:0] : _GEN_13170; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14221 = 10'h2b == _T_33 ? _ram_T_363[287:0] : _GEN_13171; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14222 = 10'h2c == _T_33 ? _ram_T_363[287:0] : _GEN_13172; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14223 = 10'h2d == _T_33 ? _ram_T_363[287:0] : _GEN_13173; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14224 = 10'h2e == _T_33 ? _ram_T_363[287:0] : _GEN_13174; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14225 = 10'h2f == _T_33 ? _ram_T_363[287:0] : _GEN_13175; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14226 = 10'h30 == _T_33 ? _ram_T_363[287:0] : _GEN_13176; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14227 = 10'h31 == _T_33 ? _ram_T_363[287:0] : _GEN_13177; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14228 = 10'h32 == _T_33 ? _ram_T_363[287:0] : _GEN_13178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14229 = 10'h33 == _T_33 ? _ram_T_363[287:0] : _GEN_13179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14230 = 10'h34 == _T_33 ? _ram_T_363[287:0] : _GEN_13180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14231 = 10'h35 == _T_33 ? _ram_T_363[287:0] : _GEN_13181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14232 = 10'h36 == _T_33 ? _ram_T_363[287:0] : _GEN_13182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14233 = 10'h37 == _T_33 ? _ram_T_363[287:0] : _GEN_13183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14234 = 10'h38 == _T_33 ? _ram_T_363[287:0] : _GEN_13184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14235 = 10'h39 == _T_33 ? _ram_T_363[287:0] : _GEN_13185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14236 = 10'h3a == _T_33 ? _ram_T_363[287:0] : _GEN_13186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14237 = 10'h3b == _T_33 ? _ram_T_363[287:0] : _GEN_13187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14238 = 10'h3c == _T_33 ? _ram_T_363[287:0] : _GEN_13188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14239 = 10'h3d == _T_33 ? _ram_T_363[287:0] : _GEN_13189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14240 = 10'h3e == _T_33 ? _ram_T_363[287:0] : _GEN_13190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14241 = 10'h3f == _T_33 ? _ram_T_363[287:0] : _GEN_13191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14242 = 10'h40 == _T_33 ? _ram_T_363[287:0] : _GEN_13192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14243 = 10'h41 == _T_33 ? _ram_T_363[287:0] : _GEN_13193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14244 = 10'h42 == _T_33 ? _ram_T_363[287:0] : _GEN_13194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14245 = 10'h43 == _T_33 ? _ram_T_363[287:0] : _GEN_13195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14246 = 10'h44 == _T_33 ? _ram_T_363[287:0] : _GEN_13196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14247 = 10'h45 == _T_33 ? _ram_T_363[287:0] : _GEN_13197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14248 = 10'h46 == _T_33 ? _ram_T_363[287:0] : _GEN_13198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14249 = 10'h47 == _T_33 ? _ram_T_363[287:0] : _GEN_13199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14250 = 10'h48 == _T_33 ? _ram_T_363[287:0] : _GEN_13200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14251 = 10'h49 == _T_33 ? _ram_T_363[287:0] : _GEN_13201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14252 = 10'h4a == _T_33 ? _ram_T_363[287:0] : _GEN_13202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14253 = 10'h4b == _T_33 ? _ram_T_363[287:0] : _GEN_13203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14254 = 10'h4c == _T_33 ? _ram_T_363[287:0] : _GEN_13204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14255 = 10'h4d == _T_33 ? _ram_T_363[287:0] : _GEN_13205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14256 = 10'h4e == _T_33 ? _ram_T_363[287:0] : _GEN_13206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14257 = 10'h4f == _T_33 ? _ram_T_363[287:0] : _GEN_13207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14258 = 10'h50 == _T_33 ? _ram_T_363[287:0] : _GEN_13208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14259 = 10'h51 == _T_33 ? _ram_T_363[287:0] : _GEN_13209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14260 = 10'h52 == _T_33 ? _ram_T_363[287:0] : _GEN_13210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14261 = 10'h53 == _T_33 ? _ram_T_363[287:0] : _GEN_13211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14262 = 10'h54 == _T_33 ? _ram_T_363[287:0] : _GEN_13212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14263 = 10'h55 == _T_33 ? _ram_T_363[287:0] : _GEN_13213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14264 = 10'h56 == _T_33 ? _ram_T_363[287:0] : _GEN_13214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14265 = 10'h57 == _T_33 ? _ram_T_363[287:0] : _GEN_13215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14266 = 10'h58 == _T_33 ? _ram_T_363[287:0] : _GEN_13216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14267 = 10'h59 == _T_33 ? _ram_T_363[287:0] : _GEN_13217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14268 = 10'h5a == _T_33 ? _ram_T_363[287:0] : _GEN_13218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14269 = 10'h5b == _T_33 ? _ram_T_363[287:0] : _GEN_13219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14270 = 10'h5c == _T_33 ? _ram_T_363[287:0] : _GEN_13220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14271 = 10'h5d == _T_33 ? _ram_T_363[287:0] : _GEN_13221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14272 = 10'h5e == _T_33 ? _ram_T_363[287:0] : _GEN_13222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14273 = 10'h5f == _T_33 ? _ram_T_363[287:0] : _GEN_13223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14274 = 10'h60 == _T_33 ? _ram_T_363[287:0] : _GEN_13224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14275 = 10'h61 == _T_33 ? _ram_T_363[287:0] : _GEN_13225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14276 = 10'h62 == _T_33 ? _ram_T_363[287:0] : _GEN_13226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14277 = 10'h63 == _T_33 ? _ram_T_363[287:0] : _GEN_13227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14278 = 10'h64 == _T_33 ? _ram_T_363[287:0] : _GEN_13228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14279 = 10'h65 == _T_33 ? _ram_T_363[287:0] : _GEN_13229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14280 = 10'h66 == _T_33 ? _ram_T_363[287:0] : _GEN_13230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14281 = 10'h67 == _T_33 ? _ram_T_363[287:0] : _GEN_13231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14282 = 10'h68 == _T_33 ? _ram_T_363[287:0] : _GEN_13232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14283 = 10'h69 == _T_33 ? _ram_T_363[287:0] : _GEN_13233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14284 = 10'h6a == _T_33 ? _ram_T_363[287:0] : _GEN_13234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14285 = 10'h6b == _T_33 ? _ram_T_363[287:0] : _GEN_13235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14286 = 10'h6c == _T_33 ? _ram_T_363[287:0] : _GEN_13236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14287 = 10'h6d == _T_33 ? _ram_T_363[287:0] : _GEN_13237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14288 = 10'h6e == _T_33 ? _ram_T_363[287:0] : _GEN_13238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14289 = 10'h6f == _T_33 ? _ram_T_363[287:0] : _GEN_13239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14290 = 10'h70 == _T_33 ? _ram_T_363[287:0] : _GEN_13240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14291 = 10'h71 == _T_33 ? _ram_T_363[287:0] : _GEN_13241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14292 = 10'h72 == _T_33 ? _ram_T_363[287:0] : _GEN_13242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14293 = 10'h73 == _T_33 ? _ram_T_363[287:0] : _GEN_13243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14294 = 10'h74 == _T_33 ? _ram_T_363[287:0] : _GEN_13244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14295 = 10'h75 == _T_33 ? _ram_T_363[287:0] : _GEN_13245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14296 = 10'h76 == _T_33 ? _ram_T_363[287:0] : _GEN_13246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14297 = 10'h77 == _T_33 ? _ram_T_363[287:0] : _GEN_13247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14298 = 10'h78 == _T_33 ? _ram_T_363[287:0] : _GEN_13248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14299 = 10'h79 == _T_33 ? _ram_T_363[287:0] : _GEN_13249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14300 = 10'h7a == _T_33 ? _ram_T_363[287:0] : _GEN_13250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14301 = 10'h7b == _T_33 ? _ram_T_363[287:0] : _GEN_13251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14302 = 10'h7c == _T_33 ? _ram_T_363[287:0] : _GEN_13252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14303 = 10'h7d == _T_33 ? _ram_T_363[287:0] : _GEN_13253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14304 = 10'h7e == _T_33 ? _ram_T_363[287:0] : _GEN_13254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14305 = 10'h7f == _T_33 ? _ram_T_363[287:0] : _GEN_13255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14306 = 10'h80 == _T_33 ? _ram_T_363[287:0] : _GEN_13256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14307 = 10'h81 == _T_33 ? _ram_T_363[287:0] : _GEN_13257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14308 = 10'h82 == _T_33 ? _ram_T_363[287:0] : _GEN_13258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14309 = 10'h83 == _T_33 ? _ram_T_363[287:0] : _GEN_13259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14310 = 10'h84 == _T_33 ? _ram_T_363[287:0] : _GEN_13260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14311 = 10'h85 == _T_33 ? _ram_T_363[287:0] : _GEN_13261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14312 = 10'h86 == _T_33 ? _ram_T_363[287:0] : _GEN_13262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14313 = 10'h87 == _T_33 ? _ram_T_363[287:0] : _GEN_13263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14314 = 10'h88 == _T_33 ? _ram_T_363[287:0] : _GEN_13264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14315 = 10'h89 == _T_33 ? _ram_T_363[287:0] : _GEN_13265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14316 = 10'h8a == _T_33 ? _ram_T_363[287:0] : _GEN_13266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14317 = 10'h8b == _T_33 ? _ram_T_363[287:0] : _GEN_13267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14318 = 10'h8c == _T_33 ? _ram_T_363[287:0] : _GEN_13268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14319 = 10'h8d == _T_33 ? _ram_T_363[287:0] : _GEN_13269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14320 = 10'h8e == _T_33 ? _ram_T_363[287:0] : _GEN_13270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14321 = 10'h8f == _T_33 ? _ram_T_363[287:0] : _GEN_13271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14322 = 10'h90 == _T_33 ? _ram_T_363[287:0] : _GEN_13272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14323 = 10'h91 == _T_33 ? _ram_T_363[287:0] : _GEN_13273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14324 = 10'h92 == _T_33 ? _ram_T_363[287:0] : _GEN_13274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14325 = 10'h93 == _T_33 ? _ram_T_363[287:0] : _GEN_13275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14326 = 10'h94 == _T_33 ? _ram_T_363[287:0] : _GEN_13276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14327 = 10'h95 == _T_33 ? _ram_T_363[287:0] : _GEN_13277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14328 = 10'h96 == _T_33 ? _ram_T_363[287:0] : _GEN_13278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14329 = 10'h97 == _T_33 ? _ram_T_363[287:0] : _GEN_13279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14330 = 10'h98 == _T_33 ? _ram_T_363[287:0] : _GEN_13280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14331 = 10'h99 == _T_33 ? _ram_T_363[287:0] : _GEN_13281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14332 = 10'h9a == _T_33 ? _ram_T_363[287:0] : _GEN_13282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14333 = 10'h9b == _T_33 ? _ram_T_363[287:0] : _GEN_13283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14334 = 10'h9c == _T_33 ? _ram_T_363[287:0] : _GEN_13284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14335 = 10'h9d == _T_33 ? _ram_T_363[287:0] : _GEN_13285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14336 = 10'h9e == _T_33 ? _ram_T_363[287:0] : _GEN_13286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14337 = 10'h9f == _T_33 ? _ram_T_363[287:0] : _GEN_13287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14338 = 10'ha0 == _T_33 ? _ram_T_363[287:0] : _GEN_13288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14339 = 10'ha1 == _T_33 ? _ram_T_363[287:0] : _GEN_13289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14340 = 10'ha2 == _T_33 ? _ram_T_363[287:0] : _GEN_13290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14341 = 10'ha3 == _T_33 ? _ram_T_363[287:0] : _GEN_13291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14342 = 10'ha4 == _T_33 ? _ram_T_363[287:0] : _GEN_13292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14343 = 10'ha5 == _T_33 ? _ram_T_363[287:0] : _GEN_13293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14344 = 10'ha6 == _T_33 ? _ram_T_363[287:0] : _GEN_13294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14345 = 10'ha7 == _T_33 ? _ram_T_363[287:0] : _GEN_13295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14346 = 10'ha8 == _T_33 ? _ram_T_363[287:0] : _GEN_13296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14347 = 10'ha9 == _T_33 ? _ram_T_363[287:0] : _GEN_13297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14348 = 10'haa == _T_33 ? _ram_T_363[287:0] : _GEN_13298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14349 = 10'hab == _T_33 ? _ram_T_363[287:0] : _GEN_13299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14350 = 10'hac == _T_33 ? _ram_T_363[287:0] : _GEN_13300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14351 = 10'had == _T_33 ? _ram_T_363[287:0] : _GEN_13301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14352 = 10'hae == _T_33 ? _ram_T_363[287:0] : _GEN_13302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14353 = 10'haf == _T_33 ? _ram_T_363[287:0] : _GEN_13303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14354 = 10'hb0 == _T_33 ? _ram_T_363[287:0] : _GEN_13304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14355 = 10'hb1 == _T_33 ? _ram_T_363[287:0] : _GEN_13305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14356 = 10'hb2 == _T_33 ? _ram_T_363[287:0] : _GEN_13306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14357 = 10'hb3 == _T_33 ? _ram_T_363[287:0] : _GEN_13307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14358 = 10'hb4 == _T_33 ? _ram_T_363[287:0] : _GEN_13308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14359 = 10'hb5 == _T_33 ? _ram_T_363[287:0] : _GEN_13309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14360 = 10'hb6 == _T_33 ? _ram_T_363[287:0] : _GEN_13310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14361 = 10'hb7 == _T_33 ? _ram_T_363[287:0] : _GEN_13311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14362 = 10'hb8 == _T_33 ? _ram_T_363[287:0] : _GEN_13312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14363 = 10'hb9 == _T_33 ? _ram_T_363[287:0] : _GEN_13313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14364 = 10'hba == _T_33 ? _ram_T_363[287:0] : _GEN_13314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14365 = 10'hbb == _T_33 ? _ram_T_363[287:0] : _GEN_13315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14366 = 10'hbc == _T_33 ? _ram_T_363[287:0] : _GEN_13316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14367 = 10'hbd == _T_33 ? _ram_T_363[287:0] : _GEN_13317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14368 = 10'hbe == _T_33 ? _ram_T_363[287:0] : _GEN_13318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14369 = 10'hbf == _T_33 ? _ram_T_363[287:0] : _GEN_13319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14370 = 10'hc0 == _T_33 ? _ram_T_363[287:0] : _GEN_13320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14371 = 10'hc1 == _T_33 ? _ram_T_363[287:0] : _GEN_13321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14372 = 10'hc2 == _T_33 ? _ram_T_363[287:0] : _GEN_13322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14373 = 10'hc3 == _T_33 ? _ram_T_363[287:0] : _GEN_13323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14374 = 10'hc4 == _T_33 ? _ram_T_363[287:0] : _GEN_13324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14375 = 10'hc5 == _T_33 ? _ram_T_363[287:0] : _GEN_13325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14376 = 10'hc6 == _T_33 ? _ram_T_363[287:0] : _GEN_13326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14377 = 10'hc7 == _T_33 ? _ram_T_363[287:0] : _GEN_13327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14378 = 10'hc8 == _T_33 ? _ram_T_363[287:0] : _GEN_13328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14379 = 10'hc9 == _T_33 ? _ram_T_363[287:0] : _GEN_13329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14380 = 10'hca == _T_33 ? _ram_T_363[287:0] : _GEN_13330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14381 = 10'hcb == _T_33 ? _ram_T_363[287:0] : _GEN_13331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14382 = 10'hcc == _T_33 ? _ram_T_363[287:0] : _GEN_13332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14383 = 10'hcd == _T_33 ? _ram_T_363[287:0] : _GEN_13333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14384 = 10'hce == _T_33 ? _ram_T_363[287:0] : _GEN_13334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14385 = 10'hcf == _T_33 ? _ram_T_363[287:0] : _GEN_13335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14386 = 10'hd0 == _T_33 ? _ram_T_363[287:0] : _GEN_13336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14387 = 10'hd1 == _T_33 ? _ram_T_363[287:0] : _GEN_13337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14388 = 10'hd2 == _T_33 ? _ram_T_363[287:0] : _GEN_13338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14389 = 10'hd3 == _T_33 ? _ram_T_363[287:0] : _GEN_13339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14390 = 10'hd4 == _T_33 ? _ram_T_363[287:0] : _GEN_13340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14391 = 10'hd5 == _T_33 ? _ram_T_363[287:0] : _GEN_13341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14392 = 10'hd6 == _T_33 ? _ram_T_363[287:0] : _GEN_13342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14393 = 10'hd7 == _T_33 ? _ram_T_363[287:0] : _GEN_13343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14394 = 10'hd8 == _T_33 ? _ram_T_363[287:0] : _GEN_13344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14395 = 10'hd9 == _T_33 ? _ram_T_363[287:0] : _GEN_13345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14396 = 10'hda == _T_33 ? _ram_T_363[287:0] : _GEN_13346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14397 = 10'hdb == _T_33 ? _ram_T_363[287:0] : _GEN_13347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14398 = 10'hdc == _T_33 ? _ram_T_363[287:0] : _GEN_13348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14399 = 10'hdd == _T_33 ? _ram_T_363[287:0] : _GEN_13349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14400 = 10'hde == _T_33 ? _ram_T_363[287:0] : _GEN_13350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14401 = 10'hdf == _T_33 ? _ram_T_363[287:0] : _GEN_13351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14402 = 10'he0 == _T_33 ? _ram_T_363[287:0] : _GEN_13352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14403 = 10'he1 == _T_33 ? _ram_T_363[287:0] : _GEN_13353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14404 = 10'he2 == _T_33 ? _ram_T_363[287:0] : _GEN_13354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14405 = 10'he3 == _T_33 ? _ram_T_363[287:0] : _GEN_13355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14406 = 10'he4 == _T_33 ? _ram_T_363[287:0] : _GEN_13356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14407 = 10'he5 == _T_33 ? _ram_T_363[287:0] : _GEN_13357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14408 = 10'he6 == _T_33 ? _ram_T_363[287:0] : _GEN_13358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14409 = 10'he7 == _T_33 ? _ram_T_363[287:0] : _GEN_13359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14410 = 10'he8 == _T_33 ? _ram_T_363[287:0] : _GEN_13360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14411 = 10'he9 == _T_33 ? _ram_T_363[287:0] : _GEN_13361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14412 = 10'hea == _T_33 ? _ram_T_363[287:0] : _GEN_13362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14413 = 10'heb == _T_33 ? _ram_T_363[287:0] : _GEN_13363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14414 = 10'hec == _T_33 ? _ram_T_363[287:0] : _GEN_13364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14415 = 10'hed == _T_33 ? _ram_T_363[287:0] : _GEN_13365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14416 = 10'hee == _T_33 ? _ram_T_363[287:0] : _GEN_13366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14417 = 10'hef == _T_33 ? _ram_T_363[287:0] : _GEN_13367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14418 = 10'hf0 == _T_33 ? _ram_T_363[287:0] : _GEN_13368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14419 = 10'hf1 == _T_33 ? _ram_T_363[287:0] : _GEN_13369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14420 = 10'hf2 == _T_33 ? _ram_T_363[287:0] : _GEN_13370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14421 = 10'hf3 == _T_33 ? _ram_T_363[287:0] : _GEN_13371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14422 = 10'hf4 == _T_33 ? _ram_T_363[287:0] : _GEN_13372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14423 = 10'hf5 == _T_33 ? _ram_T_363[287:0] : _GEN_13373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14424 = 10'hf6 == _T_33 ? _ram_T_363[287:0] : _GEN_13374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14425 = 10'hf7 == _T_33 ? _ram_T_363[287:0] : _GEN_13375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14426 = 10'hf8 == _T_33 ? _ram_T_363[287:0] : _GEN_13376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14427 = 10'hf9 == _T_33 ? _ram_T_363[287:0] : _GEN_13377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14428 = 10'hfa == _T_33 ? _ram_T_363[287:0] : _GEN_13378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14429 = 10'hfb == _T_33 ? _ram_T_363[287:0] : _GEN_13379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14430 = 10'hfc == _T_33 ? _ram_T_363[287:0] : _GEN_13380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14431 = 10'hfd == _T_33 ? _ram_T_363[287:0] : _GEN_13381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14432 = 10'hfe == _T_33 ? _ram_T_363[287:0] : _GEN_13382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14433 = 10'hff == _T_33 ? _ram_T_363[287:0] : _GEN_13383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14434 = 10'h100 == _T_33 ? _ram_T_363[287:0] : _GEN_13384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14435 = 10'h101 == _T_33 ? _ram_T_363[287:0] : _GEN_13385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14436 = 10'h102 == _T_33 ? _ram_T_363[287:0] : _GEN_13386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14437 = 10'h103 == _T_33 ? _ram_T_363[287:0] : _GEN_13387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14438 = 10'h104 == _T_33 ? _ram_T_363[287:0] : _GEN_13388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14439 = 10'h105 == _T_33 ? _ram_T_363[287:0] : _GEN_13389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14440 = 10'h106 == _T_33 ? _ram_T_363[287:0] : _GEN_13390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14441 = 10'h107 == _T_33 ? _ram_T_363[287:0] : _GEN_13391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14442 = 10'h108 == _T_33 ? _ram_T_363[287:0] : _GEN_13392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14443 = 10'h109 == _T_33 ? _ram_T_363[287:0] : _GEN_13393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14444 = 10'h10a == _T_33 ? _ram_T_363[287:0] : _GEN_13394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14445 = 10'h10b == _T_33 ? _ram_T_363[287:0] : _GEN_13395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14446 = 10'h10c == _T_33 ? _ram_T_363[287:0] : _GEN_13396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14447 = 10'h10d == _T_33 ? _ram_T_363[287:0] : _GEN_13397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14448 = 10'h10e == _T_33 ? _ram_T_363[287:0] : _GEN_13398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14449 = 10'h10f == _T_33 ? _ram_T_363[287:0] : _GEN_13399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14450 = 10'h110 == _T_33 ? _ram_T_363[287:0] : _GEN_13400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14451 = 10'h111 == _T_33 ? _ram_T_363[287:0] : _GEN_13401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14452 = 10'h112 == _T_33 ? _ram_T_363[287:0] : _GEN_13402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14453 = 10'h113 == _T_33 ? _ram_T_363[287:0] : _GEN_13403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14454 = 10'h114 == _T_33 ? _ram_T_363[287:0] : _GEN_13404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14455 = 10'h115 == _T_33 ? _ram_T_363[287:0] : _GEN_13405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14456 = 10'h116 == _T_33 ? _ram_T_363[287:0] : _GEN_13406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14457 = 10'h117 == _T_33 ? _ram_T_363[287:0] : _GEN_13407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14458 = 10'h118 == _T_33 ? _ram_T_363[287:0] : _GEN_13408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14459 = 10'h119 == _T_33 ? _ram_T_363[287:0] : _GEN_13409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14460 = 10'h11a == _T_33 ? _ram_T_363[287:0] : _GEN_13410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14461 = 10'h11b == _T_33 ? _ram_T_363[287:0] : _GEN_13411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14462 = 10'h11c == _T_33 ? _ram_T_363[287:0] : _GEN_13412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14463 = 10'h11d == _T_33 ? _ram_T_363[287:0] : _GEN_13413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14464 = 10'h11e == _T_33 ? _ram_T_363[287:0] : _GEN_13414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14465 = 10'h11f == _T_33 ? _ram_T_363[287:0] : _GEN_13415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14466 = 10'h120 == _T_33 ? _ram_T_363[287:0] : _GEN_13416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14467 = 10'h121 == _T_33 ? _ram_T_363[287:0] : _GEN_13417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14468 = 10'h122 == _T_33 ? _ram_T_363[287:0] : _GEN_13418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14469 = 10'h123 == _T_33 ? _ram_T_363[287:0] : _GEN_13419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14470 = 10'h124 == _T_33 ? _ram_T_363[287:0] : _GEN_13420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14471 = 10'h125 == _T_33 ? _ram_T_363[287:0] : _GEN_13421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14472 = 10'h126 == _T_33 ? _ram_T_363[287:0] : _GEN_13422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14473 = 10'h127 == _T_33 ? _ram_T_363[287:0] : _GEN_13423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14474 = 10'h128 == _T_33 ? _ram_T_363[287:0] : _GEN_13424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14475 = 10'h129 == _T_33 ? _ram_T_363[287:0] : _GEN_13425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14476 = 10'h12a == _T_33 ? _ram_T_363[287:0] : _GEN_13426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14477 = 10'h12b == _T_33 ? _ram_T_363[287:0] : _GEN_13427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14478 = 10'h12c == _T_33 ? _ram_T_363[287:0] : _GEN_13428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14479 = 10'h12d == _T_33 ? _ram_T_363[287:0] : _GEN_13429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14480 = 10'h12e == _T_33 ? _ram_T_363[287:0] : _GEN_13430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14481 = 10'h12f == _T_33 ? _ram_T_363[287:0] : _GEN_13431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14482 = 10'h130 == _T_33 ? _ram_T_363[287:0] : _GEN_13432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14483 = 10'h131 == _T_33 ? _ram_T_363[287:0] : _GEN_13433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14484 = 10'h132 == _T_33 ? _ram_T_363[287:0] : _GEN_13434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14485 = 10'h133 == _T_33 ? _ram_T_363[287:0] : _GEN_13435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14486 = 10'h134 == _T_33 ? _ram_T_363[287:0] : _GEN_13436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14487 = 10'h135 == _T_33 ? _ram_T_363[287:0] : _GEN_13437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14488 = 10'h136 == _T_33 ? _ram_T_363[287:0] : _GEN_13438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14489 = 10'h137 == _T_33 ? _ram_T_363[287:0] : _GEN_13439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14490 = 10'h138 == _T_33 ? _ram_T_363[287:0] : _GEN_13440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14491 = 10'h139 == _T_33 ? _ram_T_363[287:0] : _GEN_13441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14492 = 10'h13a == _T_33 ? _ram_T_363[287:0] : _GEN_13442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14493 = 10'h13b == _T_33 ? _ram_T_363[287:0] : _GEN_13443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14494 = 10'h13c == _T_33 ? _ram_T_363[287:0] : _GEN_13444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14495 = 10'h13d == _T_33 ? _ram_T_363[287:0] : _GEN_13445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14496 = 10'h13e == _T_33 ? _ram_T_363[287:0] : _GEN_13446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14497 = 10'h13f == _T_33 ? _ram_T_363[287:0] : _GEN_13447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14498 = 10'h140 == _T_33 ? _ram_T_363[287:0] : _GEN_13448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14499 = 10'h141 == _T_33 ? _ram_T_363[287:0] : _GEN_13449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14500 = 10'h142 == _T_33 ? _ram_T_363[287:0] : _GEN_13450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14501 = 10'h143 == _T_33 ? _ram_T_363[287:0] : _GEN_13451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14502 = 10'h144 == _T_33 ? _ram_T_363[287:0] : _GEN_13452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14503 = 10'h145 == _T_33 ? _ram_T_363[287:0] : _GEN_13453; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14504 = 10'h146 == _T_33 ? _ram_T_363[287:0] : _GEN_13454; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14505 = 10'h147 == _T_33 ? _ram_T_363[287:0] : _GEN_13455; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14506 = 10'h148 == _T_33 ? _ram_T_363[287:0] : _GEN_13456; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14507 = 10'h149 == _T_33 ? _ram_T_363[287:0] : _GEN_13457; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14508 = 10'h14a == _T_33 ? _ram_T_363[287:0] : _GEN_13458; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14509 = 10'h14b == _T_33 ? _ram_T_363[287:0] : _GEN_13459; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14510 = 10'h14c == _T_33 ? _ram_T_363[287:0] : _GEN_13460; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14511 = 10'h14d == _T_33 ? _ram_T_363[287:0] : _GEN_13461; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14512 = 10'h14e == _T_33 ? _ram_T_363[287:0] : _GEN_13462; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14513 = 10'h14f == _T_33 ? _ram_T_363[287:0] : _GEN_13463; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14514 = 10'h150 == _T_33 ? _ram_T_363[287:0] : _GEN_13464; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14515 = 10'h151 == _T_33 ? _ram_T_363[287:0] : _GEN_13465; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14516 = 10'h152 == _T_33 ? _ram_T_363[287:0] : _GEN_13466; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14517 = 10'h153 == _T_33 ? _ram_T_363[287:0] : _GEN_13467; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14518 = 10'h154 == _T_33 ? _ram_T_363[287:0] : _GEN_13468; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14519 = 10'h155 == _T_33 ? _ram_T_363[287:0] : _GEN_13469; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14520 = 10'h156 == _T_33 ? _ram_T_363[287:0] : _GEN_13470; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14521 = 10'h157 == _T_33 ? _ram_T_363[287:0] : _GEN_13471; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14522 = 10'h158 == _T_33 ? _ram_T_363[287:0] : _GEN_13472; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14523 = 10'h159 == _T_33 ? _ram_T_363[287:0] : _GEN_13473; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14524 = 10'h15a == _T_33 ? _ram_T_363[287:0] : _GEN_13474; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14525 = 10'h15b == _T_33 ? _ram_T_363[287:0] : _GEN_13475; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14526 = 10'h15c == _T_33 ? _ram_T_363[287:0] : _GEN_13476; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14527 = 10'h15d == _T_33 ? _ram_T_363[287:0] : _GEN_13477; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14528 = 10'h15e == _T_33 ? _ram_T_363[287:0] : _GEN_13478; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14529 = 10'h15f == _T_33 ? _ram_T_363[287:0] : _GEN_13479; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14530 = 10'h160 == _T_33 ? _ram_T_363[287:0] : _GEN_13480; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14531 = 10'h161 == _T_33 ? _ram_T_363[287:0] : _GEN_13481; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14532 = 10'h162 == _T_33 ? _ram_T_363[287:0] : _GEN_13482; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14533 = 10'h163 == _T_33 ? _ram_T_363[287:0] : _GEN_13483; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14534 = 10'h164 == _T_33 ? _ram_T_363[287:0] : _GEN_13484; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14535 = 10'h165 == _T_33 ? _ram_T_363[287:0] : _GEN_13485; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14536 = 10'h166 == _T_33 ? _ram_T_363[287:0] : _GEN_13486; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14537 = 10'h167 == _T_33 ? _ram_T_363[287:0] : _GEN_13487; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14538 = 10'h168 == _T_33 ? _ram_T_363[287:0] : _GEN_13488; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14539 = 10'h169 == _T_33 ? _ram_T_363[287:0] : _GEN_13489; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14540 = 10'h16a == _T_33 ? _ram_T_363[287:0] : _GEN_13490; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14541 = 10'h16b == _T_33 ? _ram_T_363[287:0] : _GEN_13491; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14542 = 10'h16c == _T_33 ? _ram_T_363[287:0] : _GEN_13492; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14543 = 10'h16d == _T_33 ? _ram_T_363[287:0] : _GEN_13493; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14544 = 10'h16e == _T_33 ? _ram_T_363[287:0] : _GEN_13494; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14545 = 10'h16f == _T_33 ? _ram_T_363[287:0] : _GEN_13495; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14546 = 10'h170 == _T_33 ? _ram_T_363[287:0] : _GEN_13496; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14547 = 10'h171 == _T_33 ? _ram_T_363[287:0] : _GEN_13497; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14548 = 10'h172 == _T_33 ? _ram_T_363[287:0] : _GEN_13498; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14549 = 10'h173 == _T_33 ? _ram_T_363[287:0] : _GEN_13499; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14550 = 10'h174 == _T_33 ? _ram_T_363[287:0] : _GEN_13500; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14551 = 10'h175 == _T_33 ? _ram_T_363[287:0] : _GEN_13501; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14552 = 10'h176 == _T_33 ? _ram_T_363[287:0] : _GEN_13502; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14553 = 10'h177 == _T_33 ? _ram_T_363[287:0] : _GEN_13503; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14554 = 10'h178 == _T_33 ? _ram_T_363[287:0] : _GEN_13504; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14555 = 10'h179 == _T_33 ? _ram_T_363[287:0] : _GEN_13505; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14556 = 10'h17a == _T_33 ? _ram_T_363[287:0] : _GEN_13506; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14557 = 10'h17b == _T_33 ? _ram_T_363[287:0] : _GEN_13507; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14558 = 10'h17c == _T_33 ? _ram_T_363[287:0] : _GEN_13508; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14559 = 10'h17d == _T_33 ? _ram_T_363[287:0] : _GEN_13509; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14560 = 10'h17e == _T_33 ? _ram_T_363[287:0] : _GEN_13510; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14561 = 10'h17f == _T_33 ? _ram_T_363[287:0] : _GEN_13511; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14562 = 10'h180 == _T_33 ? _ram_T_363[287:0] : _GEN_13512; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14563 = 10'h181 == _T_33 ? _ram_T_363[287:0] : _GEN_13513; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14564 = 10'h182 == _T_33 ? _ram_T_363[287:0] : _GEN_13514; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14565 = 10'h183 == _T_33 ? _ram_T_363[287:0] : _GEN_13515; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14566 = 10'h184 == _T_33 ? _ram_T_363[287:0] : _GEN_13516; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14567 = 10'h185 == _T_33 ? _ram_T_363[287:0] : _GEN_13517; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14568 = 10'h186 == _T_33 ? _ram_T_363[287:0] : _GEN_13518; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14569 = 10'h187 == _T_33 ? _ram_T_363[287:0] : _GEN_13519; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14570 = 10'h188 == _T_33 ? _ram_T_363[287:0] : _GEN_13520; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14571 = 10'h189 == _T_33 ? _ram_T_363[287:0] : _GEN_13521; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14572 = 10'h18a == _T_33 ? _ram_T_363[287:0] : _GEN_13522; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14573 = 10'h18b == _T_33 ? _ram_T_363[287:0] : _GEN_13523; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14574 = 10'h18c == _T_33 ? _ram_T_363[287:0] : _GEN_13524; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14575 = 10'h18d == _T_33 ? _ram_T_363[287:0] : _GEN_13525; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14576 = 10'h18e == _T_33 ? _ram_T_363[287:0] : _GEN_13526; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14577 = 10'h18f == _T_33 ? _ram_T_363[287:0] : _GEN_13527; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14578 = 10'h190 == _T_33 ? _ram_T_363[287:0] : _GEN_13528; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14579 = 10'h191 == _T_33 ? _ram_T_363[287:0] : _GEN_13529; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14580 = 10'h192 == _T_33 ? _ram_T_363[287:0] : _GEN_13530; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14581 = 10'h193 == _T_33 ? _ram_T_363[287:0] : _GEN_13531; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14582 = 10'h194 == _T_33 ? _ram_T_363[287:0] : _GEN_13532; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14583 = 10'h195 == _T_33 ? _ram_T_363[287:0] : _GEN_13533; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14584 = 10'h196 == _T_33 ? _ram_T_363[287:0] : _GEN_13534; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14585 = 10'h197 == _T_33 ? _ram_T_363[287:0] : _GEN_13535; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14586 = 10'h198 == _T_33 ? _ram_T_363[287:0] : _GEN_13536; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14587 = 10'h199 == _T_33 ? _ram_T_363[287:0] : _GEN_13537; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14588 = 10'h19a == _T_33 ? _ram_T_363[287:0] : _GEN_13538; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14589 = 10'h19b == _T_33 ? _ram_T_363[287:0] : _GEN_13539; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14590 = 10'h19c == _T_33 ? _ram_T_363[287:0] : _GEN_13540; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14591 = 10'h19d == _T_33 ? _ram_T_363[287:0] : _GEN_13541; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14592 = 10'h19e == _T_33 ? _ram_T_363[287:0] : _GEN_13542; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14593 = 10'h19f == _T_33 ? _ram_T_363[287:0] : _GEN_13543; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14594 = 10'h1a0 == _T_33 ? _ram_T_363[287:0] : _GEN_13544; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14595 = 10'h1a1 == _T_33 ? _ram_T_363[287:0] : _GEN_13545; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14596 = 10'h1a2 == _T_33 ? _ram_T_363[287:0] : _GEN_13546; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14597 = 10'h1a3 == _T_33 ? _ram_T_363[287:0] : _GEN_13547; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14598 = 10'h1a4 == _T_33 ? _ram_T_363[287:0] : _GEN_13548; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14599 = 10'h1a5 == _T_33 ? _ram_T_363[287:0] : _GEN_13549; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14600 = 10'h1a6 == _T_33 ? _ram_T_363[287:0] : _GEN_13550; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14601 = 10'h1a7 == _T_33 ? _ram_T_363[287:0] : _GEN_13551; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14602 = 10'h1a8 == _T_33 ? _ram_T_363[287:0] : _GEN_13552; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14603 = 10'h1a9 == _T_33 ? _ram_T_363[287:0] : _GEN_13553; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14604 = 10'h1aa == _T_33 ? _ram_T_363[287:0] : _GEN_13554; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14605 = 10'h1ab == _T_33 ? _ram_T_363[287:0] : _GEN_13555; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14606 = 10'h1ac == _T_33 ? _ram_T_363[287:0] : _GEN_13556; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14607 = 10'h1ad == _T_33 ? _ram_T_363[287:0] : _GEN_13557; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14608 = 10'h1ae == _T_33 ? _ram_T_363[287:0] : _GEN_13558; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14609 = 10'h1af == _T_33 ? _ram_T_363[287:0] : _GEN_13559; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14610 = 10'h1b0 == _T_33 ? _ram_T_363[287:0] : _GEN_13560; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14611 = 10'h1b1 == _T_33 ? _ram_T_363[287:0] : _GEN_13561; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14612 = 10'h1b2 == _T_33 ? _ram_T_363[287:0] : _GEN_13562; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14613 = 10'h1b3 == _T_33 ? _ram_T_363[287:0] : _GEN_13563; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14614 = 10'h1b4 == _T_33 ? _ram_T_363[287:0] : _GEN_13564; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14615 = 10'h1b5 == _T_33 ? _ram_T_363[287:0] : _GEN_13565; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14616 = 10'h1b6 == _T_33 ? _ram_T_363[287:0] : _GEN_13566; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14617 = 10'h1b7 == _T_33 ? _ram_T_363[287:0] : _GEN_13567; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14618 = 10'h1b8 == _T_33 ? _ram_T_363[287:0] : _GEN_13568; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14619 = 10'h1b9 == _T_33 ? _ram_T_363[287:0] : _GEN_13569; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14620 = 10'h1ba == _T_33 ? _ram_T_363[287:0] : _GEN_13570; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14621 = 10'h1bb == _T_33 ? _ram_T_363[287:0] : _GEN_13571; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14622 = 10'h1bc == _T_33 ? _ram_T_363[287:0] : _GEN_13572; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14623 = 10'h1bd == _T_33 ? _ram_T_363[287:0] : _GEN_13573; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14624 = 10'h1be == _T_33 ? _ram_T_363[287:0] : _GEN_13574; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14625 = 10'h1bf == _T_33 ? _ram_T_363[287:0] : _GEN_13575; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14626 = 10'h1c0 == _T_33 ? _ram_T_363[287:0] : _GEN_13576; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14627 = 10'h1c1 == _T_33 ? _ram_T_363[287:0] : _GEN_13577; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14628 = 10'h1c2 == _T_33 ? _ram_T_363[287:0] : _GEN_13578; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14629 = 10'h1c3 == _T_33 ? _ram_T_363[287:0] : _GEN_13579; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14630 = 10'h1c4 == _T_33 ? _ram_T_363[287:0] : _GEN_13580; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14631 = 10'h1c5 == _T_33 ? _ram_T_363[287:0] : _GEN_13581; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14632 = 10'h1c6 == _T_33 ? _ram_T_363[287:0] : _GEN_13582; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14633 = 10'h1c7 == _T_33 ? _ram_T_363[287:0] : _GEN_13583; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14634 = 10'h1c8 == _T_33 ? _ram_T_363[287:0] : _GEN_13584; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14635 = 10'h1c9 == _T_33 ? _ram_T_363[287:0] : _GEN_13585; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14636 = 10'h1ca == _T_33 ? _ram_T_363[287:0] : _GEN_13586; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14637 = 10'h1cb == _T_33 ? _ram_T_363[287:0] : _GEN_13587; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14638 = 10'h1cc == _T_33 ? _ram_T_363[287:0] : _GEN_13588; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14639 = 10'h1cd == _T_33 ? _ram_T_363[287:0] : _GEN_13589; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14640 = 10'h1ce == _T_33 ? _ram_T_363[287:0] : _GEN_13590; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14641 = 10'h1cf == _T_33 ? _ram_T_363[287:0] : _GEN_13591; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14642 = 10'h1d0 == _T_33 ? _ram_T_363[287:0] : _GEN_13592; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14643 = 10'h1d1 == _T_33 ? _ram_T_363[287:0] : _GEN_13593; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14644 = 10'h1d2 == _T_33 ? _ram_T_363[287:0] : _GEN_13594; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14645 = 10'h1d3 == _T_33 ? _ram_T_363[287:0] : _GEN_13595; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14646 = 10'h1d4 == _T_33 ? _ram_T_363[287:0] : _GEN_13596; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14647 = 10'h1d5 == _T_33 ? _ram_T_363[287:0] : _GEN_13597; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14648 = 10'h1d6 == _T_33 ? _ram_T_363[287:0] : _GEN_13598; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14649 = 10'h1d7 == _T_33 ? _ram_T_363[287:0] : _GEN_13599; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14650 = 10'h1d8 == _T_33 ? _ram_T_363[287:0] : _GEN_13600; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14651 = 10'h1d9 == _T_33 ? _ram_T_363[287:0] : _GEN_13601; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14652 = 10'h1da == _T_33 ? _ram_T_363[287:0] : _GEN_13602; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14653 = 10'h1db == _T_33 ? _ram_T_363[287:0] : _GEN_13603; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14654 = 10'h1dc == _T_33 ? _ram_T_363[287:0] : _GEN_13604; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14655 = 10'h1dd == _T_33 ? _ram_T_363[287:0] : _GEN_13605; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14656 = 10'h1de == _T_33 ? _ram_T_363[287:0] : _GEN_13606; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14657 = 10'h1df == _T_33 ? _ram_T_363[287:0] : _GEN_13607; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14658 = 10'h1e0 == _T_33 ? _ram_T_363[287:0] : _GEN_13608; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14659 = 10'h1e1 == _T_33 ? _ram_T_363[287:0] : _GEN_13609; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14660 = 10'h1e2 == _T_33 ? _ram_T_363[287:0] : _GEN_13610; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14661 = 10'h1e3 == _T_33 ? _ram_T_363[287:0] : _GEN_13611; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14662 = 10'h1e4 == _T_33 ? _ram_T_363[287:0] : _GEN_13612; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14663 = 10'h1e5 == _T_33 ? _ram_T_363[287:0] : _GEN_13613; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14664 = 10'h1e6 == _T_33 ? _ram_T_363[287:0] : _GEN_13614; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14665 = 10'h1e7 == _T_33 ? _ram_T_363[287:0] : _GEN_13615; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14666 = 10'h1e8 == _T_33 ? _ram_T_363[287:0] : _GEN_13616; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14667 = 10'h1e9 == _T_33 ? _ram_T_363[287:0] : _GEN_13617; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14668 = 10'h1ea == _T_33 ? _ram_T_363[287:0] : _GEN_13618; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14669 = 10'h1eb == _T_33 ? _ram_T_363[287:0] : _GEN_13619; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14670 = 10'h1ec == _T_33 ? _ram_T_363[287:0] : _GEN_13620; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14671 = 10'h1ed == _T_33 ? _ram_T_363[287:0] : _GEN_13621; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14672 = 10'h1ee == _T_33 ? _ram_T_363[287:0] : _GEN_13622; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14673 = 10'h1ef == _T_33 ? _ram_T_363[287:0] : _GEN_13623; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14674 = 10'h1f0 == _T_33 ? _ram_T_363[287:0] : _GEN_13624; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14675 = 10'h1f1 == _T_33 ? _ram_T_363[287:0] : _GEN_13625; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14676 = 10'h1f2 == _T_33 ? _ram_T_363[287:0] : _GEN_13626; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14677 = 10'h1f3 == _T_33 ? _ram_T_363[287:0] : _GEN_13627; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14678 = 10'h1f4 == _T_33 ? _ram_T_363[287:0] : _GEN_13628; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14679 = 10'h1f5 == _T_33 ? _ram_T_363[287:0] : _GEN_13629; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14680 = 10'h1f6 == _T_33 ? _ram_T_363[287:0] : _GEN_13630; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14681 = 10'h1f7 == _T_33 ? _ram_T_363[287:0] : _GEN_13631; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14682 = 10'h1f8 == _T_33 ? _ram_T_363[287:0] : _GEN_13632; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14683 = 10'h1f9 == _T_33 ? _ram_T_363[287:0] : _GEN_13633; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14684 = 10'h1fa == _T_33 ? _ram_T_363[287:0] : _GEN_13634; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14685 = 10'h1fb == _T_33 ? _ram_T_363[287:0] : _GEN_13635; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14686 = 10'h1fc == _T_33 ? _ram_T_363[287:0] : _GEN_13636; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14687 = 10'h1fd == _T_33 ? _ram_T_363[287:0] : _GEN_13637; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14688 = 10'h1fe == _T_33 ? _ram_T_363[287:0] : _GEN_13638; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14689 = 10'h1ff == _T_33 ? _ram_T_363[287:0] : _GEN_13639; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14690 = 10'h200 == _T_33 ? _ram_T_363[287:0] : _GEN_13640; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14691 = 10'h201 == _T_33 ? _ram_T_363[287:0] : _GEN_13641; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14692 = 10'h202 == _T_33 ? _ram_T_363[287:0] : _GEN_13642; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14693 = 10'h203 == _T_33 ? _ram_T_363[287:0] : _GEN_13643; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14694 = 10'h204 == _T_33 ? _ram_T_363[287:0] : _GEN_13644; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14695 = 10'h205 == _T_33 ? _ram_T_363[287:0] : _GEN_13645; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14696 = 10'h206 == _T_33 ? _ram_T_363[287:0] : _GEN_13646; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14697 = 10'h207 == _T_33 ? _ram_T_363[287:0] : _GEN_13647; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14698 = 10'h208 == _T_33 ? _ram_T_363[287:0] : _GEN_13648; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14699 = 10'h209 == _T_33 ? _ram_T_363[287:0] : _GEN_13649; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14700 = 10'h20a == _T_33 ? _ram_T_363[287:0] : _GEN_13650; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14701 = 10'h20b == _T_33 ? _ram_T_363[287:0] : _GEN_13651; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_14702 = 10'h20c == _T_33 ? _ram_T_363[287:0] : _GEN_13652; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_35 = h + 10'he; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_14 = vga_mem_ram_MPORT_126_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_14 = vga_mem_ram_MPORT_127_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_14 = vga_mem_ram_MPORT_128_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_14 = vga_mem_ram_MPORT_129_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_14 = vga_mem_ram_MPORT_130_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_14 = vga_mem_ram_MPORT_131_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_14 = vga_mem_ram_MPORT_132_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_14 = vga_mem_ram_MPORT_133_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_14 = vga_mem_ram_MPORT_134_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_384 = {278'h0,ram_hi_hi_hi_lo_14,ram_hi_hi_lo_14,ram_hi_lo_hi_14,ram_hi_lo_lo_14,
    ram_lo_hi_hi_hi_14,ram_lo_hi_hi_lo_14,ram_lo_hi_lo_14,ram_lo_lo_hi_14,ram_lo_lo_lo_14}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19088 = {{8191'd0}, _ram_T_384}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_388 = _GEN_19088 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_14704 = 10'h1 == _T_35 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14705 = 10'h2 == _T_35 ? ram_2 : _GEN_14704; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14706 = 10'h3 == _T_35 ? ram_3 : _GEN_14705; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14707 = 10'h4 == _T_35 ? ram_4 : _GEN_14706; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14708 = 10'h5 == _T_35 ? ram_5 : _GEN_14707; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14709 = 10'h6 == _T_35 ? ram_6 : _GEN_14708; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14710 = 10'h7 == _T_35 ? ram_7 : _GEN_14709; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14711 = 10'h8 == _T_35 ? ram_8 : _GEN_14710; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14712 = 10'h9 == _T_35 ? ram_9 : _GEN_14711; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14713 = 10'ha == _T_35 ? ram_10 : _GEN_14712; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14714 = 10'hb == _T_35 ? ram_11 : _GEN_14713; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14715 = 10'hc == _T_35 ? ram_12 : _GEN_14714; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14716 = 10'hd == _T_35 ? ram_13 : _GEN_14715; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14717 = 10'he == _T_35 ? ram_14 : _GEN_14716; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14718 = 10'hf == _T_35 ? ram_15 : _GEN_14717; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14719 = 10'h10 == _T_35 ? ram_16 : _GEN_14718; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14720 = 10'h11 == _T_35 ? ram_17 : _GEN_14719; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14721 = 10'h12 == _T_35 ? ram_18 : _GEN_14720; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14722 = 10'h13 == _T_35 ? ram_19 : _GEN_14721; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14723 = 10'h14 == _T_35 ? ram_20 : _GEN_14722; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14724 = 10'h15 == _T_35 ? ram_21 : _GEN_14723; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14725 = 10'h16 == _T_35 ? ram_22 : _GEN_14724; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14726 = 10'h17 == _T_35 ? ram_23 : _GEN_14725; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14727 = 10'h18 == _T_35 ? ram_24 : _GEN_14726; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14728 = 10'h19 == _T_35 ? ram_25 : _GEN_14727; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14729 = 10'h1a == _T_35 ? ram_26 : _GEN_14728; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14730 = 10'h1b == _T_35 ? ram_27 : _GEN_14729; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14731 = 10'h1c == _T_35 ? ram_28 : _GEN_14730; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14732 = 10'h1d == _T_35 ? ram_29 : _GEN_14731; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14733 = 10'h1e == _T_35 ? ram_30 : _GEN_14732; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14734 = 10'h1f == _T_35 ? ram_31 : _GEN_14733; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14735 = 10'h20 == _T_35 ? ram_32 : _GEN_14734; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14736 = 10'h21 == _T_35 ? ram_33 : _GEN_14735; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14737 = 10'h22 == _T_35 ? ram_34 : _GEN_14736; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14738 = 10'h23 == _T_35 ? ram_35 : _GEN_14737; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14739 = 10'h24 == _T_35 ? ram_36 : _GEN_14738; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14740 = 10'h25 == _T_35 ? ram_37 : _GEN_14739; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14741 = 10'h26 == _T_35 ? ram_38 : _GEN_14740; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14742 = 10'h27 == _T_35 ? ram_39 : _GEN_14741; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14743 = 10'h28 == _T_35 ? ram_40 : _GEN_14742; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14744 = 10'h29 == _T_35 ? ram_41 : _GEN_14743; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14745 = 10'h2a == _T_35 ? ram_42 : _GEN_14744; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14746 = 10'h2b == _T_35 ? ram_43 : _GEN_14745; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14747 = 10'h2c == _T_35 ? ram_44 : _GEN_14746; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14748 = 10'h2d == _T_35 ? ram_45 : _GEN_14747; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14749 = 10'h2e == _T_35 ? ram_46 : _GEN_14748; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14750 = 10'h2f == _T_35 ? ram_47 : _GEN_14749; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14751 = 10'h30 == _T_35 ? ram_48 : _GEN_14750; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14752 = 10'h31 == _T_35 ? ram_49 : _GEN_14751; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14753 = 10'h32 == _T_35 ? ram_50 : _GEN_14752; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14754 = 10'h33 == _T_35 ? ram_51 : _GEN_14753; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14755 = 10'h34 == _T_35 ? ram_52 : _GEN_14754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14756 = 10'h35 == _T_35 ? ram_53 : _GEN_14755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14757 = 10'h36 == _T_35 ? ram_54 : _GEN_14756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14758 = 10'h37 == _T_35 ? ram_55 : _GEN_14757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14759 = 10'h38 == _T_35 ? ram_56 : _GEN_14758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14760 = 10'h39 == _T_35 ? ram_57 : _GEN_14759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14761 = 10'h3a == _T_35 ? ram_58 : _GEN_14760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14762 = 10'h3b == _T_35 ? ram_59 : _GEN_14761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14763 = 10'h3c == _T_35 ? ram_60 : _GEN_14762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14764 = 10'h3d == _T_35 ? ram_61 : _GEN_14763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14765 = 10'h3e == _T_35 ? ram_62 : _GEN_14764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14766 = 10'h3f == _T_35 ? ram_63 : _GEN_14765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14767 = 10'h40 == _T_35 ? ram_64 : _GEN_14766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14768 = 10'h41 == _T_35 ? ram_65 : _GEN_14767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14769 = 10'h42 == _T_35 ? ram_66 : _GEN_14768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14770 = 10'h43 == _T_35 ? ram_67 : _GEN_14769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14771 = 10'h44 == _T_35 ? ram_68 : _GEN_14770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14772 = 10'h45 == _T_35 ? ram_69 : _GEN_14771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14773 = 10'h46 == _T_35 ? ram_70 : _GEN_14772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14774 = 10'h47 == _T_35 ? ram_71 : _GEN_14773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14775 = 10'h48 == _T_35 ? ram_72 : _GEN_14774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14776 = 10'h49 == _T_35 ? ram_73 : _GEN_14775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14777 = 10'h4a == _T_35 ? ram_74 : _GEN_14776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14778 = 10'h4b == _T_35 ? ram_75 : _GEN_14777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14779 = 10'h4c == _T_35 ? ram_76 : _GEN_14778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14780 = 10'h4d == _T_35 ? ram_77 : _GEN_14779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14781 = 10'h4e == _T_35 ? ram_78 : _GEN_14780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14782 = 10'h4f == _T_35 ? ram_79 : _GEN_14781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14783 = 10'h50 == _T_35 ? ram_80 : _GEN_14782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14784 = 10'h51 == _T_35 ? ram_81 : _GEN_14783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14785 = 10'h52 == _T_35 ? ram_82 : _GEN_14784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14786 = 10'h53 == _T_35 ? ram_83 : _GEN_14785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14787 = 10'h54 == _T_35 ? ram_84 : _GEN_14786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14788 = 10'h55 == _T_35 ? ram_85 : _GEN_14787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14789 = 10'h56 == _T_35 ? ram_86 : _GEN_14788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14790 = 10'h57 == _T_35 ? ram_87 : _GEN_14789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14791 = 10'h58 == _T_35 ? ram_88 : _GEN_14790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14792 = 10'h59 == _T_35 ? ram_89 : _GEN_14791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14793 = 10'h5a == _T_35 ? ram_90 : _GEN_14792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14794 = 10'h5b == _T_35 ? ram_91 : _GEN_14793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14795 = 10'h5c == _T_35 ? ram_92 : _GEN_14794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14796 = 10'h5d == _T_35 ? ram_93 : _GEN_14795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14797 = 10'h5e == _T_35 ? ram_94 : _GEN_14796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14798 = 10'h5f == _T_35 ? ram_95 : _GEN_14797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14799 = 10'h60 == _T_35 ? ram_96 : _GEN_14798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14800 = 10'h61 == _T_35 ? ram_97 : _GEN_14799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14801 = 10'h62 == _T_35 ? ram_98 : _GEN_14800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14802 = 10'h63 == _T_35 ? ram_99 : _GEN_14801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14803 = 10'h64 == _T_35 ? ram_100 : _GEN_14802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14804 = 10'h65 == _T_35 ? ram_101 : _GEN_14803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14805 = 10'h66 == _T_35 ? ram_102 : _GEN_14804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14806 = 10'h67 == _T_35 ? ram_103 : _GEN_14805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14807 = 10'h68 == _T_35 ? ram_104 : _GEN_14806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14808 = 10'h69 == _T_35 ? ram_105 : _GEN_14807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14809 = 10'h6a == _T_35 ? ram_106 : _GEN_14808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14810 = 10'h6b == _T_35 ? ram_107 : _GEN_14809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14811 = 10'h6c == _T_35 ? ram_108 : _GEN_14810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14812 = 10'h6d == _T_35 ? ram_109 : _GEN_14811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14813 = 10'h6e == _T_35 ? ram_110 : _GEN_14812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14814 = 10'h6f == _T_35 ? ram_111 : _GEN_14813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14815 = 10'h70 == _T_35 ? ram_112 : _GEN_14814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14816 = 10'h71 == _T_35 ? ram_113 : _GEN_14815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14817 = 10'h72 == _T_35 ? ram_114 : _GEN_14816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14818 = 10'h73 == _T_35 ? ram_115 : _GEN_14817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14819 = 10'h74 == _T_35 ? ram_116 : _GEN_14818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14820 = 10'h75 == _T_35 ? ram_117 : _GEN_14819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14821 = 10'h76 == _T_35 ? ram_118 : _GEN_14820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14822 = 10'h77 == _T_35 ? ram_119 : _GEN_14821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14823 = 10'h78 == _T_35 ? ram_120 : _GEN_14822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14824 = 10'h79 == _T_35 ? ram_121 : _GEN_14823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14825 = 10'h7a == _T_35 ? ram_122 : _GEN_14824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14826 = 10'h7b == _T_35 ? ram_123 : _GEN_14825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14827 = 10'h7c == _T_35 ? ram_124 : _GEN_14826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14828 = 10'h7d == _T_35 ? ram_125 : _GEN_14827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14829 = 10'h7e == _T_35 ? ram_126 : _GEN_14828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14830 = 10'h7f == _T_35 ? ram_127 : _GEN_14829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14831 = 10'h80 == _T_35 ? ram_128 : _GEN_14830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14832 = 10'h81 == _T_35 ? ram_129 : _GEN_14831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14833 = 10'h82 == _T_35 ? ram_130 : _GEN_14832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14834 = 10'h83 == _T_35 ? ram_131 : _GEN_14833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14835 = 10'h84 == _T_35 ? ram_132 : _GEN_14834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14836 = 10'h85 == _T_35 ? ram_133 : _GEN_14835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14837 = 10'h86 == _T_35 ? ram_134 : _GEN_14836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14838 = 10'h87 == _T_35 ? ram_135 : _GEN_14837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14839 = 10'h88 == _T_35 ? ram_136 : _GEN_14838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14840 = 10'h89 == _T_35 ? ram_137 : _GEN_14839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14841 = 10'h8a == _T_35 ? ram_138 : _GEN_14840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14842 = 10'h8b == _T_35 ? ram_139 : _GEN_14841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14843 = 10'h8c == _T_35 ? ram_140 : _GEN_14842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14844 = 10'h8d == _T_35 ? ram_141 : _GEN_14843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14845 = 10'h8e == _T_35 ? ram_142 : _GEN_14844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14846 = 10'h8f == _T_35 ? ram_143 : _GEN_14845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14847 = 10'h90 == _T_35 ? ram_144 : _GEN_14846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14848 = 10'h91 == _T_35 ? ram_145 : _GEN_14847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14849 = 10'h92 == _T_35 ? ram_146 : _GEN_14848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14850 = 10'h93 == _T_35 ? ram_147 : _GEN_14849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14851 = 10'h94 == _T_35 ? ram_148 : _GEN_14850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14852 = 10'h95 == _T_35 ? ram_149 : _GEN_14851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14853 = 10'h96 == _T_35 ? ram_150 : _GEN_14852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14854 = 10'h97 == _T_35 ? ram_151 : _GEN_14853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14855 = 10'h98 == _T_35 ? ram_152 : _GEN_14854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14856 = 10'h99 == _T_35 ? ram_153 : _GEN_14855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14857 = 10'h9a == _T_35 ? ram_154 : _GEN_14856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14858 = 10'h9b == _T_35 ? ram_155 : _GEN_14857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14859 = 10'h9c == _T_35 ? ram_156 : _GEN_14858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14860 = 10'h9d == _T_35 ? ram_157 : _GEN_14859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14861 = 10'h9e == _T_35 ? ram_158 : _GEN_14860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14862 = 10'h9f == _T_35 ? ram_159 : _GEN_14861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14863 = 10'ha0 == _T_35 ? ram_160 : _GEN_14862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14864 = 10'ha1 == _T_35 ? ram_161 : _GEN_14863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14865 = 10'ha2 == _T_35 ? ram_162 : _GEN_14864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14866 = 10'ha3 == _T_35 ? ram_163 : _GEN_14865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14867 = 10'ha4 == _T_35 ? ram_164 : _GEN_14866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14868 = 10'ha5 == _T_35 ? ram_165 : _GEN_14867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14869 = 10'ha6 == _T_35 ? ram_166 : _GEN_14868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14870 = 10'ha7 == _T_35 ? ram_167 : _GEN_14869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14871 = 10'ha8 == _T_35 ? ram_168 : _GEN_14870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14872 = 10'ha9 == _T_35 ? ram_169 : _GEN_14871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14873 = 10'haa == _T_35 ? ram_170 : _GEN_14872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14874 = 10'hab == _T_35 ? ram_171 : _GEN_14873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14875 = 10'hac == _T_35 ? ram_172 : _GEN_14874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14876 = 10'had == _T_35 ? ram_173 : _GEN_14875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14877 = 10'hae == _T_35 ? ram_174 : _GEN_14876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14878 = 10'haf == _T_35 ? ram_175 : _GEN_14877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14879 = 10'hb0 == _T_35 ? ram_176 : _GEN_14878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14880 = 10'hb1 == _T_35 ? ram_177 : _GEN_14879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14881 = 10'hb2 == _T_35 ? ram_178 : _GEN_14880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14882 = 10'hb3 == _T_35 ? ram_179 : _GEN_14881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14883 = 10'hb4 == _T_35 ? ram_180 : _GEN_14882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14884 = 10'hb5 == _T_35 ? ram_181 : _GEN_14883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14885 = 10'hb6 == _T_35 ? ram_182 : _GEN_14884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14886 = 10'hb7 == _T_35 ? ram_183 : _GEN_14885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14887 = 10'hb8 == _T_35 ? ram_184 : _GEN_14886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14888 = 10'hb9 == _T_35 ? ram_185 : _GEN_14887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14889 = 10'hba == _T_35 ? ram_186 : _GEN_14888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14890 = 10'hbb == _T_35 ? ram_187 : _GEN_14889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14891 = 10'hbc == _T_35 ? ram_188 : _GEN_14890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14892 = 10'hbd == _T_35 ? ram_189 : _GEN_14891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14893 = 10'hbe == _T_35 ? ram_190 : _GEN_14892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14894 = 10'hbf == _T_35 ? ram_191 : _GEN_14893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14895 = 10'hc0 == _T_35 ? ram_192 : _GEN_14894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14896 = 10'hc1 == _T_35 ? ram_193 : _GEN_14895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14897 = 10'hc2 == _T_35 ? ram_194 : _GEN_14896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14898 = 10'hc3 == _T_35 ? ram_195 : _GEN_14897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14899 = 10'hc4 == _T_35 ? ram_196 : _GEN_14898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14900 = 10'hc5 == _T_35 ? ram_197 : _GEN_14899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14901 = 10'hc6 == _T_35 ? ram_198 : _GEN_14900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14902 = 10'hc7 == _T_35 ? ram_199 : _GEN_14901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14903 = 10'hc8 == _T_35 ? ram_200 : _GEN_14902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14904 = 10'hc9 == _T_35 ? ram_201 : _GEN_14903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14905 = 10'hca == _T_35 ? ram_202 : _GEN_14904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14906 = 10'hcb == _T_35 ? ram_203 : _GEN_14905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14907 = 10'hcc == _T_35 ? ram_204 : _GEN_14906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14908 = 10'hcd == _T_35 ? ram_205 : _GEN_14907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14909 = 10'hce == _T_35 ? ram_206 : _GEN_14908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14910 = 10'hcf == _T_35 ? ram_207 : _GEN_14909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14911 = 10'hd0 == _T_35 ? ram_208 : _GEN_14910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14912 = 10'hd1 == _T_35 ? ram_209 : _GEN_14911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14913 = 10'hd2 == _T_35 ? ram_210 : _GEN_14912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14914 = 10'hd3 == _T_35 ? ram_211 : _GEN_14913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14915 = 10'hd4 == _T_35 ? ram_212 : _GEN_14914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14916 = 10'hd5 == _T_35 ? ram_213 : _GEN_14915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14917 = 10'hd6 == _T_35 ? ram_214 : _GEN_14916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14918 = 10'hd7 == _T_35 ? ram_215 : _GEN_14917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14919 = 10'hd8 == _T_35 ? ram_216 : _GEN_14918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14920 = 10'hd9 == _T_35 ? ram_217 : _GEN_14919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14921 = 10'hda == _T_35 ? ram_218 : _GEN_14920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14922 = 10'hdb == _T_35 ? ram_219 : _GEN_14921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14923 = 10'hdc == _T_35 ? ram_220 : _GEN_14922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14924 = 10'hdd == _T_35 ? ram_221 : _GEN_14923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14925 = 10'hde == _T_35 ? ram_222 : _GEN_14924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14926 = 10'hdf == _T_35 ? ram_223 : _GEN_14925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14927 = 10'he0 == _T_35 ? ram_224 : _GEN_14926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14928 = 10'he1 == _T_35 ? ram_225 : _GEN_14927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14929 = 10'he2 == _T_35 ? ram_226 : _GEN_14928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14930 = 10'he3 == _T_35 ? ram_227 : _GEN_14929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14931 = 10'he4 == _T_35 ? ram_228 : _GEN_14930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14932 = 10'he5 == _T_35 ? ram_229 : _GEN_14931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14933 = 10'he6 == _T_35 ? ram_230 : _GEN_14932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14934 = 10'he7 == _T_35 ? ram_231 : _GEN_14933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14935 = 10'he8 == _T_35 ? ram_232 : _GEN_14934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14936 = 10'he9 == _T_35 ? ram_233 : _GEN_14935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14937 = 10'hea == _T_35 ? ram_234 : _GEN_14936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14938 = 10'heb == _T_35 ? ram_235 : _GEN_14937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14939 = 10'hec == _T_35 ? ram_236 : _GEN_14938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14940 = 10'hed == _T_35 ? ram_237 : _GEN_14939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14941 = 10'hee == _T_35 ? ram_238 : _GEN_14940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14942 = 10'hef == _T_35 ? ram_239 : _GEN_14941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14943 = 10'hf0 == _T_35 ? ram_240 : _GEN_14942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14944 = 10'hf1 == _T_35 ? ram_241 : _GEN_14943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14945 = 10'hf2 == _T_35 ? ram_242 : _GEN_14944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14946 = 10'hf3 == _T_35 ? ram_243 : _GEN_14945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14947 = 10'hf4 == _T_35 ? ram_244 : _GEN_14946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14948 = 10'hf5 == _T_35 ? ram_245 : _GEN_14947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14949 = 10'hf6 == _T_35 ? ram_246 : _GEN_14948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14950 = 10'hf7 == _T_35 ? ram_247 : _GEN_14949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14951 = 10'hf8 == _T_35 ? ram_248 : _GEN_14950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14952 = 10'hf9 == _T_35 ? ram_249 : _GEN_14951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14953 = 10'hfa == _T_35 ? ram_250 : _GEN_14952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14954 = 10'hfb == _T_35 ? ram_251 : _GEN_14953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14955 = 10'hfc == _T_35 ? ram_252 : _GEN_14954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14956 = 10'hfd == _T_35 ? ram_253 : _GEN_14955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14957 = 10'hfe == _T_35 ? ram_254 : _GEN_14956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14958 = 10'hff == _T_35 ? ram_255 : _GEN_14957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14959 = 10'h100 == _T_35 ? ram_256 : _GEN_14958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14960 = 10'h101 == _T_35 ? ram_257 : _GEN_14959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14961 = 10'h102 == _T_35 ? ram_258 : _GEN_14960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14962 = 10'h103 == _T_35 ? ram_259 : _GEN_14961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14963 = 10'h104 == _T_35 ? ram_260 : _GEN_14962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14964 = 10'h105 == _T_35 ? ram_261 : _GEN_14963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14965 = 10'h106 == _T_35 ? ram_262 : _GEN_14964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14966 = 10'h107 == _T_35 ? ram_263 : _GEN_14965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14967 = 10'h108 == _T_35 ? ram_264 : _GEN_14966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14968 = 10'h109 == _T_35 ? ram_265 : _GEN_14967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14969 = 10'h10a == _T_35 ? ram_266 : _GEN_14968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14970 = 10'h10b == _T_35 ? ram_267 : _GEN_14969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14971 = 10'h10c == _T_35 ? ram_268 : _GEN_14970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14972 = 10'h10d == _T_35 ? ram_269 : _GEN_14971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14973 = 10'h10e == _T_35 ? ram_270 : _GEN_14972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14974 = 10'h10f == _T_35 ? ram_271 : _GEN_14973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14975 = 10'h110 == _T_35 ? ram_272 : _GEN_14974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14976 = 10'h111 == _T_35 ? ram_273 : _GEN_14975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14977 = 10'h112 == _T_35 ? ram_274 : _GEN_14976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14978 = 10'h113 == _T_35 ? ram_275 : _GEN_14977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14979 = 10'h114 == _T_35 ? ram_276 : _GEN_14978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14980 = 10'h115 == _T_35 ? ram_277 : _GEN_14979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14981 = 10'h116 == _T_35 ? ram_278 : _GEN_14980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14982 = 10'h117 == _T_35 ? ram_279 : _GEN_14981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14983 = 10'h118 == _T_35 ? ram_280 : _GEN_14982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14984 = 10'h119 == _T_35 ? ram_281 : _GEN_14983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14985 = 10'h11a == _T_35 ? ram_282 : _GEN_14984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14986 = 10'h11b == _T_35 ? ram_283 : _GEN_14985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14987 = 10'h11c == _T_35 ? ram_284 : _GEN_14986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14988 = 10'h11d == _T_35 ? ram_285 : _GEN_14987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14989 = 10'h11e == _T_35 ? ram_286 : _GEN_14988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14990 = 10'h11f == _T_35 ? ram_287 : _GEN_14989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14991 = 10'h120 == _T_35 ? ram_288 : _GEN_14990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14992 = 10'h121 == _T_35 ? ram_289 : _GEN_14991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14993 = 10'h122 == _T_35 ? ram_290 : _GEN_14992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14994 = 10'h123 == _T_35 ? ram_291 : _GEN_14993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14995 = 10'h124 == _T_35 ? ram_292 : _GEN_14994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14996 = 10'h125 == _T_35 ? ram_293 : _GEN_14995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14997 = 10'h126 == _T_35 ? ram_294 : _GEN_14996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14998 = 10'h127 == _T_35 ? ram_295 : _GEN_14997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_14999 = 10'h128 == _T_35 ? ram_296 : _GEN_14998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15000 = 10'h129 == _T_35 ? ram_297 : _GEN_14999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15001 = 10'h12a == _T_35 ? ram_298 : _GEN_15000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15002 = 10'h12b == _T_35 ? ram_299 : _GEN_15001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15003 = 10'h12c == _T_35 ? ram_300 : _GEN_15002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15004 = 10'h12d == _T_35 ? ram_301 : _GEN_15003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15005 = 10'h12e == _T_35 ? ram_302 : _GEN_15004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15006 = 10'h12f == _T_35 ? ram_303 : _GEN_15005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15007 = 10'h130 == _T_35 ? ram_304 : _GEN_15006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15008 = 10'h131 == _T_35 ? ram_305 : _GEN_15007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15009 = 10'h132 == _T_35 ? ram_306 : _GEN_15008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15010 = 10'h133 == _T_35 ? ram_307 : _GEN_15009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15011 = 10'h134 == _T_35 ? ram_308 : _GEN_15010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15012 = 10'h135 == _T_35 ? ram_309 : _GEN_15011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15013 = 10'h136 == _T_35 ? ram_310 : _GEN_15012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15014 = 10'h137 == _T_35 ? ram_311 : _GEN_15013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15015 = 10'h138 == _T_35 ? ram_312 : _GEN_15014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15016 = 10'h139 == _T_35 ? ram_313 : _GEN_15015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15017 = 10'h13a == _T_35 ? ram_314 : _GEN_15016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15018 = 10'h13b == _T_35 ? ram_315 : _GEN_15017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15019 = 10'h13c == _T_35 ? ram_316 : _GEN_15018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15020 = 10'h13d == _T_35 ? ram_317 : _GEN_15019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15021 = 10'h13e == _T_35 ? ram_318 : _GEN_15020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15022 = 10'h13f == _T_35 ? ram_319 : _GEN_15021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15023 = 10'h140 == _T_35 ? ram_320 : _GEN_15022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15024 = 10'h141 == _T_35 ? ram_321 : _GEN_15023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15025 = 10'h142 == _T_35 ? ram_322 : _GEN_15024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15026 = 10'h143 == _T_35 ? ram_323 : _GEN_15025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15027 = 10'h144 == _T_35 ? ram_324 : _GEN_15026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15028 = 10'h145 == _T_35 ? ram_325 : _GEN_15027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15029 = 10'h146 == _T_35 ? ram_326 : _GEN_15028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15030 = 10'h147 == _T_35 ? ram_327 : _GEN_15029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15031 = 10'h148 == _T_35 ? ram_328 : _GEN_15030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15032 = 10'h149 == _T_35 ? ram_329 : _GEN_15031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15033 = 10'h14a == _T_35 ? ram_330 : _GEN_15032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15034 = 10'h14b == _T_35 ? ram_331 : _GEN_15033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15035 = 10'h14c == _T_35 ? ram_332 : _GEN_15034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15036 = 10'h14d == _T_35 ? ram_333 : _GEN_15035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15037 = 10'h14e == _T_35 ? ram_334 : _GEN_15036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15038 = 10'h14f == _T_35 ? ram_335 : _GEN_15037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15039 = 10'h150 == _T_35 ? ram_336 : _GEN_15038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15040 = 10'h151 == _T_35 ? ram_337 : _GEN_15039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15041 = 10'h152 == _T_35 ? ram_338 : _GEN_15040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15042 = 10'h153 == _T_35 ? ram_339 : _GEN_15041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15043 = 10'h154 == _T_35 ? ram_340 : _GEN_15042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15044 = 10'h155 == _T_35 ? ram_341 : _GEN_15043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15045 = 10'h156 == _T_35 ? ram_342 : _GEN_15044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15046 = 10'h157 == _T_35 ? ram_343 : _GEN_15045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15047 = 10'h158 == _T_35 ? ram_344 : _GEN_15046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15048 = 10'h159 == _T_35 ? ram_345 : _GEN_15047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15049 = 10'h15a == _T_35 ? ram_346 : _GEN_15048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15050 = 10'h15b == _T_35 ? ram_347 : _GEN_15049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15051 = 10'h15c == _T_35 ? ram_348 : _GEN_15050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15052 = 10'h15d == _T_35 ? ram_349 : _GEN_15051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15053 = 10'h15e == _T_35 ? ram_350 : _GEN_15052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15054 = 10'h15f == _T_35 ? ram_351 : _GEN_15053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15055 = 10'h160 == _T_35 ? ram_352 : _GEN_15054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15056 = 10'h161 == _T_35 ? ram_353 : _GEN_15055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15057 = 10'h162 == _T_35 ? ram_354 : _GEN_15056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15058 = 10'h163 == _T_35 ? ram_355 : _GEN_15057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15059 = 10'h164 == _T_35 ? ram_356 : _GEN_15058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15060 = 10'h165 == _T_35 ? ram_357 : _GEN_15059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15061 = 10'h166 == _T_35 ? ram_358 : _GEN_15060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15062 = 10'h167 == _T_35 ? ram_359 : _GEN_15061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15063 = 10'h168 == _T_35 ? ram_360 : _GEN_15062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15064 = 10'h169 == _T_35 ? ram_361 : _GEN_15063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15065 = 10'h16a == _T_35 ? ram_362 : _GEN_15064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15066 = 10'h16b == _T_35 ? ram_363 : _GEN_15065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15067 = 10'h16c == _T_35 ? ram_364 : _GEN_15066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15068 = 10'h16d == _T_35 ? ram_365 : _GEN_15067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15069 = 10'h16e == _T_35 ? ram_366 : _GEN_15068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15070 = 10'h16f == _T_35 ? ram_367 : _GEN_15069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15071 = 10'h170 == _T_35 ? ram_368 : _GEN_15070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15072 = 10'h171 == _T_35 ? ram_369 : _GEN_15071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15073 = 10'h172 == _T_35 ? ram_370 : _GEN_15072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15074 = 10'h173 == _T_35 ? ram_371 : _GEN_15073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15075 = 10'h174 == _T_35 ? ram_372 : _GEN_15074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15076 = 10'h175 == _T_35 ? ram_373 : _GEN_15075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15077 = 10'h176 == _T_35 ? ram_374 : _GEN_15076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15078 = 10'h177 == _T_35 ? ram_375 : _GEN_15077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15079 = 10'h178 == _T_35 ? ram_376 : _GEN_15078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15080 = 10'h179 == _T_35 ? ram_377 : _GEN_15079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15081 = 10'h17a == _T_35 ? ram_378 : _GEN_15080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15082 = 10'h17b == _T_35 ? ram_379 : _GEN_15081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15083 = 10'h17c == _T_35 ? ram_380 : _GEN_15082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15084 = 10'h17d == _T_35 ? ram_381 : _GEN_15083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15085 = 10'h17e == _T_35 ? ram_382 : _GEN_15084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15086 = 10'h17f == _T_35 ? ram_383 : _GEN_15085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15087 = 10'h180 == _T_35 ? ram_384 : _GEN_15086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15088 = 10'h181 == _T_35 ? ram_385 : _GEN_15087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15089 = 10'h182 == _T_35 ? ram_386 : _GEN_15088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15090 = 10'h183 == _T_35 ? ram_387 : _GEN_15089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15091 = 10'h184 == _T_35 ? ram_388 : _GEN_15090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15092 = 10'h185 == _T_35 ? ram_389 : _GEN_15091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15093 = 10'h186 == _T_35 ? ram_390 : _GEN_15092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15094 = 10'h187 == _T_35 ? ram_391 : _GEN_15093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15095 = 10'h188 == _T_35 ? ram_392 : _GEN_15094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15096 = 10'h189 == _T_35 ? ram_393 : _GEN_15095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15097 = 10'h18a == _T_35 ? ram_394 : _GEN_15096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15098 = 10'h18b == _T_35 ? ram_395 : _GEN_15097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15099 = 10'h18c == _T_35 ? ram_396 : _GEN_15098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15100 = 10'h18d == _T_35 ? ram_397 : _GEN_15099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15101 = 10'h18e == _T_35 ? ram_398 : _GEN_15100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15102 = 10'h18f == _T_35 ? ram_399 : _GEN_15101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15103 = 10'h190 == _T_35 ? ram_400 : _GEN_15102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15104 = 10'h191 == _T_35 ? ram_401 : _GEN_15103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15105 = 10'h192 == _T_35 ? ram_402 : _GEN_15104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15106 = 10'h193 == _T_35 ? ram_403 : _GEN_15105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15107 = 10'h194 == _T_35 ? ram_404 : _GEN_15106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15108 = 10'h195 == _T_35 ? ram_405 : _GEN_15107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15109 = 10'h196 == _T_35 ? ram_406 : _GEN_15108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15110 = 10'h197 == _T_35 ? ram_407 : _GEN_15109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15111 = 10'h198 == _T_35 ? ram_408 : _GEN_15110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15112 = 10'h199 == _T_35 ? ram_409 : _GEN_15111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15113 = 10'h19a == _T_35 ? ram_410 : _GEN_15112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15114 = 10'h19b == _T_35 ? ram_411 : _GEN_15113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15115 = 10'h19c == _T_35 ? ram_412 : _GEN_15114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15116 = 10'h19d == _T_35 ? ram_413 : _GEN_15115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15117 = 10'h19e == _T_35 ? ram_414 : _GEN_15116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15118 = 10'h19f == _T_35 ? ram_415 : _GEN_15117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15119 = 10'h1a0 == _T_35 ? ram_416 : _GEN_15118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15120 = 10'h1a1 == _T_35 ? ram_417 : _GEN_15119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15121 = 10'h1a2 == _T_35 ? ram_418 : _GEN_15120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15122 = 10'h1a3 == _T_35 ? ram_419 : _GEN_15121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15123 = 10'h1a4 == _T_35 ? ram_420 : _GEN_15122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15124 = 10'h1a5 == _T_35 ? ram_421 : _GEN_15123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15125 = 10'h1a6 == _T_35 ? ram_422 : _GEN_15124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15126 = 10'h1a7 == _T_35 ? ram_423 : _GEN_15125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15127 = 10'h1a8 == _T_35 ? ram_424 : _GEN_15126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15128 = 10'h1a9 == _T_35 ? ram_425 : _GEN_15127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15129 = 10'h1aa == _T_35 ? ram_426 : _GEN_15128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15130 = 10'h1ab == _T_35 ? ram_427 : _GEN_15129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15131 = 10'h1ac == _T_35 ? ram_428 : _GEN_15130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15132 = 10'h1ad == _T_35 ? ram_429 : _GEN_15131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15133 = 10'h1ae == _T_35 ? ram_430 : _GEN_15132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15134 = 10'h1af == _T_35 ? ram_431 : _GEN_15133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15135 = 10'h1b0 == _T_35 ? ram_432 : _GEN_15134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15136 = 10'h1b1 == _T_35 ? ram_433 : _GEN_15135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15137 = 10'h1b2 == _T_35 ? ram_434 : _GEN_15136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15138 = 10'h1b3 == _T_35 ? ram_435 : _GEN_15137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15139 = 10'h1b4 == _T_35 ? ram_436 : _GEN_15138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15140 = 10'h1b5 == _T_35 ? ram_437 : _GEN_15139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15141 = 10'h1b6 == _T_35 ? ram_438 : _GEN_15140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15142 = 10'h1b7 == _T_35 ? ram_439 : _GEN_15141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15143 = 10'h1b8 == _T_35 ? ram_440 : _GEN_15142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15144 = 10'h1b9 == _T_35 ? ram_441 : _GEN_15143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15145 = 10'h1ba == _T_35 ? ram_442 : _GEN_15144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15146 = 10'h1bb == _T_35 ? ram_443 : _GEN_15145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15147 = 10'h1bc == _T_35 ? ram_444 : _GEN_15146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15148 = 10'h1bd == _T_35 ? ram_445 : _GEN_15147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15149 = 10'h1be == _T_35 ? ram_446 : _GEN_15148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15150 = 10'h1bf == _T_35 ? ram_447 : _GEN_15149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15151 = 10'h1c0 == _T_35 ? ram_448 : _GEN_15150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15152 = 10'h1c1 == _T_35 ? ram_449 : _GEN_15151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15153 = 10'h1c2 == _T_35 ? ram_450 : _GEN_15152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15154 = 10'h1c3 == _T_35 ? ram_451 : _GEN_15153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15155 = 10'h1c4 == _T_35 ? ram_452 : _GEN_15154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15156 = 10'h1c5 == _T_35 ? ram_453 : _GEN_15155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15157 = 10'h1c6 == _T_35 ? ram_454 : _GEN_15156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15158 = 10'h1c7 == _T_35 ? ram_455 : _GEN_15157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15159 = 10'h1c8 == _T_35 ? ram_456 : _GEN_15158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15160 = 10'h1c9 == _T_35 ? ram_457 : _GEN_15159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15161 = 10'h1ca == _T_35 ? ram_458 : _GEN_15160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15162 = 10'h1cb == _T_35 ? ram_459 : _GEN_15161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15163 = 10'h1cc == _T_35 ? ram_460 : _GEN_15162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15164 = 10'h1cd == _T_35 ? ram_461 : _GEN_15163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15165 = 10'h1ce == _T_35 ? ram_462 : _GEN_15164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15166 = 10'h1cf == _T_35 ? ram_463 : _GEN_15165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15167 = 10'h1d0 == _T_35 ? ram_464 : _GEN_15166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15168 = 10'h1d1 == _T_35 ? ram_465 : _GEN_15167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15169 = 10'h1d2 == _T_35 ? ram_466 : _GEN_15168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15170 = 10'h1d3 == _T_35 ? ram_467 : _GEN_15169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15171 = 10'h1d4 == _T_35 ? ram_468 : _GEN_15170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15172 = 10'h1d5 == _T_35 ? ram_469 : _GEN_15171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15173 = 10'h1d6 == _T_35 ? ram_470 : _GEN_15172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15174 = 10'h1d7 == _T_35 ? ram_471 : _GEN_15173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15175 = 10'h1d8 == _T_35 ? ram_472 : _GEN_15174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15176 = 10'h1d9 == _T_35 ? ram_473 : _GEN_15175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15177 = 10'h1da == _T_35 ? ram_474 : _GEN_15176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15178 = 10'h1db == _T_35 ? ram_475 : _GEN_15177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15179 = 10'h1dc == _T_35 ? ram_476 : _GEN_15178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15180 = 10'h1dd == _T_35 ? ram_477 : _GEN_15179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15181 = 10'h1de == _T_35 ? ram_478 : _GEN_15180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15182 = 10'h1df == _T_35 ? ram_479 : _GEN_15181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15183 = 10'h1e0 == _T_35 ? ram_480 : _GEN_15182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15184 = 10'h1e1 == _T_35 ? ram_481 : _GEN_15183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15185 = 10'h1e2 == _T_35 ? ram_482 : _GEN_15184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15186 = 10'h1e3 == _T_35 ? ram_483 : _GEN_15185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15187 = 10'h1e4 == _T_35 ? ram_484 : _GEN_15186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15188 = 10'h1e5 == _T_35 ? ram_485 : _GEN_15187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15189 = 10'h1e6 == _T_35 ? ram_486 : _GEN_15188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15190 = 10'h1e7 == _T_35 ? ram_487 : _GEN_15189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15191 = 10'h1e8 == _T_35 ? ram_488 : _GEN_15190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15192 = 10'h1e9 == _T_35 ? ram_489 : _GEN_15191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15193 = 10'h1ea == _T_35 ? ram_490 : _GEN_15192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15194 = 10'h1eb == _T_35 ? ram_491 : _GEN_15193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15195 = 10'h1ec == _T_35 ? ram_492 : _GEN_15194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15196 = 10'h1ed == _T_35 ? ram_493 : _GEN_15195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15197 = 10'h1ee == _T_35 ? ram_494 : _GEN_15196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15198 = 10'h1ef == _T_35 ? ram_495 : _GEN_15197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15199 = 10'h1f0 == _T_35 ? ram_496 : _GEN_15198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15200 = 10'h1f1 == _T_35 ? ram_497 : _GEN_15199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15201 = 10'h1f2 == _T_35 ? ram_498 : _GEN_15200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15202 = 10'h1f3 == _T_35 ? ram_499 : _GEN_15201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15203 = 10'h1f4 == _T_35 ? ram_500 : _GEN_15202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15204 = 10'h1f5 == _T_35 ? ram_501 : _GEN_15203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15205 = 10'h1f6 == _T_35 ? ram_502 : _GEN_15204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15206 = 10'h1f7 == _T_35 ? ram_503 : _GEN_15205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15207 = 10'h1f8 == _T_35 ? ram_504 : _GEN_15206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15208 = 10'h1f9 == _T_35 ? ram_505 : _GEN_15207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15209 = 10'h1fa == _T_35 ? ram_506 : _GEN_15208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15210 = 10'h1fb == _T_35 ? ram_507 : _GEN_15209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15211 = 10'h1fc == _T_35 ? ram_508 : _GEN_15210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15212 = 10'h1fd == _T_35 ? ram_509 : _GEN_15211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15213 = 10'h1fe == _T_35 ? ram_510 : _GEN_15212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15214 = 10'h1ff == _T_35 ? ram_511 : _GEN_15213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15215 = 10'h200 == _T_35 ? ram_512 : _GEN_15214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15216 = 10'h201 == _T_35 ? ram_513 : _GEN_15215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15217 = 10'h202 == _T_35 ? ram_514 : _GEN_15216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15218 = 10'h203 == _T_35 ? ram_515 : _GEN_15217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15219 = 10'h204 == _T_35 ? ram_516 : _GEN_15218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15220 = 10'h205 == _T_35 ? ram_517 : _GEN_15219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15221 = 10'h206 == _T_35 ? ram_518 : _GEN_15220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15222 = 10'h207 == _T_35 ? ram_519 : _GEN_15221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15223 = 10'h208 == _T_35 ? ram_520 : _GEN_15222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15224 = 10'h209 == _T_35 ? ram_521 : _GEN_15223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15225 = 10'h20a == _T_35 ? ram_522 : _GEN_15224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15226 = 10'h20b == _T_35 ? ram_523 : _GEN_15225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15227 = 10'h20c == _T_35 ? ram_524 : _GEN_15226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19089 = {{8190'd0}, _GEN_15227}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_389 = _GEN_19089 ^ _ram_T_388; // @[vga.scala 64:41]
  wire [287:0] _GEN_15228 = 10'h0 == _T_35 ? _ram_T_389[287:0] : _GEN_14178; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15229 = 10'h1 == _T_35 ? _ram_T_389[287:0] : _GEN_14179; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15230 = 10'h2 == _T_35 ? _ram_T_389[287:0] : _GEN_14180; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15231 = 10'h3 == _T_35 ? _ram_T_389[287:0] : _GEN_14181; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15232 = 10'h4 == _T_35 ? _ram_T_389[287:0] : _GEN_14182; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15233 = 10'h5 == _T_35 ? _ram_T_389[287:0] : _GEN_14183; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15234 = 10'h6 == _T_35 ? _ram_T_389[287:0] : _GEN_14184; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15235 = 10'h7 == _T_35 ? _ram_T_389[287:0] : _GEN_14185; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15236 = 10'h8 == _T_35 ? _ram_T_389[287:0] : _GEN_14186; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15237 = 10'h9 == _T_35 ? _ram_T_389[287:0] : _GEN_14187; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15238 = 10'ha == _T_35 ? _ram_T_389[287:0] : _GEN_14188; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15239 = 10'hb == _T_35 ? _ram_T_389[287:0] : _GEN_14189; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15240 = 10'hc == _T_35 ? _ram_T_389[287:0] : _GEN_14190; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15241 = 10'hd == _T_35 ? _ram_T_389[287:0] : _GEN_14191; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15242 = 10'he == _T_35 ? _ram_T_389[287:0] : _GEN_14192; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15243 = 10'hf == _T_35 ? _ram_T_389[287:0] : _GEN_14193; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15244 = 10'h10 == _T_35 ? _ram_T_389[287:0] : _GEN_14194; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15245 = 10'h11 == _T_35 ? _ram_T_389[287:0] : _GEN_14195; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15246 = 10'h12 == _T_35 ? _ram_T_389[287:0] : _GEN_14196; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15247 = 10'h13 == _T_35 ? _ram_T_389[287:0] : _GEN_14197; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15248 = 10'h14 == _T_35 ? _ram_T_389[287:0] : _GEN_14198; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15249 = 10'h15 == _T_35 ? _ram_T_389[287:0] : _GEN_14199; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15250 = 10'h16 == _T_35 ? _ram_T_389[287:0] : _GEN_14200; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15251 = 10'h17 == _T_35 ? _ram_T_389[287:0] : _GEN_14201; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15252 = 10'h18 == _T_35 ? _ram_T_389[287:0] : _GEN_14202; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15253 = 10'h19 == _T_35 ? _ram_T_389[287:0] : _GEN_14203; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15254 = 10'h1a == _T_35 ? _ram_T_389[287:0] : _GEN_14204; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15255 = 10'h1b == _T_35 ? _ram_T_389[287:0] : _GEN_14205; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15256 = 10'h1c == _T_35 ? _ram_T_389[287:0] : _GEN_14206; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15257 = 10'h1d == _T_35 ? _ram_T_389[287:0] : _GEN_14207; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15258 = 10'h1e == _T_35 ? _ram_T_389[287:0] : _GEN_14208; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15259 = 10'h1f == _T_35 ? _ram_T_389[287:0] : _GEN_14209; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15260 = 10'h20 == _T_35 ? _ram_T_389[287:0] : _GEN_14210; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15261 = 10'h21 == _T_35 ? _ram_T_389[287:0] : _GEN_14211; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15262 = 10'h22 == _T_35 ? _ram_T_389[287:0] : _GEN_14212; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15263 = 10'h23 == _T_35 ? _ram_T_389[287:0] : _GEN_14213; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15264 = 10'h24 == _T_35 ? _ram_T_389[287:0] : _GEN_14214; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15265 = 10'h25 == _T_35 ? _ram_T_389[287:0] : _GEN_14215; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15266 = 10'h26 == _T_35 ? _ram_T_389[287:0] : _GEN_14216; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15267 = 10'h27 == _T_35 ? _ram_T_389[287:0] : _GEN_14217; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15268 = 10'h28 == _T_35 ? _ram_T_389[287:0] : _GEN_14218; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15269 = 10'h29 == _T_35 ? _ram_T_389[287:0] : _GEN_14219; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15270 = 10'h2a == _T_35 ? _ram_T_389[287:0] : _GEN_14220; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15271 = 10'h2b == _T_35 ? _ram_T_389[287:0] : _GEN_14221; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15272 = 10'h2c == _T_35 ? _ram_T_389[287:0] : _GEN_14222; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15273 = 10'h2d == _T_35 ? _ram_T_389[287:0] : _GEN_14223; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15274 = 10'h2e == _T_35 ? _ram_T_389[287:0] : _GEN_14224; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15275 = 10'h2f == _T_35 ? _ram_T_389[287:0] : _GEN_14225; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15276 = 10'h30 == _T_35 ? _ram_T_389[287:0] : _GEN_14226; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15277 = 10'h31 == _T_35 ? _ram_T_389[287:0] : _GEN_14227; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15278 = 10'h32 == _T_35 ? _ram_T_389[287:0] : _GEN_14228; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15279 = 10'h33 == _T_35 ? _ram_T_389[287:0] : _GEN_14229; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15280 = 10'h34 == _T_35 ? _ram_T_389[287:0] : _GEN_14230; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15281 = 10'h35 == _T_35 ? _ram_T_389[287:0] : _GEN_14231; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15282 = 10'h36 == _T_35 ? _ram_T_389[287:0] : _GEN_14232; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15283 = 10'h37 == _T_35 ? _ram_T_389[287:0] : _GEN_14233; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15284 = 10'h38 == _T_35 ? _ram_T_389[287:0] : _GEN_14234; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15285 = 10'h39 == _T_35 ? _ram_T_389[287:0] : _GEN_14235; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15286 = 10'h3a == _T_35 ? _ram_T_389[287:0] : _GEN_14236; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15287 = 10'h3b == _T_35 ? _ram_T_389[287:0] : _GEN_14237; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15288 = 10'h3c == _T_35 ? _ram_T_389[287:0] : _GEN_14238; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15289 = 10'h3d == _T_35 ? _ram_T_389[287:0] : _GEN_14239; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15290 = 10'h3e == _T_35 ? _ram_T_389[287:0] : _GEN_14240; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15291 = 10'h3f == _T_35 ? _ram_T_389[287:0] : _GEN_14241; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15292 = 10'h40 == _T_35 ? _ram_T_389[287:0] : _GEN_14242; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15293 = 10'h41 == _T_35 ? _ram_T_389[287:0] : _GEN_14243; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15294 = 10'h42 == _T_35 ? _ram_T_389[287:0] : _GEN_14244; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15295 = 10'h43 == _T_35 ? _ram_T_389[287:0] : _GEN_14245; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15296 = 10'h44 == _T_35 ? _ram_T_389[287:0] : _GEN_14246; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15297 = 10'h45 == _T_35 ? _ram_T_389[287:0] : _GEN_14247; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15298 = 10'h46 == _T_35 ? _ram_T_389[287:0] : _GEN_14248; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15299 = 10'h47 == _T_35 ? _ram_T_389[287:0] : _GEN_14249; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15300 = 10'h48 == _T_35 ? _ram_T_389[287:0] : _GEN_14250; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15301 = 10'h49 == _T_35 ? _ram_T_389[287:0] : _GEN_14251; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15302 = 10'h4a == _T_35 ? _ram_T_389[287:0] : _GEN_14252; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15303 = 10'h4b == _T_35 ? _ram_T_389[287:0] : _GEN_14253; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15304 = 10'h4c == _T_35 ? _ram_T_389[287:0] : _GEN_14254; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15305 = 10'h4d == _T_35 ? _ram_T_389[287:0] : _GEN_14255; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15306 = 10'h4e == _T_35 ? _ram_T_389[287:0] : _GEN_14256; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15307 = 10'h4f == _T_35 ? _ram_T_389[287:0] : _GEN_14257; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15308 = 10'h50 == _T_35 ? _ram_T_389[287:0] : _GEN_14258; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15309 = 10'h51 == _T_35 ? _ram_T_389[287:0] : _GEN_14259; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15310 = 10'h52 == _T_35 ? _ram_T_389[287:0] : _GEN_14260; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15311 = 10'h53 == _T_35 ? _ram_T_389[287:0] : _GEN_14261; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15312 = 10'h54 == _T_35 ? _ram_T_389[287:0] : _GEN_14262; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15313 = 10'h55 == _T_35 ? _ram_T_389[287:0] : _GEN_14263; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15314 = 10'h56 == _T_35 ? _ram_T_389[287:0] : _GEN_14264; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15315 = 10'h57 == _T_35 ? _ram_T_389[287:0] : _GEN_14265; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15316 = 10'h58 == _T_35 ? _ram_T_389[287:0] : _GEN_14266; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15317 = 10'h59 == _T_35 ? _ram_T_389[287:0] : _GEN_14267; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15318 = 10'h5a == _T_35 ? _ram_T_389[287:0] : _GEN_14268; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15319 = 10'h5b == _T_35 ? _ram_T_389[287:0] : _GEN_14269; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15320 = 10'h5c == _T_35 ? _ram_T_389[287:0] : _GEN_14270; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15321 = 10'h5d == _T_35 ? _ram_T_389[287:0] : _GEN_14271; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15322 = 10'h5e == _T_35 ? _ram_T_389[287:0] : _GEN_14272; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15323 = 10'h5f == _T_35 ? _ram_T_389[287:0] : _GEN_14273; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15324 = 10'h60 == _T_35 ? _ram_T_389[287:0] : _GEN_14274; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15325 = 10'h61 == _T_35 ? _ram_T_389[287:0] : _GEN_14275; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15326 = 10'h62 == _T_35 ? _ram_T_389[287:0] : _GEN_14276; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15327 = 10'h63 == _T_35 ? _ram_T_389[287:0] : _GEN_14277; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15328 = 10'h64 == _T_35 ? _ram_T_389[287:0] : _GEN_14278; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15329 = 10'h65 == _T_35 ? _ram_T_389[287:0] : _GEN_14279; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15330 = 10'h66 == _T_35 ? _ram_T_389[287:0] : _GEN_14280; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15331 = 10'h67 == _T_35 ? _ram_T_389[287:0] : _GEN_14281; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15332 = 10'h68 == _T_35 ? _ram_T_389[287:0] : _GEN_14282; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15333 = 10'h69 == _T_35 ? _ram_T_389[287:0] : _GEN_14283; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15334 = 10'h6a == _T_35 ? _ram_T_389[287:0] : _GEN_14284; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15335 = 10'h6b == _T_35 ? _ram_T_389[287:0] : _GEN_14285; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15336 = 10'h6c == _T_35 ? _ram_T_389[287:0] : _GEN_14286; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15337 = 10'h6d == _T_35 ? _ram_T_389[287:0] : _GEN_14287; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15338 = 10'h6e == _T_35 ? _ram_T_389[287:0] : _GEN_14288; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15339 = 10'h6f == _T_35 ? _ram_T_389[287:0] : _GEN_14289; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15340 = 10'h70 == _T_35 ? _ram_T_389[287:0] : _GEN_14290; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15341 = 10'h71 == _T_35 ? _ram_T_389[287:0] : _GEN_14291; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15342 = 10'h72 == _T_35 ? _ram_T_389[287:0] : _GEN_14292; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15343 = 10'h73 == _T_35 ? _ram_T_389[287:0] : _GEN_14293; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15344 = 10'h74 == _T_35 ? _ram_T_389[287:0] : _GEN_14294; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15345 = 10'h75 == _T_35 ? _ram_T_389[287:0] : _GEN_14295; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15346 = 10'h76 == _T_35 ? _ram_T_389[287:0] : _GEN_14296; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15347 = 10'h77 == _T_35 ? _ram_T_389[287:0] : _GEN_14297; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15348 = 10'h78 == _T_35 ? _ram_T_389[287:0] : _GEN_14298; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15349 = 10'h79 == _T_35 ? _ram_T_389[287:0] : _GEN_14299; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15350 = 10'h7a == _T_35 ? _ram_T_389[287:0] : _GEN_14300; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15351 = 10'h7b == _T_35 ? _ram_T_389[287:0] : _GEN_14301; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15352 = 10'h7c == _T_35 ? _ram_T_389[287:0] : _GEN_14302; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15353 = 10'h7d == _T_35 ? _ram_T_389[287:0] : _GEN_14303; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15354 = 10'h7e == _T_35 ? _ram_T_389[287:0] : _GEN_14304; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15355 = 10'h7f == _T_35 ? _ram_T_389[287:0] : _GEN_14305; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15356 = 10'h80 == _T_35 ? _ram_T_389[287:0] : _GEN_14306; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15357 = 10'h81 == _T_35 ? _ram_T_389[287:0] : _GEN_14307; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15358 = 10'h82 == _T_35 ? _ram_T_389[287:0] : _GEN_14308; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15359 = 10'h83 == _T_35 ? _ram_T_389[287:0] : _GEN_14309; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15360 = 10'h84 == _T_35 ? _ram_T_389[287:0] : _GEN_14310; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15361 = 10'h85 == _T_35 ? _ram_T_389[287:0] : _GEN_14311; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15362 = 10'h86 == _T_35 ? _ram_T_389[287:0] : _GEN_14312; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15363 = 10'h87 == _T_35 ? _ram_T_389[287:0] : _GEN_14313; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15364 = 10'h88 == _T_35 ? _ram_T_389[287:0] : _GEN_14314; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15365 = 10'h89 == _T_35 ? _ram_T_389[287:0] : _GEN_14315; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15366 = 10'h8a == _T_35 ? _ram_T_389[287:0] : _GEN_14316; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15367 = 10'h8b == _T_35 ? _ram_T_389[287:0] : _GEN_14317; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15368 = 10'h8c == _T_35 ? _ram_T_389[287:0] : _GEN_14318; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15369 = 10'h8d == _T_35 ? _ram_T_389[287:0] : _GEN_14319; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15370 = 10'h8e == _T_35 ? _ram_T_389[287:0] : _GEN_14320; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15371 = 10'h8f == _T_35 ? _ram_T_389[287:0] : _GEN_14321; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15372 = 10'h90 == _T_35 ? _ram_T_389[287:0] : _GEN_14322; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15373 = 10'h91 == _T_35 ? _ram_T_389[287:0] : _GEN_14323; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15374 = 10'h92 == _T_35 ? _ram_T_389[287:0] : _GEN_14324; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15375 = 10'h93 == _T_35 ? _ram_T_389[287:0] : _GEN_14325; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15376 = 10'h94 == _T_35 ? _ram_T_389[287:0] : _GEN_14326; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15377 = 10'h95 == _T_35 ? _ram_T_389[287:0] : _GEN_14327; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15378 = 10'h96 == _T_35 ? _ram_T_389[287:0] : _GEN_14328; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15379 = 10'h97 == _T_35 ? _ram_T_389[287:0] : _GEN_14329; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15380 = 10'h98 == _T_35 ? _ram_T_389[287:0] : _GEN_14330; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15381 = 10'h99 == _T_35 ? _ram_T_389[287:0] : _GEN_14331; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15382 = 10'h9a == _T_35 ? _ram_T_389[287:0] : _GEN_14332; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15383 = 10'h9b == _T_35 ? _ram_T_389[287:0] : _GEN_14333; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15384 = 10'h9c == _T_35 ? _ram_T_389[287:0] : _GEN_14334; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15385 = 10'h9d == _T_35 ? _ram_T_389[287:0] : _GEN_14335; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15386 = 10'h9e == _T_35 ? _ram_T_389[287:0] : _GEN_14336; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15387 = 10'h9f == _T_35 ? _ram_T_389[287:0] : _GEN_14337; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15388 = 10'ha0 == _T_35 ? _ram_T_389[287:0] : _GEN_14338; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15389 = 10'ha1 == _T_35 ? _ram_T_389[287:0] : _GEN_14339; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15390 = 10'ha2 == _T_35 ? _ram_T_389[287:0] : _GEN_14340; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15391 = 10'ha3 == _T_35 ? _ram_T_389[287:0] : _GEN_14341; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15392 = 10'ha4 == _T_35 ? _ram_T_389[287:0] : _GEN_14342; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15393 = 10'ha5 == _T_35 ? _ram_T_389[287:0] : _GEN_14343; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15394 = 10'ha6 == _T_35 ? _ram_T_389[287:0] : _GEN_14344; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15395 = 10'ha7 == _T_35 ? _ram_T_389[287:0] : _GEN_14345; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15396 = 10'ha8 == _T_35 ? _ram_T_389[287:0] : _GEN_14346; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15397 = 10'ha9 == _T_35 ? _ram_T_389[287:0] : _GEN_14347; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15398 = 10'haa == _T_35 ? _ram_T_389[287:0] : _GEN_14348; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15399 = 10'hab == _T_35 ? _ram_T_389[287:0] : _GEN_14349; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15400 = 10'hac == _T_35 ? _ram_T_389[287:0] : _GEN_14350; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15401 = 10'had == _T_35 ? _ram_T_389[287:0] : _GEN_14351; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15402 = 10'hae == _T_35 ? _ram_T_389[287:0] : _GEN_14352; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15403 = 10'haf == _T_35 ? _ram_T_389[287:0] : _GEN_14353; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15404 = 10'hb0 == _T_35 ? _ram_T_389[287:0] : _GEN_14354; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15405 = 10'hb1 == _T_35 ? _ram_T_389[287:0] : _GEN_14355; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15406 = 10'hb2 == _T_35 ? _ram_T_389[287:0] : _GEN_14356; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15407 = 10'hb3 == _T_35 ? _ram_T_389[287:0] : _GEN_14357; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15408 = 10'hb4 == _T_35 ? _ram_T_389[287:0] : _GEN_14358; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15409 = 10'hb5 == _T_35 ? _ram_T_389[287:0] : _GEN_14359; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15410 = 10'hb6 == _T_35 ? _ram_T_389[287:0] : _GEN_14360; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15411 = 10'hb7 == _T_35 ? _ram_T_389[287:0] : _GEN_14361; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15412 = 10'hb8 == _T_35 ? _ram_T_389[287:0] : _GEN_14362; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15413 = 10'hb9 == _T_35 ? _ram_T_389[287:0] : _GEN_14363; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15414 = 10'hba == _T_35 ? _ram_T_389[287:0] : _GEN_14364; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15415 = 10'hbb == _T_35 ? _ram_T_389[287:0] : _GEN_14365; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15416 = 10'hbc == _T_35 ? _ram_T_389[287:0] : _GEN_14366; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15417 = 10'hbd == _T_35 ? _ram_T_389[287:0] : _GEN_14367; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15418 = 10'hbe == _T_35 ? _ram_T_389[287:0] : _GEN_14368; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15419 = 10'hbf == _T_35 ? _ram_T_389[287:0] : _GEN_14369; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15420 = 10'hc0 == _T_35 ? _ram_T_389[287:0] : _GEN_14370; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15421 = 10'hc1 == _T_35 ? _ram_T_389[287:0] : _GEN_14371; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15422 = 10'hc2 == _T_35 ? _ram_T_389[287:0] : _GEN_14372; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15423 = 10'hc3 == _T_35 ? _ram_T_389[287:0] : _GEN_14373; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15424 = 10'hc4 == _T_35 ? _ram_T_389[287:0] : _GEN_14374; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15425 = 10'hc5 == _T_35 ? _ram_T_389[287:0] : _GEN_14375; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15426 = 10'hc6 == _T_35 ? _ram_T_389[287:0] : _GEN_14376; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15427 = 10'hc7 == _T_35 ? _ram_T_389[287:0] : _GEN_14377; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15428 = 10'hc8 == _T_35 ? _ram_T_389[287:0] : _GEN_14378; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15429 = 10'hc9 == _T_35 ? _ram_T_389[287:0] : _GEN_14379; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15430 = 10'hca == _T_35 ? _ram_T_389[287:0] : _GEN_14380; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15431 = 10'hcb == _T_35 ? _ram_T_389[287:0] : _GEN_14381; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15432 = 10'hcc == _T_35 ? _ram_T_389[287:0] : _GEN_14382; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15433 = 10'hcd == _T_35 ? _ram_T_389[287:0] : _GEN_14383; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15434 = 10'hce == _T_35 ? _ram_T_389[287:0] : _GEN_14384; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15435 = 10'hcf == _T_35 ? _ram_T_389[287:0] : _GEN_14385; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15436 = 10'hd0 == _T_35 ? _ram_T_389[287:0] : _GEN_14386; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15437 = 10'hd1 == _T_35 ? _ram_T_389[287:0] : _GEN_14387; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15438 = 10'hd2 == _T_35 ? _ram_T_389[287:0] : _GEN_14388; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15439 = 10'hd3 == _T_35 ? _ram_T_389[287:0] : _GEN_14389; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15440 = 10'hd4 == _T_35 ? _ram_T_389[287:0] : _GEN_14390; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15441 = 10'hd5 == _T_35 ? _ram_T_389[287:0] : _GEN_14391; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15442 = 10'hd6 == _T_35 ? _ram_T_389[287:0] : _GEN_14392; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15443 = 10'hd7 == _T_35 ? _ram_T_389[287:0] : _GEN_14393; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15444 = 10'hd8 == _T_35 ? _ram_T_389[287:0] : _GEN_14394; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15445 = 10'hd9 == _T_35 ? _ram_T_389[287:0] : _GEN_14395; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15446 = 10'hda == _T_35 ? _ram_T_389[287:0] : _GEN_14396; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15447 = 10'hdb == _T_35 ? _ram_T_389[287:0] : _GEN_14397; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15448 = 10'hdc == _T_35 ? _ram_T_389[287:0] : _GEN_14398; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15449 = 10'hdd == _T_35 ? _ram_T_389[287:0] : _GEN_14399; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15450 = 10'hde == _T_35 ? _ram_T_389[287:0] : _GEN_14400; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15451 = 10'hdf == _T_35 ? _ram_T_389[287:0] : _GEN_14401; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15452 = 10'he0 == _T_35 ? _ram_T_389[287:0] : _GEN_14402; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15453 = 10'he1 == _T_35 ? _ram_T_389[287:0] : _GEN_14403; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15454 = 10'he2 == _T_35 ? _ram_T_389[287:0] : _GEN_14404; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15455 = 10'he3 == _T_35 ? _ram_T_389[287:0] : _GEN_14405; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15456 = 10'he4 == _T_35 ? _ram_T_389[287:0] : _GEN_14406; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15457 = 10'he5 == _T_35 ? _ram_T_389[287:0] : _GEN_14407; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15458 = 10'he6 == _T_35 ? _ram_T_389[287:0] : _GEN_14408; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15459 = 10'he7 == _T_35 ? _ram_T_389[287:0] : _GEN_14409; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15460 = 10'he8 == _T_35 ? _ram_T_389[287:0] : _GEN_14410; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15461 = 10'he9 == _T_35 ? _ram_T_389[287:0] : _GEN_14411; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15462 = 10'hea == _T_35 ? _ram_T_389[287:0] : _GEN_14412; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15463 = 10'heb == _T_35 ? _ram_T_389[287:0] : _GEN_14413; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15464 = 10'hec == _T_35 ? _ram_T_389[287:0] : _GEN_14414; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15465 = 10'hed == _T_35 ? _ram_T_389[287:0] : _GEN_14415; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15466 = 10'hee == _T_35 ? _ram_T_389[287:0] : _GEN_14416; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15467 = 10'hef == _T_35 ? _ram_T_389[287:0] : _GEN_14417; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15468 = 10'hf0 == _T_35 ? _ram_T_389[287:0] : _GEN_14418; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15469 = 10'hf1 == _T_35 ? _ram_T_389[287:0] : _GEN_14419; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15470 = 10'hf2 == _T_35 ? _ram_T_389[287:0] : _GEN_14420; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15471 = 10'hf3 == _T_35 ? _ram_T_389[287:0] : _GEN_14421; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15472 = 10'hf4 == _T_35 ? _ram_T_389[287:0] : _GEN_14422; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15473 = 10'hf5 == _T_35 ? _ram_T_389[287:0] : _GEN_14423; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15474 = 10'hf6 == _T_35 ? _ram_T_389[287:0] : _GEN_14424; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15475 = 10'hf7 == _T_35 ? _ram_T_389[287:0] : _GEN_14425; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15476 = 10'hf8 == _T_35 ? _ram_T_389[287:0] : _GEN_14426; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15477 = 10'hf9 == _T_35 ? _ram_T_389[287:0] : _GEN_14427; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15478 = 10'hfa == _T_35 ? _ram_T_389[287:0] : _GEN_14428; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15479 = 10'hfb == _T_35 ? _ram_T_389[287:0] : _GEN_14429; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15480 = 10'hfc == _T_35 ? _ram_T_389[287:0] : _GEN_14430; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15481 = 10'hfd == _T_35 ? _ram_T_389[287:0] : _GEN_14431; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15482 = 10'hfe == _T_35 ? _ram_T_389[287:0] : _GEN_14432; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15483 = 10'hff == _T_35 ? _ram_T_389[287:0] : _GEN_14433; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15484 = 10'h100 == _T_35 ? _ram_T_389[287:0] : _GEN_14434; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15485 = 10'h101 == _T_35 ? _ram_T_389[287:0] : _GEN_14435; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15486 = 10'h102 == _T_35 ? _ram_T_389[287:0] : _GEN_14436; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15487 = 10'h103 == _T_35 ? _ram_T_389[287:0] : _GEN_14437; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15488 = 10'h104 == _T_35 ? _ram_T_389[287:0] : _GEN_14438; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15489 = 10'h105 == _T_35 ? _ram_T_389[287:0] : _GEN_14439; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15490 = 10'h106 == _T_35 ? _ram_T_389[287:0] : _GEN_14440; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15491 = 10'h107 == _T_35 ? _ram_T_389[287:0] : _GEN_14441; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15492 = 10'h108 == _T_35 ? _ram_T_389[287:0] : _GEN_14442; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15493 = 10'h109 == _T_35 ? _ram_T_389[287:0] : _GEN_14443; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15494 = 10'h10a == _T_35 ? _ram_T_389[287:0] : _GEN_14444; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15495 = 10'h10b == _T_35 ? _ram_T_389[287:0] : _GEN_14445; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15496 = 10'h10c == _T_35 ? _ram_T_389[287:0] : _GEN_14446; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15497 = 10'h10d == _T_35 ? _ram_T_389[287:0] : _GEN_14447; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15498 = 10'h10e == _T_35 ? _ram_T_389[287:0] : _GEN_14448; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15499 = 10'h10f == _T_35 ? _ram_T_389[287:0] : _GEN_14449; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15500 = 10'h110 == _T_35 ? _ram_T_389[287:0] : _GEN_14450; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15501 = 10'h111 == _T_35 ? _ram_T_389[287:0] : _GEN_14451; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15502 = 10'h112 == _T_35 ? _ram_T_389[287:0] : _GEN_14452; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15503 = 10'h113 == _T_35 ? _ram_T_389[287:0] : _GEN_14453; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15504 = 10'h114 == _T_35 ? _ram_T_389[287:0] : _GEN_14454; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15505 = 10'h115 == _T_35 ? _ram_T_389[287:0] : _GEN_14455; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15506 = 10'h116 == _T_35 ? _ram_T_389[287:0] : _GEN_14456; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15507 = 10'h117 == _T_35 ? _ram_T_389[287:0] : _GEN_14457; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15508 = 10'h118 == _T_35 ? _ram_T_389[287:0] : _GEN_14458; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15509 = 10'h119 == _T_35 ? _ram_T_389[287:0] : _GEN_14459; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15510 = 10'h11a == _T_35 ? _ram_T_389[287:0] : _GEN_14460; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15511 = 10'h11b == _T_35 ? _ram_T_389[287:0] : _GEN_14461; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15512 = 10'h11c == _T_35 ? _ram_T_389[287:0] : _GEN_14462; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15513 = 10'h11d == _T_35 ? _ram_T_389[287:0] : _GEN_14463; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15514 = 10'h11e == _T_35 ? _ram_T_389[287:0] : _GEN_14464; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15515 = 10'h11f == _T_35 ? _ram_T_389[287:0] : _GEN_14465; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15516 = 10'h120 == _T_35 ? _ram_T_389[287:0] : _GEN_14466; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15517 = 10'h121 == _T_35 ? _ram_T_389[287:0] : _GEN_14467; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15518 = 10'h122 == _T_35 ? _ram_T_389[287:0] : _GEN_14468; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15519 = 10'h123 == _T_35 ? _ram_T_389[287:0] : _GEN_14469; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15520 = 10'h124 == _T_35 ? _ram_T_389[287:0] : _GEN_14470; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15521 = 10'h125 == _T_35 ? _ram_T_389[287:0] : _GEN_14471; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15522 = 10'h126 == _T_35 ? _ram_T_389[287:0] : _GEN_14472; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15523 = 10'h127 == _T_35 ? _ram_T_389[287:0] : _GEN_14473; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15524 = 10'h128 == _T_35 ? _ram_T_389[287:0] : _GEN_14474; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15525 = 10'h129 == _T_35 ? _ram_T_389[287:0] : _GEN_14475; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15526 = 10'h12a == _T_35 ? _ram_T_389[287:0] : _GEN_14476; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15527 = 10'h12b == _T_35 ? _ram_T_389[287:0] : _GEN_14477; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15528 = 10'h12c == _T_35 ? _ram_T_389[287:0] : _GEN_14478; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15529 = 10'h12d == _T_35 ? _ram_T_389[287:0] : _GEN_14479; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15530 = 10'h12e == _T_35 ? _ram_T_389[287:0] : _GEN_14480; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15531 = 10'h12f == _T_35 ? _ram_T_389[287:0] : _GEN_14481; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15532 = 10'h130 == _T_35 ? _ram_T_389[287:0] : _GEN_14482; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15533 = 10'h131 == _T_35 ? _ram_T_389[287:0] : _GEN_14483; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15534 = 10'h132 == _T_35 ? _ram_T_389[287:0] : _GEN_14484; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15535 = 10'h133 == _T_35 ? _ram_T_389[287:0] : _GEN_14485; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15536 = 10'h134 == _T_35 ? _ram_T_389[287:0] : _GEN_14486; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15537 = 10'h135 == _T_35 ? _ram_T_389[287:0] : _GEN_14487; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15538 = 10'h136 == _T_35 ? _ram_T_389[287:0] : _GEN_14488; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15539 = 10'h137 == _T_35 ? _ram_T_389[287:0] : _GEN_14489; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15540 = 10'h138 == _T_35 ? _ram_T_389[287:0] : _GEN_14490; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15541 = 10'h139 == _T_35 ? _ram_T_389[287:0] : _GEN_14491; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15542 = 10'h13a == _T_35 ? _ram_T_389[287:0] : _GEN_14492; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15543 = 10'h13b == _T_35 ? _ram_T_389[287:0] : _GEN_14493; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15544 = 10'h13c == _T_35 ? _ram_T_389[287:0] : _GEN_14494; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15545 = 10'h13d == _T_35 ? _ram_T_389[287:0] : _GEN_14495; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15546 = 10'h13e == _T_35 ? _ram_T_389[287:0] : _GEN_14496; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15547 = 10'h13f == _T_35 ? _ram_T_389[287:0] : _GEN_14497; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15548 = 10'h140 == _T_35 ? _ram_T_389[287:0] : _GEN_14498; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15549 = 10'h141 == _T_35 ? _ram_T_389[287:0] : _GEN_14499; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15550 = 10'h142 == _T_35 ? _ram_T_389[287:0] : _GEN_14500; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15551 = 10'h143 == _T_35 ? _ram_T_389[287:0] : _GEN_14501; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15552 = 10'h144 == _T_35 ? _ram_T_389[287:0] : _GEN_14502; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15553 = 10'h145 == _T_35 ? _ram_T_389[287:0] : _GEN_14503; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15554 = 10'h146 == _T_35 ? _ram_T_389[287:0] : _GEN_14504; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15555 = 10'h147 == _T_35 ? _ram_T_389[287:0] : _GEN_14505; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15556 = 10'h148 == _T_35 ? _ram_T_389[287:0] : _GEN_14506; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15557 = 10'h149 == _T_35 ? _ram_T_389[287:0] : _GEN_14507; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15558 = 10'h14a == _T_35 ? _ram_T_389[287:0] : _GEN_14508; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15559 = 10'h14b == _T_35 ? _ram_T_389[287:0] : _GEN_14509; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15560 = 10'h14c == _T_35 ? _ram_T_389[287:0] : _GEN_14510; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15561 = 10'h14d == _T_35 ? _ram_T_389[287:0] : _GEN_14511; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15562 = 10'h14e == _T_35 ? _ram_T_389[287:0] : _GEN_14512; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15563 = 10'h14f == _T_35 ? _ram_T_389[287:0] : _GEN_14513; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15564 = 10'h150 == _T_35 ? _ram_T_389[287:0] : _GEN_14514; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15565 = 10'h151 == _T_35 ? _ram_T_389[287:0] : _GEN_14515; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15566 = 10'h152 == _T_35 ? _ram_T_389[287:0] : _GEN_14516; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15567 = 10'h153 == _T_35 ? _ram_T_389[287:0] : _GEN_14517; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15568 = 10'h154 == _T_35 ? _ram_T_389[287:0] : _GEN_14518; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15569 = 10'h155 == _T_35 ? _ram_T_389[287:0] : _GEN_14519; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15570 = 10'h156 == _T_35 ? _ram_T_389[287:0] : _GEN_14520; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15571 = 10'h157 == _T_35 ? _ram_T_389[287:0] : _GEN_14521; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15572 = 10'h158 == _T_35 ? _ram_T_389[287:0] : _GEN_14522; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15573 = 10'h159 == _T_35 ? _ram_T_389[287:0] : _GEN_14523; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15574 = 10'h15a == _T_35 ? _ram_T_389[287:0] : _GEN_14524; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15575 = 10'h15b == _T_35 ? _ram_T_389[287:0] : _GEN_14525; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15576 = 10'h15c == _T_35 ? _ram_T_389[287:0] : _GEN_14526; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15577 = 10'h15d == _T_35 ? _ram_T_389[287:0] : _GEN_14527; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15578 = 10'h15e == _T_35 ? _ram_T_389[287:0] : _GEN_14528; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15579 = 10'h15f == _T_35 ? _ram_T_389[287:0] : _GEN_14529; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15580 = 10'h160 == _T_35 ? _ram_T_389[287:0] : _GEN_14530; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15581 = 10'h161 == _T_35 ? _ram_T_389[287:0] : _GEN_14531; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15582 = 10'h162 == _T_35 ? _ram_T_389[287:0] : _GEN_14532; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15583 = 10'h163 == _T_35 ? _ram_T_389[287:0] : _GEN_14533; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15584 = 10'h164 == _T_35 ? _ram_T_389[287:0] : _GEN_14534; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15585 = 10'h165 == _T_35 ? _ram_T_389[287:0] : _GEN_14535; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15586 = 10'h166 == _T_35 ? _ram_T_389[287:0] : _GEN_14536; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15587 = 10'h167 == _T_35 ? _ram_T_389[287:0] : _GEN_14537; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15588 = 10'h168 == _T_35 ? _ram_T_389[287:0] : _GEN_14538; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15589 = 10'h169 == _T_35 ? _ram_T_389[287:0] : _GEN_14539; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15590 = 10'h16a == _T_35 ? _ram_T_389[287:0] : _GEN_14540; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15591 = 10'h16b == _T_35 ? _ram_T_389[287:0] : _GEN_14541; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15592 = 10'h16c == _T_35 ? _ram_T_389[287:0] : _GEN_14542; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15593 = 10'h16d == _T_35 ? _ram_T_389[287:0] : _GEN_14543; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15594 = 10'h16e == _T_35 ? _ram_T_389[287:0] : _GEN_14544; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15595 = 10'h16f == _T_35 ? _ram_T_389[287:0] : _GEN_14545; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15596 = 10'h170 == _T_35 ? _ram_T_389[287:0] : _GEN_14546; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15597 = 10'h171 == _T_35 ? _ram_T_389[287:0] : _GEN_14547; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15598 = 10'h172 == _T_35 ? _ram_T_389[287:0] : _GEN_14548; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15599 = 10'h173 == _T_35 ? _ram_T_389[287:0] : _GEN_14549; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15600 = 10'h174 == _T_35 ? _ram_T_389[287:0] : _GEN_14550; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15601 = 10'h175 == _T_35 ? _ram_T_389[287:0] : _GEN_14551; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15602 = 10'h176 == _T_35 ? _ram_T_389[287:0] : _GEN_14552; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15603 = 10'h177 == _T_35 ? _ram_T_389[287:0] : _GEN_14553; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15604 = 10'h178 == _T_35 ? _ram_T_389[287:0] : _GEN_14554; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15605 = 10'h179 == _T_35 ? _ram_T_389[287:0] : _GEN_14555; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15606 = 10'h17a == _T_35 ? _ram_T_389[287:0] : _GEN_14556; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15607 = 10'h17b == _T_35 ? _ram_T_389[287:0] : _GEN_14557; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15608 = 10'h17c == _T_35 ? _ram_T_389[287:0] : _GEN_14558; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15609 = 10'h17d == _T_35 ? _ram_T_389[287:0] : _GEN_14559; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15610 = 10'h17e == _T_35 ? _ram_T_389[287:0] : _GEN_14560; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15611 = 10'h17f == _T_35 ? _ram_T_389[287:0] : _GEN_14561; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15612 = 10'h180 == _T_35 ? _ram_T_389[287:0] : _GEN_14562; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15613 = 10'h181 == _T_35 ? _ram_T_389[287:0] : _GEN_14563; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15614 = 10'h182 == _T_35 ? _ram_T_389[287:0] : _GEN_14564; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15615 = 10'h183 == _T_35 ? _ram_T_389[287:0] : _GEN_14565; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15616 = 10'h184 == _T_35 ? _ram_T_389[287:0] : _GEN_14566; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15617 = 10'h185 == _T_35 ? _ram_T_389[287:0] : _GEN_14567; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15618 = 10'h186 == _T_35 ? _ram_T_389[287:0] : _GEN_14568; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15619 = 10'h187 == _T_35 ? _ram_T_389[287:0] : _GEN_14569; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15620 = 10'h188 == _T_35 ? _ram_T_389[287:0] : _GEN_14570; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15621 = 10'h189 == _T_35 ? _ram_T_389[287:0] : _GEN_14571; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15622 = 10'h18a == _T_35 ? _ram_T_389[287:0] : _GEN_14572; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15623 = 10'h18b == _T_35 ? _ram_T_389[287:0] : _GEN_14573; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15624 = 10'h18c == _T_35 ? _ram_T_389[287:0] : _GEN_14574; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15625 = 10'h18d == _T_35 ? _ram_T_389[287:0] : _GEN_14575; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15626 = 10'h18e == _T_35 ? _ram_T_389[287:0] : _GEN_14576; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15627 = 10'h18f == _T_35 ? _ram_T_389[287:0] : _GEN_14577; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15628 = 10'h190 == _T_35 ? _ram_T_389[287:0] : _GEN_14578; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15629 = 10'h191 == _T_35 ? _ram_T_389[287:0] : _GEN_14579; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15630 = 10'h192 == _T_35 ? _ram_T_389[287:0] : _GEN_14580; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15631 = 10'h193 == _T_35 ? _ram_T_389[287:0] : _GEN_14581; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15632 = 10'h194 == _T_35 ? _ram_T_389[287:0] : _GEN_14582; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15633 = 10'h195 == _T_35 ? _ram_T_389[287:0] : _GEN_14583; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15634 = 10'h196 == _T_35 ? _ram_T_389[287:0] : _GEN_14584; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15635 = 10'h197 == _T_35 ? _ram_T_389[287:0] : _GEN_14585; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15636 = 10'h198 == _T_35 ? _ram_T_389[287:0] : _GEN_14586; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15637 = 10'h199 == _T_35 ? _ram_T_389[287:0] : _GEN_14587; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15638 = 10'h19a == _T_35 ? _ram_T_389[287:0] : _GEN_14588; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15639 = 10'h19b == _T_35 ? _ram_T_389[287:0] : _GEN_14589; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15640 = 10'h19c == _T_35 ? _ram_T_389[287:0] : _GEN_14590; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15641 = 10'h19d == _T_35 ? _ram_T_389[287:0] : _GEN_14591; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15642 = 10'h19e == _T_35 ? _ram_T_389[287:0] : _GEN_14592; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15643 = 10'h19f == _T_35 ? _ram_T_389[287:0] : _GEN_14593; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15644 = 10'h1a0 == _T_35 ? _ram_T_389[287:0] : _GEN_14594; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15645 = 10'h1a1 == _T_35 ? _ram_T_389[287:0] : _GEN_14595; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15646 = 10'h1a2 == _T_35 ? _ram_T_389[287:0] : _GEN_14596; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15647 = 10'h1a3 == _T_35 ? _ram_T_389[287:0] : _GEN_14597; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15648 = 10'h1a4 == _T_35 ? _ram_T_389[287:0] : _GEN_14598; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15649 = 10'h1a5 == _T_35 ? _ram_T_389[287:0] : _GEN_14599; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15650 = 10'h1a6 == _T_35 ? _ram_T_389[287:0] : _GEN_14600; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15651 = 10'h1a7 == _T_35 ? _ram_T_389[287:0] : _GEN_14601; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15652 = 10'h1a8 == _T_35 ? _ram_T_389[287:0] : _GEN_14602; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15653 = 10'h1a9 == _T_35 ? _ram_T_389[287:0] : _GEN_14603; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15654 = 10'h1aa == _T_35 ? _ram_T_389[287:0] : _GEN_14604; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15655 = 10'h1ab == _T_35 ? _ram_T_389[287:0] : _GEN_14605; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15656 = 10'h1ac == _T_35 ? _ram_T_389[287:0] : _GEN_14606; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15657 = 10'h1ad == _T_35 ? _ram_T_389[287:0] : _GEN_14607; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15658 = 10'h1ae == _T_35 ? _ram_T_389[287:0] : _GEN_14608; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15659 = 10'h1af == _T_35 ? _ram_T_389[287:0] : _GEN_14609; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15660 = 10'h1b0 == _T_35 ? _ram_T_389[287:0] : _GEN_14610; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15661 = 10'h1b1 == _T_35 ? _ram_T_389[287:0] : _GEN_14611; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15662 = 10'h1b2 == _T_35 ? _ram_T_389[287:0] : _GEN_14612; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15663 = 10'h1b3 == _T_35 ? _ram_T_389[287:0] : _GEN_14613; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15664 = 10'h1b4 == _T_35 ? _ram_T_389[287:0] : _GEN_14614; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15665 = 10'h1b5 == _T_35 ? _ram_T_389[287:0] : _GEN_14615; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15666 = 10'h1b6 == _T_35 ? _ram_T_389[287:0] : _GEN_14616; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15667 = 10'h1b7 == _T_35 ? _ram_T_389[287:0] : _GEN_14617; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15668 = 10'h1b8 == _T_35 ? _ram_T_389[287:0] : _GEN_14618; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15669 = 10'h1b9 == _T_35 ? _ram_T_389[287:0] : _GEN_14619; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15670 = 10'h1ba == _T_35 ? _ram_T_389[287:0] : _GEN_14620; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15671 = 10'h1bb == _T_35 ? _ram_T_389[287:0] : _GEN_14621; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15672 = 10'h1bc == _T_35 ? _ram_T_389[287:0] : _GEN_14622; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15673 = 10'h1bd == _T_35 ? _ram_T_389[287:0] : _GEN_14623; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15674 = 10'h1be == _T_35 ? _ram_T_389[287:0] : _GEN_14624; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15675 = 10'h1bf == _T_35 ? _ram_T_389[287:0] : _GEN_14625; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15676 = 10'h1c0 == _T_35 ? _ram_T_389[287:0] : _GEN_14626; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15677 = 10'h1c1 == _T_35 ? _ram_T_389[287:0] : _GEN_14627; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15678 = 10'h1c2 == _T_35 ? _ram_T_389[287:0] : _GEN_14628; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15679 = 10'h1c3 == _T_35 ? _ram_T_389[287:0] : _GEN_14629; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15680 = 10'h1c4 == _T_35 ? _ram_T_389[287:0] : _GEN_14630; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15681 = 10'h1c5 == _T_35 ? _ram_T_389[287:0] : _GEN_14631; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15682 = 10'h1c6 == _T_35 ? _ram_T_389[287:0] : _GEN_14632; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15683 = 10'h1c7 == _T_35 ? _ram_T_389[287:0] : _GEN_14633; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15684 = 10'h1c8 == _T_35 ? _ram_T_389[287:0] : _GEN_14634; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15685 = 10'h1c9 == _T_35 ? _ram_T_389[287:0] : _GEN_14635; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15686 = 10'h1ca == _T_35 ? _ram_T_389[287:0] : _GEN_14636; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15687 = 10'h1cb == _T_35 ? _ram_T_389[287:0] : _GEN_14637; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15688 = 10'h1cc == _T_35 ? _ram_T_389[287:0] : _GEN_14638; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15689 = 10'h1cd == _T_35 ? _ram_T_389[287:0] : _GEN_14639; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15690 = 10'h1ce == _T_35 ? _ram_T_389[287:0] : _GEN_14640; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15691 = 10'h1cf == _T_35 ? _ram_T_389[287:0] : _GEN_14641; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15692 = 10'h1d0 == _T_35 ? _ram_T_389[287:0] : _GEN_14642; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15693 = 10'h1d1 == _T_35 ? _ram_T_389[287:0] : _GEN_14643; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15694 = 10'h1d2 == _T_35 ? _ram_T_389[287:0] : _GEN_14644; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15695 = 10'h1d3 == _T_35 ? _ram_T_389[287:0] : _GEN_14645; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15696 = 10'h1d4 == _T_35 ? _ram_T_389[287:0] : _GEN_14646; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15697 = 10'h1d5 == _T_35 ? _ram_T_389[287:0] : _GEN_14647; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15698 = 10'h1d6 == _T_35 ? _ram_T_389[287:0] : _GEN_14648; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15699 = 10'h1d7 == _T_35 ? _ram_T_389[287:0] : _GEN_14649; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15700 = 10'h1d8 == _T_35 ? _ram_T_389[287:0] : _GEN_14650; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15701 = 10'h1d9 == _T_35 ? _ram_T_389[287:0] : _GEN_14651; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15702 = 10'h1da == _T_35 ? _ram_T_389[287:0] : _GEN_14652; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15703 = 10'h1db == _T_35 ? _ram_T_389[287:0] : _GEN_14653; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15704 = 10'h1dc == _T_35 ? _ram_T_389[287:0] : _GEN_14654; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15705 = 10'h1dd == _T_35 ? _ram_T_389[287:0] : _GEN_14655; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15706 = 10'h1de == _T_35 ? _ram_T_389[287:0] : _GEN_14656; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15707 = 10'h1df == _T_35 ? _ram_T_389[287:0] : _GEN_14657; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15708 = 10'h1e0 == _T_35 ? _ram_T_389[287:0] : _GEN_14658; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15709 = 10'h1e1 == _T_35 ? _ram_T_389[287:0] : _GEN_14659; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15710 = 10'h1e2 == _T_35 ? _ram_T_389[287:0] : _GEN_14660; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15711 = 10'h1e3 == _T_35 ? _ram_T_389[287:0] : _GEN_14661; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15712 = 10'h1e4 == _T_35 ? _ram_T_389[287:0] : _GEN_14662; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15713 = 10'h1e5 == _T_35 ? _ram_T_389[287:0] : _GEN_14663; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15714 = 10'h1e6 == _T_35 ? _ram_T_389[287:0] : _GEN_14664; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15715 = 10'h1e7 == _T_35 ? _ram_T_389[287:0] : _GEN_14665; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15716 = 10'h1e8 == _T_35 ? _ram_T_389[287:0] : _GEN_14666; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15717 = 10'h1e9 == _T_35 ? _ram_T_389[287:0] : _GEN_14667; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15718 = 10'h1ea == _T_35 ? _ram_T_389[287:0] : _GEN_14668; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15719 = 10'h1eb == _T_35 ? _ram_T_389[287:0] : _GEN_14669; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15720 = 10'h1ec == _T_35 ? _ram_T_389[287:0] : _GEN_14670; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15721 = 10'h1ed == _T_35 ? _ram_T_389[287:0] : _GEN_14671; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15722 = 10'h1ee == _T_35 ? _ram_T_389[287:0] : _GEN_14672; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15723 = 10'h1ef == _T_35 ? _ram_T_389[287:0] : _GEN_14673; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15724 = 10'h1f0 == _T_35 ? _ram_T_389[287:0] : _GEN_14674; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15725 = 10'h1f1 == _T_35 ? _ram_T_389[287:0] : _GEN_14675; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15726 = 10'h1f2 == _T_35 ? _ram_T_389[287:0] : _GEN_14676; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15727 = 10'h1f3 == _T_35 ? _ram_T_389[287:0] : _GEN_14677; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15728 = 10'h1f4 == _T_35 ? _ram_T_389[287:0] : _GEN_14678; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15729 = 10'h1f5 == _T_35 ? _ram_T_389[287:0] : _GEN_14679; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15730 = 10'h1f6 == _T_35 ? _ram_T_389[287:0] : _GEN_14680; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15731 = 10'h1f7 == _T_35 ? _ram_T_389[287:0] : _GEN_14681; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15732 = 10'h1f8 == _T_35 ? _ram_T_389[287:0] : _GEN_14682; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15733 = 10'h1f9 == _T_35 ? _ram_T_389[287:0] : _GEN_14683; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15734 = 10'h1fa == _T_35 ? _ram_T_389[287:0] : _GEN_14684; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15735 = 10'h1fb == _T_35 ? _ram_T_389[287:0] : _GEN_14685; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15736 = 10'h1fc == _T_35 ? _ram_T_389[287:0] : _GEN_14686; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15737 = 10'h1fd == _T_35 ? _ram_T_389[287:0] : _GEN_14687; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15738 = 10'h1fe == _T_35 ? _ram_T_389[287:0] : _GEN_14688; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15739 = 10'h1ff == _T_35 ? _ram_T_389[287:0] : _GEN_14689; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15740 = 10'h200 == _T_35 ? _ram_T_389[287:0] : _GEN_14690; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15741 = 10'h201 == _T_35 ? _ram_T_389[287:0] : _GEN_14691; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15742 = 10'h202 == _T_35 ? _ram_T_389[287:0] : _GEN_14692; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15743 = 10'h203 == _T_35 ? _ram_T_389[287:0] : _GEN_14693; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15744 = 10'h204 == _T_35 ? _ram_T_389[287:0] : _GEN_14694; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15745 = 10'h205 == _T_35 ? _ram_T_389[287:0] : _GEN_14695; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15746 = 10'h206 == _T_35 ? _ram_T_389[287:0] : _GEN_14696; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15747 = 10'h207 == _T_35 ? _ram_T_389[287:0] : _GEN_14697; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15748 = 10'h208 == _T_35 ? _ram_T_389[287:0] : _GEN_14698; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15749 = 10'h209 == _T_35 ? _ram_T_389[287:0] : _GEN_14699; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15750 = 10'h20a == _T_35 ? _ram_T_389[287:0] : _GEN_14700; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15751 = 10'h20b == _T_35 ? _ram_T_389[287:0] : _GEN_14701; // @[vga.scala 64:24 vga.scala 64:24]
  wire [287:0] _GEN_15752 = 10'h20c == _T_35 ? _ram_T_389[287:0] : _GEN_14702; // @[vga.scala 64:24 vga.scala 64:24]
  wire [9:0] _T_37 = h + 10'hf; // @[vga.scala 64:14]
  wire  ram_hi_hi_hi_lo_15 = vga_mem_ram_MPORT_135_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_15 = vga_mem_ram_MPORT_136_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_15 = vga_mem_ram_MPORT_137_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_15 = vga_mem_ram_MPORT_138_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_15 = vga_mem_ram_MPORT_139_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_15 = vga_mem_ram_MPORT_140_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_15 = vga_mem_ram_MPORT_141_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_15 = vga_mem_ram_MPORT_142_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_15 = vga_mem_ram_MPORT_143_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_410 = {278'h0,ram_hi_hi_hi_lo_15,ram_hi_hi_lo_15,ram_hi_lo_hi_15,ram_hi_lo_lo_15,
    ram_lo_hi_hi_hi_15,ram_lo_hi_hi_lo_15,ram_lo_hi_lo_15,ram_lo_lo_hi_15,ram_lo_lo_lo_15}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19090 = {{8191'd0}, _ram_T_410}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_414 = _GEN_19090 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_15754 = 10'h1 == _T_37 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15755 = 10'h2 == _T_37 ? ram_2 : _GEN_15754; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15756 = 10'h3 == _T_37 ? ram_3 : _GEN_15755; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15757 = 10'h4 == _T_37 ? ram_4 : _GEN_15756; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15758 = 10'h5 == _T_37 ? ram_5 : _GEN_15757; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15759 = 10'h6 == _T_37 ? ram_6 : _GEN_15758; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15760 = 10'h7 == _T_37 ? ram_7 : _GEN_15759; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15761 = 10'h8 == _T_37 ? ram_8 : _GEN_15760; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15762 = 10'h9 == _T_37 ? ram_9 : _GEN_15761; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15763 = 10'ha == _T_37 ? ram_10 : _GEN_15762; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15764 = 10'hb == _T_37 ? ram_11 : _GEN_15763; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15765 = 10'hc == _T_37 ? ram_12 : _GEN_15764; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15766 = 10'hd == _T_37 ? ram_13 : _GEN_15765; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15767 = 10'he == _T_37 ? ram_14 : _GEN_15766; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15768 = 10'hf == _T_37 ? ram_15 : _GEN_15767; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15769 = 10'h10 == _T_37 ? ram_16 : _GEN_15768; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15770 = 10'h11 == _T_37 ? ram_17 : _GEN_15769; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15771 = 10'h12 == _T_37 ? ram_18 : _GEN_15770; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15772 = 10'h13 == _T_37 ? ram_19 : _GEN_15771; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15773 = 10'h14 == _T_37 ? ram_20 : _GEN_15772; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15774 = 10'h15 == _T_37 ? ram_21 : _GEN_15773; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15775 = 10'h16 == _T_37 ? ram_22 : _GEN_15774; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15776 = 10'h17 == _T_37 ? ram_23 : _GEN_15775; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15777 = 10'h18 == _T_37 ? ram_24 : _GEN_15776; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15778 = 10'h19 == _T_37 ? ram_25 : _GEN_15777; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15779 = 10'h1a == _T_37 ? ram_26 : _GEN_15778; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15780 = 10'h1b == _T_37 ? ram_27 : _GEN_15779; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15781 = 10'h1c == _T_37 ? ram_28 : _GEN_15780; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15782 = 10'h1d == _T_37 ? ram_29 : _GEN_15781; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15783 = 10'h1e == _T_37 ? ram_30 : _GEN_15782; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15784 = 10'h1f == _T_37 ? ram_31 : _GEN_15783; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15785 = 10'h20 == _T_37 ? ram_32 : _GEN_15784; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15786 = 10'h21 == _T_37 ? ram_33 : _GEN_15785; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15787 = 10'h22 == _T_37 ? ram_34 : _GEN_15786; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15788 = 10'h23 == _T_37 ? ram_35 : _GEN_15787; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15789 = 10'h24 == _T_37 ? ram_36 : _GEN_15788; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15790 = 10'h25 == _T_37 ? ram_37 : _GEN_15789; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15791 = 10'h26 == _T_37 ? ram_38 : _GEN_15790; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15792 = 10'h27 == _T_37 ? ram_39 : _GEN_15791; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15793 = 10'h28 == _T_37 ? ram_40 : _GEN_15792; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15794 = 10'h29 == _T_37 ? ram_41 : _GEN_15793; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15795 = 10'h2a == _T_37 ? ram_42 : _GEN_15794; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15796 = 10'h2b == _T_37 ? ram_43 : _GEN_15795; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15797 = 10'h2c == _T_37 ? ram_44 : _GEN_15796; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15798 = 10'h2d == _T_37 ? ram_45 : _GEN_15797; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15799 = 10'h2e == _T_37 ? ram_46 : _GEN_15798; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15800 = 10'h2f == _T_37 ? ram_47 : _GEN_15799; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15801 = 10'h30 == _T_37 ? ram_48 : _GEN_15800; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15802 = 10'h31 == _T_37 ? ram_49 : _GEN_15801; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15803 = 10'h32 == _T_37 ? ram_50 : _GEN_15802; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15804 = 10'h33 == _T_37 ? ram_51 : _GEN_15803; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15805 = 10'h34 == _T_37 ? ram_52 : _GEN_15804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15806 = 10'h35 == _T_37 ? ram_53 : _GEN_15805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15807 = 10'h36 == _T_37 ? ram_54 : _GEN_15806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15808 = 10'h37 == _T_37 ? ram_55 : _GEN_15807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15809 = 10'h38 == _T_37 ? ram_56 : _GEN_15808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15810 = 10'h39 == _T_37 ? ram_57 : _GEN_15809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15811 = 10'h3a == _T_37 ? ram_58 : _GEN_15810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15812 = 10'h3b == _T_37 ? ram_59 : _GEN_15811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15813 = 10'h3c == _T_37 ? ram_60 : _GEN_15812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15814 = 10'h3d == _T_37 ? ram_61 : _GEN_15813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15815 = 10'h3e == _T_37 ? ram_62 : _GEN_15814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15816 = 10'h3f == _T_37 ? ram_63 : _GEN_15815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15817 = 10'h40 == _T_37 ? ram_64 : _GEN_15816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15818 = 10'h41 == _T_37 ? ram_65 : _GEN_15817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15819 = 10'h42 == _T_37 ? ram_66 : _GEN_15818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15820 = 10'h43 == _T_37 ? ram_67 : _GEN_15819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15821 = 10'h44 == _T_37 ? ram_68 : _GEN_15820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15822 = 10'h45 == _T_37 ? ram_69 : _GEN_15821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15823 = 10'h46 == _T_37 ? ram_70 : _GEN_15822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15824 = 10'h47 == _T_37 ? ram_71 : _GEN_15823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15825 = 10'h48 == _T_37 ? ram_72 : _GEN_15824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15826 = 10'h49 == _T_37 ? ram_73 : _GEN_15825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15827 = 10'h4a == _T_37 ? ram_74 : _GEN_15826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15828 = 10'h4b == _T_37 ? ram_75 : _GEN_15827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15829 = 10'h4c == _T_37 ? ram_76 : _GEN_15828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15830 = 10'h4d == _T_37 ? ram_77 : _GEN_15829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15831 = 10'h4e == _T_37 ? ram_78 : _GEN_15830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15832 = 10'h4f == _T_37 ? ram_79 : _GEN_15831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15833 = 10'h50 == _T_37 ? ram_80 : _GEN_15832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15834 = 10'h51 == _T_37 ? ram_81 : _GEN_15833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15835 = 10'h52 == _T_37 ? ram_82 : _GEN_15834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15836 = 10'h53 == _T_37 ? ram_83 : _GEN_15835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15837 = 10'h54 == _T_37 ? ram_84 : _GEN_15836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15838 = 10'h55 == _T_37 ? ram_85 : _GEN_15837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15839 = 10'h56 == _T_37 ? ram_86 : _GEN_15838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15840 = 10'h57 == _T_37 ? ram_87 : _GEN_15839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15841 = 10'h58 == _T_37 ? ram_88 : _GEN_15840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15842 = 10'h59 == _T_37 ? ram_89 : _GEN_15841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15843 = 10'h5a == _T_37 ? ram_90 : _GEN_15842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15844 = 10'h5b == _T_37 ? ram_91 : _GEN_15843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15845 = 10'h5c == _T_37 ? ram_92 : _GEN_15844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15846 = 10'h5d == _T_37 ? ram_93 : _GEN_15845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15847 = 10'h5e == _T_37 ? ram_94 : _GEN_15846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15848 = 10'h5f == _T_37 ? ram_95 : _GEN_15847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15849 = 10'h60 == _T_37 ? ram_96 : _GEN_15848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15850 = 10'h61 == _T_37 ? ram_97 : _GEN_15849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15851 = 10'h62 == _T_37 ? ram_98 : _GEN_15850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15852 = 10'h63 == _T_37 ? ram_99 : _GEN_15851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15853 = 10'h64 == _T_37 ? ram_100 : _GEN_15852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15854 = 10'h65 == _T_37 ? ram_101 : _GEN_15853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15855 = 10'h66 == _T_37 ? ram_102 : _GEN_15854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15856 = 10'h67 == _T_37 ? ram_103 : _GEN_15855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15857 = 10'h68 == _T_37 ? ram_104 : _GEN_15856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15858 = 10'h69 == _T_37 ? ram_105 : _GEN_15857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15859 = 10'h6a == _T_37 ? ram_106 : _GEN_15858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15860 = 10'h6b == _T_37 ? ram_107 : _GEN_15859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15861 = 10'h6c == _T_37 ? ram_108 : _GEN_15860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15862 = 10'h6d == _T_37 ? ram_109 : _GEN_15861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15863 = 10'h6e == _T_37 ? ram_110 : _GEN_15862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15864 = 10'h6f == _T_37 ? ram_111 : _GEN_15863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15865 = 10'h70 == _T_37 ? ram_112 : _GEN_15864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15866 = 10'h71 == _T_37 ? ram_113 : _GEN_15865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15867 = 10'h72 == _T_37 ? ram_114 : _GEN_15866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15868 = 10'h73 == _T_37 ? ram_115 : _GEN_15867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15869 = 10'h74 == _T_37 ? ram_116 : _GEN_15868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15870 = 10'h75 == _T_37 ? ram_117 : _GEN_15869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15871 = 10'h76 == _T_37 ? ram_118 : _GEN_15870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15872 = 10'h77 == _T_37 ? ram_119 : _GEN_15871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15873 = 10'h78 == _T_37 ? ram_120 : _GEN_15872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15874 = 10'h79 == _T_37 ? ram_121 : _GEN_15873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15875 = 10'h7a == _T_37 ? ram_122 : _GEN_15874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15876 = 10'h7b == _T_37 ? ram_123 : _GEN_15875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15877 = 10'h7c == _T_37 ? ram_124 : _GEN_15876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15878 = 10'h7d == _T_37 ? ram_125 : _GEN_15877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15879 = 10'h7e == _T_37 ? ram_126 : _GEN_15878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15880 = 10'h7f == _T_37 ? ram_127 : _GEN_15879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15881 = 10'h80 == _T_37 ? ram_128 : _GEN_15880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15882 = 10'h81 == _T_37 ? ram_129 : _GEN_15881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15883 = 10'h82 == _T_37 ? ram_130 : _GEN_15882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15884 = 10'h83 == _T_37 ? ram_131 : _GEN_15883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15885 = 10'h84 == _T_37 ? ram_132 : _GEN_15884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15886 = 10'h85 == _T_37 ? ram_133 : _GEN_15885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15887 = 10'h86 == _T_37 ? ram_134 : _GEN_15886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15888 = 10'h87 == _T_37 ? ram_135 : _GEN_15887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15889 = 10'h88 == _T_37 ? ram_136 : _GEN_15888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15890 = 10'h89 == _T_37 ? ram_137 : _GEN_15889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15891 = 10'h8a == _T_37 ? ram_138 : _GEN_15890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15892 = 10'h8b == _T_37 ? ram_139 : _GEN_15891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15893 = 10'h8c == _T_37 ? ram_140 : _GEN_15892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15894 = 10'h8d == _T_37 ? ram_141 : _GEN_15893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15895 = 10'h8e == _T_37 ? ram_142 : _GEN_15894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15896 = 10'h8f == _T_37 ? ram_143 : _GEN_15895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15897 = 10'h90 == _T_37 ? ram_144 : _GEN_15896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15898 = 10'h91 == _T_37 ? ram_145 : _GEN_15897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15899 = 10'h92 == _T_37 ? ram_146 : _GEN_15898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15900 = 10'h93 == _T_37 ? ram_147 : _GEN_15899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15901 = 10'h94 == _T_37 ? ram_148 : _GEN_15900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15902 = 10'h95 == _T_37 ? ram_149 : _GEN_15901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15903 = 10'h96 == _T_37 ? ram_150 : _GEN_15902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15904 = 10'h97 == _T_37 ? ram_151 : _GEN_15903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15905 = 10'h98 == _T_37 ? ram_152 : _GEN_15904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15906 = 10'h99 == _T_37 ? ram_153 : _GEN_15905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15907 = 10'h9a == _T_37 ? ram_154 : _GEN_15906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15908 = 10'h9b == _T_37 ? ram_155 : _GEN_15907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15909 = 10'h9c == _T_37 ? ram_156 : _GEN_15908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15910 = 10'h9d == _T_37 ? ram_157 : _GEN_15909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15911 = 10'h9e == _T_37 ? ram_158 : _GEN_15910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15912 = 10'h9f == _T_37 ? ram_159 : _GEN_15911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15913 = 10'ha0 == _T_37 ? ram_160 : _GEN_15912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15914 = 10'ha1 == _T_37 ? ram_161 : _GEN_15913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15915 = 10'ha2 == _T_37 ? ram_162 : _GEN_15914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15916 = 10'ha3 == _T_37 ? ram_163 : _GEN_15915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15917 = 10'ha4 == _T_37 ? ram_164 : _GEN_15916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15918 = 10'ha5 == _T_37 ? ram_165 : _GEN_15917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15919 = 10'ha6 == _T_37 ? ram_166 : _GEN_15918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15920 = 10'ha7 == _T_37 ? ram_167 : _GEN_15919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15921 = 10'ha8 == _T_37 ? ram_168 : _GEN_15920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15922 = 10'ha9 == _T_37 ? ram_169 : _GEN_15921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15923 = 10'haa == _T_37 ? ram_170 : _GEN_15922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15924 = 10'hab == _T_37 ? ram_171 : _GEN_15923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15925 = 10'hac == _T_37 ? ram_172 : _GEN_15924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15926 = 10'had == _T_37 ? ram_173 : _GEN_15925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15927 = 10'hae == _T_37 ? ram_174 : _GEN_15926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15928 = 10'haf == _T_37 ? ram_175 : _GEN_15927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15929 = 10'hb0 == _T_37 ? ram_176 : _GEN_15928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15930 = 10'hb1 == _T_37 ? ram_177 : _GEN_15929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15931 = 10'hb2 == _T_37 ? ram_178 : _GEN_15930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15932 = 10'hb3 == _T_37 ? ram_179 : _GEN_15931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15933 = 10'hb4 == _T_37 ? ram_180 : _GEN_15932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15934 = 10'hb5 == _T_37 ? ram_181 : _GEN_15933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15935 = 10'hb6 == _T_37 ? ram_182 : _GEN_15934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15936 = 10'hb7 == _T_37 ? ram_183 : _GEN_15935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15937 = 10'hb8 == _T_37 ? ram_184 : _GEN_15936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15938 = 10'hb9 == _T_37 ? ram_185 : _GEN_15937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15939 = 10'hba == _T_37 ? ram_186 : _GEN_15938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15940 = 10'hbb == _T_37 ? ram_187 : _GEN_15939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15941 = 10'hbc == _T_37 ? ram_188 : _GEN_15940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15942 = 10'hbd == _T_37 ? ram_189 : _GEN_15941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15943 = 10'hbe == _T_37 ? ram_190 : _GEN_15942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15944 = 10'hbf == _T_37 ? ram_191 : _GEN_15943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15945 = 10'hc0 == _T_37 ? ram_192 : _GEN_15944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15946 = 10'hc1 == _T_37 ? ram_193 : _GEN_15945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15947 = 10'hc2 == _T_37 ? ram_194 : _GEN_15946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15948 = 10'hc3 == _T_37 ? ram_195 : _GEN_15947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15949 = 10'hc4 == _T_37 ? ram_196 : _GEN_15948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15950 = 10'hc5 == _T_37 ? ram_197 : _GEN_15949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15951 = 10'hc6 == _T_37 ? ram_198 : _GEN_15950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15952 = 10'hc7 == _T_37 ? ram_199 : _GEN_15951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15953 = 10'hc8 == _T_37 ? ram_200 : _GEN_15952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15954 = 10'hc9 == _T_37 ? ram_201 : _GEN_15953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15955 = 10'hca == _T_37 ? ram_202 : _GEN_15954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15956 = 10'hcb == _T_37 ? ram_203 : _GEN_15955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15957 = 10'hcc == _T_37 ? ram_204 : _GEN_15956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15958 = 10'hcd == _T_37 ? ram_205 : _GEN_15957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15959 = 10'hce == _T_37 ? ram_206 : _GEN_15958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15960 = 10'hcf == _T_37 ? ram_207 : _GEN_15959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15961 = 10'hd0 == _T_37 ? ram_208 : _GEN_15960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15962 = 10'hd1 == _T_37 ? ram_209 : _GEN_15961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15963 = 10'hd2 == _T_37 ? ram_210 : _GEN_15962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15964 = 10'hd3 == _T_37 ? ram_211 : _GEN_15963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15965 = 10'hd4 == _T_37 ? ram_212 : _GEN_15964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15966 = 10'hd5 == _T_37 ? ram_213 : _GEN_15965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15967 = 10'hd6 == _T_37 ? ram_214 : _GEN_15966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15968 = 10'hd7 == _T_37 ? ram_215 : _GEN_15967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15969 = 10'hd8 == _T_37 ? ram_216 : _GEN_15968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15970 = 10'hd9 == _T_37 ? ram_217 : _GEN_15969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15971 = 10'hda == _T_37 ? ram_218 : _GEN_15970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15972 = 10'hdb == _T_37 ? ram_219 : _GEN_15971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15973 = 10'hdc == _T_37 ? ram_220 : _GEN_15972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15974 = 10'hdd == _T_37 ? ram_221 : _GEN_15973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15975 = 10'hde == _T_37 ? ram_222 : _GEN_15974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15976 = 10'hdf == _T_37 ? ram_223 : _GEN_15975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15977 = 10'he0 == _T_37 ? ram_224 : _GEN_15976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15978 = 10'he1 == _T_37 ? ram_225 : _GEN_15977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15979 = 10'he2 == _T_37 ? ram_226 : _GEN_15978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15980 = 10'he3 == _T_37 ? ram_227 : _GEN_15979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15981 = 10'he4 == _T_37 ? ram_228 : _GEN_15980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15982 = 10'he5 == _T_37 ? ram_229 : _GEN_15981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15983 = 10'he6 == _T_37 ? ram_230 : _GEN_15982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15984 = 10'he7 == _T_37 ? ram_231 : _GEN_15983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15985 = 10'he8 == _T_37 ? ram_232 : _GEN_15984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15986 = 10'he9 == _T_37 ? ram_233 : _GEN_15985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15987 = 10'hea == _T_37 ? ram_234 : _GEN_15986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15988 = 10'heb == _T_37 ? ram_235 : _GEN_15987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15989 = 10'hec == _T_37 ? ram_236 : _GEN_15988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15990 = 10'hed == _T_37 ? ram_237 : _GEN_15989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15991 = 10'hee == _T_37 ? ram_238 : _GEN_15990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15992 = 10'hef == _T_37 ? ram_239 : _GEN_15991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15993 = 10'hf0 == _T_37 ? ram_240 : _GEN_15992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15994 = 10'hf1 == _T_37 ? ram_241 : _GEN_15993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15995 = 10'hf2 == _T_37 ? ram_242 : _GEN_15994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15996 = 10'hf3 == _T_37 ? ram_243 : _GEN_15995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15997 = 10'hf4 == _T_37 ? ram_244 : _GEN_15996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15998 = 10'hf5 == _T_37 ? ram_245 : _GEN_15997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_15999 = 10'hf6 == _T_37 ? ram_246 : _GEN_15998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16000 = 10'hf7 == _T_37 ? ram_247 : _GEN_15999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16001 = 10'hf8 == _T_37 ? ram_248 : _GEN_16000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16002 = 10'hf9 == _T_37 ? ram_249 : _GEN_16001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16003 = 10'hfa == _T_37 ? ram_250 : _GEN_16002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16004 = 10'hfb == _T_37 ? ram_251 : _GEN_16003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16005 = 10'hfc == _T_37 ? ram_252 : _GEN_16004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16006 = 10'hfd == _T_37 ? ram_253 : _GEN_16005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16007 = 10'hfe == _T_37 ? ram_254 : _GEN_16006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16008 = 10'hff == _T_37 ? ram_255 : _GEN_16007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16009 = 10'h100 == _T_37 ? ram_256 : _GEN_16008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16010 = 10'h101 == _T_37 ? ram_257 : _GEN_16009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16011 = 10'h102 == _T_37 ? ram_258 : _GEN_16010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16012 = 10'h103 == _T_37 ? ram_259 : _GEN_16011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16013 = 10'h104 == _T_37 ? ram_260 : _GEN_16012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16014 = 10'h105 == _T_37 ? ram_261 : _GEN_16013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16015 = 10'h106 == _T_37 ? ram_262 : _GEN_16014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16016 = 10'h107 == _T_37 ? ram_263 : _GEN_16015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16017 = 10'h108 == _T_37 ? ram_264 : _GEN_16016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16018 = 10'h109 == _T_37 ? ram_265 : _GEN_16017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16019 = 10'h10a == _T_37 ? ram_266 : _GEN_16018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16020 = 10'h10b == _T_37 ? ram_267 : _GEN_16019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16021 = 10'h10c == _T_37 ? ram_268 : _GEN_16020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16022 = 10'h10d == _T_37 ? ram_269 : _GEN_16021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16023 = 10'h10e == _T_37 ? ram_270 : _GEN_16022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16024 = 10'h10f == _T_37 ? ram_271 : _GEN_16023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16025 = 10'h110 == _T_37 ? ram_272 : _GEN_16024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16026 = 10'h111 == _T_37 ? ram_273 : _GEN_16025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16027 = 10'h112 == _T_37 ? ram_274 : _GEN_16026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16028 = 10'h113 == _T_37 ? ram_275 : _GEN_16027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16029 = 10'h114 == _T_37 ? ram_276 : _GEN_16028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16030 = 10'h115 == _T_37 ? ram_277 : _GEN_16029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16031 = 10'h116 == _T_37 ? ram_278 : _GEN_16030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16032 = 10'h117 == _T_37 ? ram_279 : _GEN_16031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16033 = 10'h118 == _T_37 ? ram_280 : _GEN_16032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16034 = 10'h119 == _T_37 ? ram_281 : _GEN_16033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16035 = 10'h11a == _T_37 ? ram_282 : _GEN_16034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16036 = 10'h11b == _T_37 ? ram_283 : _GEN_16035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16037 = 10'h11c == _T_37 ? ram_284 : _GEN_16036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16038 = 10'h11d == _T_37 ? ram_285 : _GEN_16037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16039 = 10'h11e == _T_37 ? ram_286 : _GEN_16038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16040 = 10'h11f == _T_37 ? ram_287 : _GEN_16039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16041 = 10'h120 == _T_37 ? ram_288 : _GEN_16040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16042 = 10'h121 == _T_37 ? ram_289 : _GEN_16041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16043 = 10'h122 == _T_37 ? ram_290 : _GEN_16042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16044 = 10'h123 == _T_37 ? ram_291 : _GEN_16043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16045 = 10'h124 == _T_37 ? ram_292 : _GEN_16044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16046 = 10'h125 == _T_37 ? ram_293 : _GEN_16045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16047 = 10'h126 == _T_37 ? ram_294 : _GEN_16046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16048 = 10'h127 == _T_37 ? ram_295 : _GEN_16047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16049 = 10'h128 == _T_37 ? ram_296 : _GEN_16048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16050 = 10'h129 == _T_37 ? ram_297 : _GEN_16049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16051 = 10'h12a == _T_37 ? ram_298 : _GEN_16050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16052 = 10'h12b == _T_37 ? ram_299 : _GEN_16051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16053 = 10'h12c == _T_37 ? ram_300 : _GEN_16052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16054 = 10'h12d == _T_37 ? ram_301 : _GEN_16053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16055 = 10'h12e == _T_37 ? ram_302 : _GEN_16054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16056 = 10'h12f == _T_37 ? ram_303 : _GEN_16055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16057 = 10'h130 == _T_37 ? ram_304 : _GEN_16056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16058 = 10'h131 == _T_37 ? ram_305 : _GEN_16057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16059 = 10'h132 == _T_37 ? ram_306 : _GEN_16058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16060 = 10'h133 == _T_37 ? ram_307 : _GEN_16059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16061 = 10'h134 == _T_37 ? ram_308 : _GEN_16060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16062 = 10'h135 == _T_37 ? ram_309 : _GEN_16061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16063 = 10'h136 == _T_37 ? ram_310 : _GEN_16062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16064 = 10'h137 == _T_37 ? ram_311 : _GEN_16063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16065 = 10'h138 == _T_37 ? ram_312 : _GEN_16064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16066 = 10'h139 == _T_37 ? ram_313 : _GEN_16065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16067 = 10'h13a == _T_37 ? ram_314 : _GEN_16066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16068 = 10'h13b == _T_37 ? ram_315 : _GEN_16067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16069 = 10'h13c == _T_37 ? ram_316 : _GEN_16068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16070 = 10'h13d == _T_37 ? ram_317 : _GEN_16069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16071 = 10'h13e == _T_37 ? ram_318 : _GEN_16070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16072 = 10'h13f == _T_37 ? ram_319 : _GEN_16071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16073 = 10'h140 == _T_37 ? ram_320 : _GEN_16072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16074 = 10'h141 == _T_37 ? ram_321 : _GEN_16073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16075 = 10'h142 == _T_37 ? ram_322 : _GEN_16074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16076 = 10'h143 == _T_37 ? ram_323 : _GEN_16075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16077 = 10'h144 == _T_37 ? ram_324 : _GEN_16076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16078 = 10'h145 == _T_37 ? ram_325 : _GEN_16077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16079 = 10'h146 == _T_37 ? ram_326 : _GEN_16078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16080 = 10'h147 == _T_37 ? ram_327 : _GEN_16079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16081 = 10'h148 == _T_37 ? ram_328 : _GEN_16080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16082 = 10'h149 == _T_37 ? ram_329 : _GEN_16081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16083 = 10'h14a == _T_37 ? ram_330 : _GEN_16082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16084 = 10'h14b == _T_37 ? ram_331 : _GEN_16083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16085 = 10'h14c == _T_37 ? ram_332 : _GEN_16084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16086 = 10'h14d == _T_37 ? ram_333 : _GEN_16085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16087 = 10'h14e == _T_37 ? ram_334 : _GEN_16086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16088 = 10'h14f == _T_37 ? ram_335 : _GEN_16087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16089 = 10'h150 == _T_37 ? ram_336 : _GEN_16088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16090 = 10'h151 == _T_37 ? ram_337 : _GEN_16089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16091 = 10'h152 == _T_37 ? ram_338 : _GEN_16090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16092 = 10'h153 == _T_37 ? ram_339 : _GEN_16091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16093 = 10'h154 == _T_37 ? ram_340 : _GEN_16092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16094 = 10'h155 == _T_37 ? ram_341 : _GEN_16093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16095 = 10'h156 == _T_37 ? ram_342 : _GEN_16094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16096 = 10'h157 == _T_37 ? ram_343 : _GEN_16095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16097 = 10'h158 == _T_37 ? ram_344 : _GEN_16096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16098 = 10'h159 == _T_37 ? ram_345 : _GEN_16097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16099 = 10'h15a == _T_37 ? ram_346 : _GEN_16098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16100 = 10'h15b == _T_37 ? ram_347 : _GEN_16099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16101 = 10'h15c == _T_37 ? ram_348 : _GEN_16100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16102 = 10'h15d == _T_37 ? ram_349 : _GEN_16101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16103 = 10'h15e == _T_37 ? ram_350 : _GEN_16102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16104 = 10'h15f == _T_37 ? ram_351 : _GEN_16103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16105 = 10'h160 == _T_37 ? ram_352 : _GEN_16104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16106 = 10'h161 == _T_37 ? ram_353 : _GEN_16105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16107 = 10'h162 == _T_37 ? ram_354 : _GEN_16106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16108 = 10'h163 == _T_37 ? ram_355 : _GEN_16107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16109 = 10'h164 == _T_37 ? ram_356 : _GEN_16108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16110 = 10'h165 == _T_37 ? ram_357 : _GEN_16109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16111 = 10'h166 == _T_37 ? ram_358 : _GEN_16110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16112 = 10'h167 == _T_37 ? ram_359 : _GEN_16111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16113 = 10'h168 == _T_37 ? ram_360 : _GEN_16112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16114 = 10'h169 == _T_37 ? ram_361 : _GEN_16113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16115 = 10'h16a == _T_37 ? ram_362 : _GEN_16114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16116 = 10'h16b == _T_37 ? ram_363 : _GEN_16115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16117 = 10'h16c == _T_37 ? ram_364 : _GEN_16116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16118 = 10'h16d == _T_37 ? ram_365 : _GEN_16117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16119 = 10'h16e == _T_37 ? ram_366 : _GEN_16118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16120 = 10'h16f == _T_37 ? ram_367 : _GEN_16119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16121 = 10'h170 == _T_37 ? ram_368 : _GEN_16120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16122 = 10'h171 == _T_37 ? ram_369 : _GEN_16121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16123 = 10'h172 == _T_37 ? ram_370 : _GEN_16122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16124 = 10'h173 == _T_37 ? ram_371 : _GEN_16123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16125 = 10'h174 == _T_37 ? ram_372 : _GEN_16124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16126 = 10'h175 == _T_37 ? ram_373 : _GEN_16125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16127 = 10'h176 == _T_37 ? ram_374 : _GEN_16126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16128 = 10'h177 == _T_37 ? ram_375 : _GEN_16127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16129 = 10'h178 == _T_37 ? ram_376 : _GEN_16128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16130 = 10'h179 == _T_37 ? ram_377 : _GEN_16129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16131 = 10'h17a == _T_37 ? ram_378 : _GEN_16130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16132 = 10'h17b == _T_37 ? ram_379 : _GEN_16131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16133 = 10'h17c == _T_37 ? ram_380 : _GEN_16132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16134 = 10'h17d == _T_37 ? ram_381 : _GEN_16133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16135 = 10'h17e == _T_37 ? ram_382 : _GEN_16134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16136 = 10'h17f == _T_37 ? ram_383 : _GEN_16135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16137 = 10'h180 == _T_37 ? ram_384 : _GEN_16136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16138 = 10'h181 == _T_37 ? ram_385 : _GEN_16137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16139 = 10'h182 == _T_37 ? ram_386 : _GEN_16138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16140 = 10'h183 == _T_37 ? ram_387 : _GEN_16139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16141 = 10'h184 == _T_37 ? ram_388 : _GEN_16140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16142 = 10'h185 == _T_37 ? ram_389 : _GEN_16141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16143 = 10'h186 == _T_37 ? ram_390 : _GEN_16142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16144 = 10'h187 == _T_37 ? ram_391 : _GEN_16143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16145 = 10'h188 == _T_37 ? ram_392 : _GEN_16144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16146 = 10'h189 == _T_37 ? ram_393 : _GEN_16145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16147 = 10'h18a == _T_37 ? ram_394 : _GEN_16146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16148 = 10'h18b == _T_37 ? ram_395 : _GEN_16147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16149 = 10'h18c == _T_37 ? ram_396 : _GEN_16148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16150 = 10'h18d == _T_37 ? ram_397 : _GEN_16149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16151 = 10'h18e == _T_37 ? ram_398 : _GEN_16150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16152 = 10'h18f == _T_37 ? ram_399 : _GEN_16151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16153 = 10'h190 == _T_37 ? ram_400 : _GEN_16152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16154 = 10'h191 == _T_37 ? ram_401 : _GEN_16153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16155 = 10'h192 == _T_37 ? ram_402 : _GEN_16154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16156 = 10'h193 == _T_37 ? ram_403 : _GEN_16155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16157 = 10'h194 == _T_37 ? ram_404 : _GEN_16156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16158 = 10'h195 == _T_37 ? ram_405 : _GEN_16157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16159 = 10'h196 == _T_37 ? ram_406 : _GEN_16158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16160 = 10'h197 == _T_37 ? ram_407 : _GEN_16159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16161 = 10'h198 == _T_37 ? ram_408 : _GEN_16160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16162 = 10'h199 == _T_37 ? ram_409 : _GEN_16161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16163 = 10'h19a == _T_37 ? ram_410 : _GEN_16162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16164 = 10'h19b == _T_37 ? ram_411 : _GEN_16163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16165 = 10'h19c == _T_37 ? ram_412 : _GEN_16164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16166 = 10'h19d == _T_37 ? ram_413 : _GEN_16165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16167 = 10'h19e == _T_37 ? ram_414 : _GEN_16166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16168 = 10'h19f == _T_37 ? ram_415 : _GEN_16167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16169 = 10'h1a0 == _T_37 ? ram_416 : _GEN_16168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16170 = 10'h1a1 == _T_37 ? ram_417 : _GEN_16169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16171 = 10'h1a2 == _T_37 ? ram_418 : _GEN_16170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16172 = 10'h1a3 == _T_37 ? ram_419 : _GEN_16171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16173 = 10'h1a4 == _T_37 ? ram_420 : _GEN_16172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16174 = 10'h1a5 == _T_37 ? ram_421 : _GEN_16173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16175 = 10'h1a6 == _T_37 ? ram_422 : _GEN_16174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16176 = 10'h1a7 == _T_37 ? ram_423 : _GEN_16175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16177 = 10'h1a8 == _T_37 ? ram_424 : _GEN_16176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16178 = 10'h1a9 == _T_37 ? ram_425 : _GEN_16177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16179 = 10'h1aa == _T_37 ? ram_426 : _GEN_16178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16180 = 10'h1ab == _T_37 ? ram_427 : _GEN_16179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16181 = 10'h1ac == _T_37 ? ram_428 : _GEN_16180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16182 = 10'h1ad == _T_37 ? ram_429 : _GEN_16181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16183 = 10'h1ae == _T_37 ? ram_430 : _GEN_16182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16184 = 10'h1af == _T_37 ? ram_431 : _GEN_16183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16185 = 10'h1b0 == _T_37 ? ram_432 : _GEN_16184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16186 = 10'h1b1 == _T_37 ? ram_433 : _GEN_16185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16187 = 10'h1b2 == _T_37 ? ram_434 : _GEN_16186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16188 = 10'h1b3 == _T_37 ? ram_435 : _GEN_16187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16189 = 10'h1b4 == _T_37 ? ram_436 : _GEN_16188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16190 = 10'h1b5 == _T_37 ? ram_437 : _GEN_16189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16191 = 10'h1b6 == _T_37 ? ram_438 : _GEN_16190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16192 = 10'h1b7 == _T_37 ? ram_439 : _GEN_16191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16193 = 10'h1b8 == _T_37 ? ram_440 : _GEN_16192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16194 = 10'h1b9 == _T_37 ? ram_441 : _GEN_16193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16195 = 10'h1ba == _T_37 ? ram_442 : _GEN_16194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16196 = 10'h1bb == _T_37 ? ram_443 : _GEN_16195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16197 = 10'h1bc == _T_37 ? ram_444 : _GEN_16196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16198 = 10'h1bd == _T_37 ? ram_445 : _GEN_16197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16199 = 10'h1be == _T_37 ? ram_446 : _GEN_16198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16200 = 10'h1bf == _T_37 ? ram_447 : _GEN_16199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16201 = 10'h1c0 == _T_37 ? ram_448 : _GEN_16200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16202 = 10'h1c1 == _T_37 ? ram_449 : _GEN_16201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16203 = 10'h1c2 == _T_37 ? ram_450 : _GEN_16202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16204 = 10'h1c3 == _T_37 ? ram_451 : _GEN_16203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16205 = 10'h1c4 == _T_37 ? ram_452 : _GEN_16204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16206 = 10'h1c5 == _T_37 ? ram_453 : _GEN_16205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16207 = 10'h1c6 == _T_37 ? ram_454 : _GEN_16206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16208 = 10'h1c7 == _T_37 ? ram_455 : _GEN_16207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16209 = 10'h1c8 == _T_37 ? ram_456 : _GEN_16208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16210 = 10'h1c9 == _T_37 ? ram_457 : _GEN_16209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16211 = 10'h1ca == _T_37 ? ram_458 : _GEN_16210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16212 = 10'h1cb == _T_37 ? ram_459 : _GEN_16211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16213 = 10'h1cc == _T_37 ? ram_460 : _GEN_16212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16214 = 10'h1cd == _T_37 ? ram_461 : _GEN_16213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16215 = 10'h1ce == _T_37 ? ram_462 : _GEN_16214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16216 = 10'h1cf == _T_37 ? ram_463 : _GEN_16215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16217 = 10'h1d0 == _T_37 ? ram_464 : _GEN_16216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16218 = 10'h1d1 == _T_37 ? ram_465 : _GEN_16217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16219 = 10'h1d2 == _T_37 ? ram_466 : _GEN_16218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16220 = 10'h1d3 == _T_37 ? ram_467 : _GEN_16219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16221 = 10'h1d4 == _T_37 ? ram_468 : _GEN_16220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16222 = 10'h1d5 == _T_37 ? ram_469 : _GEN_16221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16223 = 10'h1d6 == _T_37 ? ram_470 : _GEN_16222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16224 = 10'h1d7 == _T_37 ? ram_471 : _GEN_16223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16225 = 10'h1d8 == _T_37 ? ram_472 : _GEN_16224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16226 = 10'h1d9 == _T_37 ? ram_473 : _GEN_16225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16227 = 10'h1da == _T_37 ? ram_474 : _GEN_16226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16228 = 10'h1db == _T_37 ? ram_475 : _GEN_16227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16229 = 10'h1dc == _T_37 ? ram_476 : _GEN_16228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16230 = 10'h1dd == _T_37 ? ram_477 : _GEN_16229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16231 = 10'h1de == _T_37 ? ram_478 : _GEN_16230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16232 = 10'h1df == _T_37 ? ram_479 : _GEN_16231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16233 = 10'h1e0 == _T_37 ? ram_480 : _GEN_16232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16234 = 10'h1e1 == _T_37 ? ram_481 : _GEN_16233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16235 = 10'h1e2 == _T_37 ? ram_482 : _GEN_16234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16236 = 10'h1e3 == _T_37 ? ram_483 : _GEN_16235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16237 = 10'h1e4 == _T_37 ? ram_484 : _GEN_16236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16238 = 10'h1e5 == _T_37 ? ram_485 : _GEN_16237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16239 = 10'h1e6 == _T_37 ? ram_486 : _GEN_16238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16240 = 10'h1e7 == _T_37 ? ram_487 : _GEN_16239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16241 = 10'h1e8 == _T_37 ? ram_488 : _GEN_16240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16242 = 10'h1e9 == _T_37 ? ram_489 : _GEN_16241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16243 = 10'h1ea == _T_37 ? ram_490 : _GEN_16242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16244 = 10'h1eb == _T_37 ? ram_491 : _GEN_16243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16245 = 10'h1ec == _T_37 ? ram_492 : _GEN_16244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16246 = 10'h1ed == _T_37 ? ram_493 : _GEN_16245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16247 = 10'h1ee == _T_37 ? ram_494 : _GEN_16246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16248 = 10'h1ef == _T_37 ? ram_495 : _GEN_16247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16249 = 10'h1f0 == _T_37 ? ram_496 : _GEN_16248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16250 = 10'h1f1 == _T_37 ? ram_497 : _GEN_16249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16251 = 10'h1f2 == _T_37 ? ram_498 : _GEN_16250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16252 = 10'h1f3 == _T_37 ? ram_499 : _GEN_16251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16253 = 10'h1f4 == _T_37 ? ram_500 : _GEN_16252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16254 = 10'h1f5 == _T_37 ? ram_501 : _GEN_16253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16255 = 10'h1f6 == _T_37 ? ram_502 : _GEN_16254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16256 = 10'h1f7 == _T_37 ? ram_503 : _GEN_16255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16257 = 10'h1f8 == _T_37 ? ram_504 : _GEN_16256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16258 = 10'h1f9 == _T_37 ? ram_505 : _GEN_16257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16259 = 10'h1fa == _T_37 ? ram_506 : _GEN_16258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16260 = 10'h1fb == _T_37 ? ram_507 : _GEN_16259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16261 = 10'h1fc == _T_37 ? ram_508 : _GEN_16260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16262 = 10'h1fd == _T_37 ? ram_509 : _GEN_16261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16263 = 10'h1fe == _T_37 ? ram_510 : _GEN_16262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16264 = 10'h1ff == _T_37 ? ram_511 : _GEN_16263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16265 = 10'h200 == _T_37 ? ram_512 : _GEN_16264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16266 = 10'h201 == _T_37 ? ram_513 : _GEN_16265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16267 = 10'h202 == _T_37 ? ram_514 : _GEN_16266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16268 = 10'h203 == _T_37 ? ram_515 : _GEN_16267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16269 = 10'h204 == _T_37 ? ram_516 : _GEN_16268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16270 = 10'h205 == _T_37 ? ram_517 : _GEN_16269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16271 = 10'h206 == _T_37 ? ram_518 : _GEN_16270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16272 = 10'h207 == _T_37 ? ram_519 : _GEN_16271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16273 = 10'h208 == _T_37 ? ram_520 : _GEN_16272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16274 = 10'h209 == _T_37 ? ram_521 : _GEN_16273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16275 = 10'h20a == _T_37 ? ram_522 : _GEN_16274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16276 = 10'h20b == _T_37 ? ram_523 : _GEN_16275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16277 = 10'h20c == _T_37 ? ram_524 : _GEN_16276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19091 = {{8190'd0}, _GEN_16277}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_415 = _GEN_19091 ^ _ram_T_414; // @[vga.scala 64:41]
  wire  ram_hi_hi_hi_lo_16 = vga_mem_ram_MPORT_144_data[0]; // @[vga.scala 64:83]
  wire  ram_hi_hi_lo_16 = vga_mem_ram_MPORT_145_data[1]; // @[vga.scala 64:109]
  wire  ram_hi_lo_hi_16 = vga_mem_ram_MPORT_146_data[2]; // @[vga.scala 64:135]
  wire  ram_hi_lo_lo_16 = vga_mem_ram_MPORT_147_data[3]; // @[vga.scala 64:161]
  wire  ram_lo_hi_hi_hi_16 = vga_mem_ram_MPORT_148_data[4]; // @[vga.scala 64:187]
  wire  ram_lo_hi_hi_lo_16 = vga_mem_ram_MPORT_149_data[5]; // @[vga.scala 64:213]
  wire  ram_lo_hi_lo_16 = vga_mem_ram_MPORT_150_data[6]; // @[vga.scala 64:239]
  wire  ram_lo_lo_hi_16 = vga_mem_ram_MPORT_151_data[7]; // @[vga.scala 64:265]
  wire  ram_lo_lo_lo_16 = vga_mem_ram_MPORT_152_data[8]; // @[vga.scala 64:291]
  wire [286:0] _ram_T_436 = {278'h0,ram_hi_hi_hi_lo_16,ram_hi_hi_lo_16,ram_hi_lo_hi_16,ram_hi_lo_lo_16,
    ram_lo_hi_hi_hi_16,ram_lo_hi_hi_lo_16,ram_lo_hi_lo_16,ram_lo_lo_hi_16,ram_lo_lo_lo_16}; // @[Cat.scala 30:58]
  wire [8477:0] _GEN_19092 = {{8191'd0}, _ram_T_436}; // @[vga.scala 64:295]
  wire [8477:0] _ram_T_440 = _GEN_19092 << _ram_T_23; // @[vga.scala 64:295]
  wire [287:0] _GEN_16804 = 10'h1 == _h_T_1 ? ram_1 : ram_0; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16805 = 10'h2 == _h_T_1 ? ram_2 : _GEN_16804; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16806 = 10'h3 == _h_T_1 ? ram_3 : _GEN_16805; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16807 = 10'h4 == _h_T_1 ? ram_4 : _GEN_16806; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16808 = 10'h5 == _h_T_1 ? ram_5 : _GEN_16807; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16809 = 10'h6 == _h_T_1 ? ram_6 : _GEN_16808; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16810 = 10'h7 == _h_T_1 ? ram_7 : _GEN_16809; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16811 = 10'h8 == _h_T_1 ? ram_8 : _GEN_16810; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16812 = 10'h9 == _h_T_1 ? ram_9 : _GEN_16811; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16813 = 10'ha == _h_T_1 ? ram_10 : _GEN_16812; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16814 = 10'hb == _h_T_1 ? ram_11 : _GEN_16813; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16815 = 10'hc == _h_T_1 ? ram_12 : _GEN_16814; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16816 = 10'hd == _h_T_1 ? ram_13 : _GEN_16815; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16817 = 10'he == _h_T_1 ? ram_14 : _GEN_16816; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16818 = 10'hf == _h_T_1 ? ram_15 : _GEN_16817; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16819 = 10'h10 == _h_T_1 ? ram_16 : _GEN_16818; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16820 = 10'h11 == _h_T_1 ? ram_17 : _GEN_16819; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16821 = 10'h12 == _h_T_1 ? ram_18 : _GEN_16820; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16822 = 10'h13 == _h_T_1 ? ram_19 : _GEN_16821; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16823 = 10'h14 == _h_T_1 ? ram_20 : _GEN_16822; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16824 = 10'h15 == _h_T_1 ? ram_21 : _GEN_16823; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16825 = 10'h16 == _h_T_1 ? ram_22 : _GEN_16824; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16826 = 10'h17 == _h_T_1 ? ram_23 : _GEN_16825; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16827 = 10'h18 == _h_T_1 ? ram_24 : _GEN_16826; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16828 = 10'h19 == _h_T_1 ? ram_25 : _GEN_16827; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16829 = 10'h1a == _h_T_1 ? ram_26 : _GEN_16828; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16830 = 10'h1b == _h_T_1 ? ram_27 : _GEN_16829; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16831 = 10'h1c == _h_T_1 ? ram_28 : _GEN_16830; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16832 = 10'h1d == _h_T_1 ? ram_29 : _GEN_16831; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16833 = 10'h1e == _h_T_1 ? ram_30 : _GEN_16832; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16834 = 10'h1f == _h_T_1 ? ram_31 : _GEN_16833; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16835 = 10'h20 == _h_T_1 ? ram_32 : _GEN_16834; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16836 = 10'h21 == _h_T_1 ? ram_33 : _GEN_16835; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16837 = 10'h22 == _h_T_1 ? ram_34 : _GEN_16836; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16838 = 10'h23 == _h_T_1 ? ram_35 : _GEN_16837; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16839 = 10'h24 == _h_T_1 ? ram_36 : _GEN_16838; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16840 = 10'h25 == _h_T_1 ? ram_37 : _GEN_16839; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16841 = 10'h26 == _h_T_1 ? ram_38 : _GEN_16840; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16842 = 10'h27 == _h_T_1 ? ram_39 : _GEN_16841; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16843 = 10'h28 == _h_T_1 ? ram_40 : _GEN_16842; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16844 = 10'h29 == _h_T_1 ? ram_41 : _GEN_16843; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16845 = 10'h2a == _h_T_1 ? ram_42 : _GEN_16844; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16846 = 10'h2b == _h_T_1 ? ram_43 : _GEN_16845; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16847 = 10'h2c == _h_T_1 ? ram_44 : _GEN_16846; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16848 = 10'h2d == _h_T_1 ? ram_45 : _GEN_16847; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16849 = 10'h2e == _h_T_1 ? ram_46 : _GEN_16848; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16850 = 10'h2f == _h_T_1 ? ram_47 : _GEN_16849; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16851 = 10'h30 == _h_T_1 ? ram_48 : _GEN_16850; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16852 = 10'h31 == _h_T_1 ? ram_49 : _GEN_16851; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16853 = 10'h32 == _h_T_1 ? ram_50 : _GEN_16852; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16854 = 10'h33 == _h_T_1 ? ram_51 : _GEN_16853; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16855 = 10'h34 == _h_T_1 ? ram_52 : _GEN_16854; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16856 = 10'h35 == _h_T_1 ? ram_53 : _GEN_16855; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16857 = 10'h36 == _h_T_1 ? ram_54 : _GEN_16856; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16858 = 10'h37 == _h_T_1 ? ram_55 : _GEN_16857; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16859 = 10'h38 == _h_T_1 ? ram_56 : _GEN_16858; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16860 = 10'h39 == _h_T_1 ? ram_57 : _GEN_16859; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16861 = 10'h3a == _h_T_1 ? ram_58 : _GEN_16860; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16862 = 10'h3b == _h_T_1 ? ram_59 : _GEN_16861; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16863 = 10'h3c == _h_T_1 ? ram_60 : _GEN_16862; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16864 = 10'h3d == _h_T_1 ? ram_61 : _GEN_16863; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16865 = 10'h3e == _h_T_1 ? ram_62 : _GEN_16864; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16866 = 10'h3f == _h_T_1 ? ram_63 : _GEN_16865; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16867 = 10'h40 == _h_T_1 ? ram_64 : _GEN_16866; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16868 = 10'h41 == _h_T_1 ? ram_65 : _GEN_16867; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16869 = 10'h42 == _h_T_1 ? ram_66 : _GEN_16868; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16870 = 10'h43 == _h_T_1 ? ram_67 : _GEN_16869; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16871 = 10'h44 == _h_T_1 ? ram_68 : _GEN_16870; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16872 = 10'h45 == _h_T_1 ? ram_69 : _GEN_16871; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16873 = 10'h46 == _h_T_1 ? ram_70 : _GEN_16872; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16874 = 10'h47 == _h_T_1 ? ram_71 : _GEN_16873; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16875 = 10'h48 == _h_T_1 ? ram_72 : _GEN_16874; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16876 = 10'h49 == _h_T_1 ? ram_73 : _GEN_16875; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16877 = 10'h4a == _h_T_1 ? ram_74 : _GEN_16876; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16878 = 10'h4b == _h_T_1 ? ram_75 : _GEN_16877; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16879 = 10'h4c == _h_T_1 ? ram_76 : _GEN_16878; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16880 = 10'h4d == _h_T_1 ? ram_77 : _GEN_16879; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16881 = 10'h4e == _h_T_1 ? ram_78 : _GEN_16880; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16882 = 10'h4f == _h_T_1 ? ram_79 : _GEN_16881; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16883 = 10'h50 == _h_T_1 ? ram_80 : _GEN_16882; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16884 = 10'h51 == _h_T_1 ? ram_81 : _GEN_16883; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16885 = 10'h52 == _h_T_1 ? ram_82 : _GEN_16884; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16886 = 10'h53 == _h_T_1 ? ram_83 : _GEN_16885; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16887 = 10'h54 == _h_T_1 ? ram_84 : _GEN_16886; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16888 = 10'h55 == _h_T_1 ? ram_85 : _GEN_16887; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16889 = 10'h56 == _h_T_1 ? ram_86 : _GEN_16888; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16890 = 10'h57 == _h_T_1 ? ram_87 : _GEN_16889; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16891 = 10'h58 == _h_T_1 ? ram_88 : _GEN_16890; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16892 = 10'h59 == _h_T_1 ? ram_89 : _GEN_16891; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16893 = 10'h5a == _h_T_1 ? ram_90 : _GEN_16892; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16894 = 10'h5b == _h_T_1 ? ram_91 : _GEN_16893; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16895 = 10'h5c == _h_T_1 ? ram_92 : _GEN_16894; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16896 = 10'h5d == _h_T_1 ? ram_93 : _GEN_16895; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16897 = 10'h5e == _h_T_1 ? ram_94 : _GEN_16896; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16898 = 10'h5f == _h_T_1 ? ram_95 : _GEN_16897; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16899 = 10'h60 == _h_T_1 ? ram_96 : _GEN_16898; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16900 = 10'h61 == _h_T_1 ? ram_97 : _GEN_16899; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16901 = 10'h62 == _h_T_1 ? ram_98 : _GEN_16900; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16902 = 10'h63 == _h_T_1 ? ram_99 : _GEN_16901; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16903 = 10'h64 == _h_T_1 ? ram_100 : _GEN_16902; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16904 = 10'h65 == _h_T_1 ? ram_101 : _GEN_16903; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16905 = 10'h66 == _h_T_1 ? ram_102 : _GEN_16904; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16906 = 10'h67 == _h_T_1 ? ram_103 : _GEN_16905; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16907 = 10'h68 == _h_T_1 ? ram_104 : _GEN_16906; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16908 = 10'h69 == _h_T_1 ? ram_105 : _GEN_16907; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16909 = 10'h6a == _h_T_1 ? ram_106 : _GEN_16908; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16910 = 10'h6b == _h_T_1 ? ram_107 : _GEN_16909; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16911 = 10'h6c == _h_T_1 ? ram_108 : _GEN_16910; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16912 = 10'h6d == _h_T_1 ? ram_109 : _GEN_16911; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16913 = 10'h6e == _h_T_1 ? ram_110 : _GEN_16912; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16914 = 10'h6f == _h_T_1 ? ram_111 : _GEN_16913; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16915 = 10'h70 == _h_T_1 ? ram_112 : _GEN_16914; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16916 = 10'h71 == _h_T_1 ? ram_113 : _GEN_16915; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16917 = 10'h72 == _h_T_1 ? ram_114 : _GEN_16916; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16918 = 10'h73 == _h_T_1 ? ram_115 : _GEN_16917; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16919 = 10'h74 == _h_T_1 ? ram_116 : _GEN_16918; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16920 = 10'h75 == _h_T_1 ? ram_117 : _GEN_16919; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16921 = 10'h76 == _h_T_1 ? ram_118 : _GEN_16920; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16922 = 10'h77 == _h_T_1 ? ram_119 : _GEN_16921; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16923 = 10'h78 == _h_T_1 ? ram_120 : _GEN_16922; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16924 = 10'h79 == _h_T_1 ? ram_121 : _GEN_16923; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16925 = 10'h7a == _h_T_1 ? ram_122 : _GEN_16924; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16926 = 10'h7b == _h_T_1 ? ram_123 : _GEN_16925; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16927 = 10'h7c == _h_T_1 ? ram_124 : _GEN_16926; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16928 = 10'h7d == _h_T_1 ? ram_125 : _GEN_16927; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16929 = 10'h7e == _h_T_1 ? ram_126 : _GEN_16928; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16930 = 10'h7f == _h_T_1 ? ram_127 : _GEN_16929; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16931 = 10'h80 == _h_T_1 ? ram_128 : _GEN_16930; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16932 = 10'h81 == _h_T_1 ? ram_129 : _GEN_16931; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16933 = 10'h82 == _h_T_1 ? ram_130 : _GEN_16932; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16934 = 10'h83 == _h_T_1 ? ram_131 : _GEN_16933; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16935 = 10'h84 == _h_T_1 ? ram_132 : _GEN_16934; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16936 = 10'h85 == _h_T_1 ? ram_133 : _GEN_16935; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16937 = 10'h86 == _h_T_1 ? ram_134 : _GEN_16936; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16938 = 10'h87 == _h_T_1 ? ram_135 : _GEN_16937; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16939 = 10'h88 == _h_T_1 ? ram_136 : _GEN_16938; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16940 = 10'h89 == _h_T_1 ? ram_137 : _GEN_16939; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16941 = 10'h8a == _h_T_1 ? ram_138 : _GEN_16940; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16942 = 10'h8b == _h_T_1 ? ram_139 : _GEN_16941; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16943 = 10'h8c == _h_T_1 ? ram_140 : _GEN_16942; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16944 = 10'h8d == _h_T_1 ? ram_141 : _GEN_16943; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16945 = 10'h8e == _h_T_1 ? ram_142 : _GEN_16944; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16946 = 10'h8f == _h_T_1 ? ram_143 : _GEN_16945; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16947 = 10'h90 == _h_T_1 ? ram_144 : _GEN_16946; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16948 = 10'h91 == _h_T_1 ? ram_145 : _GEN_16947; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16949 = 10'h92 == _h_T_1 ? ram_146 : _GEN_16948; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16950 = 10'h93 == _h_T_1 ? ram_147 : _GEN_16949; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16951 = 10'h94 == _h_T_1 ? ram_148 : _GEN_16950; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16952 = 10'h95 == _h_T_1 ? ram_149 : _GEN_16951; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16953 = 10'h96 == _h_T_1 ? ram_150 : _GEN_16952; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16954 = 10'h97 == _h_T_1 ? ram_151 : _GEN_16953; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16955 = 10'h98 == _h_T_1 ? ram_152 : _GEN_16954; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16956 = 10'h99 == _h_T_1 ? ram_153 : _GEN_16955; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16957 = 10'h9a == _h_T_1 ? ram_154 : _GEN_16956; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16958 = 10'h9b == _h_T_1 ? ram_155 : _GEN_16957; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16959 = 10'h9c == _h_T_1 ? ram_156 : _GEN_16958; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16960 = 10'h9d == _h_T_1 ? ram_157 : _GEN_16959; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16961 = 10'h9e == _h_T_1 ? ram_158 : _GEN_16960; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16962 = 10'h9f == _h_T_1 ? ram_159 : _GEN_16961; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16963 = 10'ha0 == _h_T_1 ? ram_160 : _GEN_16962; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16964 = 10'ha1 == _h_T_1 ? ram_161 : _GEN_16963; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16965 = 10'ha2 == _h_T_1 ? ram_162 : _GEN_16964; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16966 = 10'ha3 == _h_T_1 ? ram_163 : _GEN_16965; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16967 = 10'ha4 == _h_T_1 ? ram_164 : _GEN_16966; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16968 = 10'ha5 == _h_T_1 ? ram_165 : _GEN_16967; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16969 = 10'ha6 == _h_T_1 ? ram_166 : _GEN_16968; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16970 = 10'ha7 == _h_T_1 ? ram_167 : _GEN_16969; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16971 = 10'ha8 == _h_T_1 ? ram_168 : _GEN_16970; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16972 = 10'ha9 == _h_T_1 ? ram_169 : _GEN_16971; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16973 = 10'haa == _h_T_1 ? ram_170 : _GEN_16972; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16974 = 10'hab == _h_T_1 ? ram_171 : _GEN_16973; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16975 = 10'hac == _h_T_1 ? ram_172 : _GEN_16974; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16976 = 10'had == _h_T_1 ? ram_173 : _GEN_16975; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16977 = 10'hae == _h_T_1 ? ram_174 : _GEN_16976; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16978 = 10'haf == _h_T_1 ? ram_175 : _GEN_16977; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16979 = 10'hb0 == _h_T_1 ? ram_176 : _GEN_16978; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16980 = 10'hb1 == _h_T_1 ? ram_177 : _GEN_16979; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16981 = 10'hb2 == _h_T_1 ? ram_178 : _GEN_16980; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16982 = 10'hb3 == _h_T_1 ? ram_179 : _GEN_16981; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16983 = 10'hb4 == _h_T_1 ? ram_180 : _GEN_16982; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16984 = 10'hb5 == _h_T_1 ? ram_181 : _GEN_16983; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16985 = 10'hb6 == _h_T_1 ? ram_182 : _GEN_16984; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16986 = 10'hb7 == _h_T_1 ? ram_183 : _GEN_16985; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16987 = 10'hb8 == _h_T_1 ? ram_184 : _GEN_16986; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16988 = 10'hb9 == _h_T_1 ? ram_185 : _GEN_16987; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16989 = 10'hba == _h_T_1 ? ram_186 : _GEN_16988; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16990 = 10'hbb == _h_T_1 ? ram_187 : _GEN_16989; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16991 = 10'hbc == _h_T_1 ? ram_188 : _GEN_16990; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16992 = 10'hbd == _h_T_1 ? ram_189 : _GEN_16991; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16993 = 10'hbe == _h_T_1 ? ram_190 : _GEN_16992; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16994 = 10'hbf == _h_T_1 ? ram_191 : _GEN_16993; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16995 = 10'hc0 == _h_T_1 ? ram_192 : _GEN_16994; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16996 = 10'hc1 == _h_T_1 ? ram_193 : _GEN_16995; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16997 = 10'hc2 == _h_T_1 ? ram_194 : _GEN_16996; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16998 = 10'hc3 == _h_T_1 ? ram_195 : _GEN_16997; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_16999 = 10'hc4 == _h_T_1 ? ram_196 : _GEN_16998; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17000 = 10'hc5 == _h_T_1 ? ram_197 : _GEN_16999; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17001 = 10'hc6 == _h_T_1 ? ram_198 : _GEN_17000; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17002 = 10'hc7 == _h_T_1 ? ram_199 : _GEN_17001; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17003 = 10'hc8 == _h_T_1 ? ram_200 : _GEN_17002; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17004 = 10'hc9 == _h_T_1 ? ram_201 : _GEN_17003; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17005 = 10'hca == _h_T_1 ? ram_202 : _GEN_17004; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17006 = 10'hcb == _h_T_1 ? ram_203 : _GEN_17005; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17007 = 10'hcc == _h_T_1 ? ram_204 : _GEN_17006; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17008 = 10'hcd == _h_T_1 ? ram_205 : _GEN_17007; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17009 = 10'hce == _h_T_1 ? ram_206 : _GEN_17008; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17010 = 10'hcf == _h_T_1 ? ram_207 : _GEN_17009; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17011 = 10'hd0 == _h_T_1 ? ram_208 : _GEN_17010; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17012 = 10'hd1 == _h_T_1 ? ram_209 : _GEN_17011; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17013 = 10'hd2 == _h_T_1 ? ram_210 : _GEN_17012; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17014 = 10'hd3 == _h_T_1 ? ram_211 : _GEN_17013; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17015 = 10'hd4 == _h_T_1 ? ram_212 : _GEN_17014; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17016 = 10'hd5 == _h_T_1 ? ram_213 : _GEN_17015; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17017 = 10'hd6 == _h_T_1 ? ram_214 : _GEN_17016; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17018 = 10'hd7 == _h_T_1 ? ram_215 : _GEN_17017; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17019 = 10'hd8 == _h_T_1 ? ram_216 : _GEN_17018; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17020 = 10'hd9 == _h_T_1 ? ram_217 : _GEN_17019; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17021 = 10'hda == _h_T_1 ? ram_218 : _GEN_17020; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17022 = 10'hdb == _h_T_1 ? ram_219 : _GEN_17021; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17023 = 10'hdc == _h_T_1 ? ram_220 : _GEN_17022; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17024 = 10'hdd == _h_T_1 ? ram_221 : _GEN_17023; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17025 = 10'hde == _h_T_1 ? ram_222 : _GEN_17024; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17026 = 10'hdf == _h_T_1 ? ram_223 : _GEN_17025; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17027 = 10'he0 == _h_T_1 ? ram_224 : _GEN_17026; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17028 = 10'he1 == _h_T_1 ? ram_225 : _GEN_17027; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17029 = 10'he2 == _h_T_1 ? ram_226 : _GEN_17028; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17030 = 10'he3 == _h_T_1 ? ram_227 : _GEN_17029; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17031 = 10'he4 == _h_T_1 ? ram_228 : _GEN_17030; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17032 = 10'he5 == _h_T_1 ? ram_229 : _GEN_17031; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17033 = 10'he6 == _h_T_1 ? ram_230 : _GEN_17032; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17034 = 10'he7 == _h_T_1 ? ram_231 : _GEN_17033; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17035 = 10'he8 == _h_T_1 ? ram_232 : _GEN_17034; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17036 = 10'he9 == _h_T_1 ? ram_233 : _GEN_17035; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17037 = 10'hea == _h_T_1 ? ram_234 : _GEN_17036; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17038 = 10'heb == _h_T_1 ? ram_235 : _GEN_17037; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17039 = 10'hec == _h_T_1 ? ram_236 : _GEN_17038; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17040 = 10'hed == _h_T_1 ? ram_237 : _GEN_17039; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17041 = 10'hee == _h_T_1 ? ram_238 : _GEN_17040; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17042 = 10'hef == _h_T_1 ? ram_239 : _GEN_17041; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17043 = 10'hf0 == _h_T_1 ? ram_240 : _GEN_17042; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17044 = 10'hf1 == _h_T_1 ? ram_241 : _GEN_17043; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17045 = 10'hf2 == _h_T_1 ? ram_242 : _GEN_17044; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17046 = 10'hf3 == _h_T_1 ? ram_243 : _GEN_17045; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17047 = 10'hf4 == _h_T_1 ? ram_244 : _GEN_17046; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17048 = 10'hf5 == _h_T_1 ? ram_245 : _GEN_17047; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17049 = 10'hf6 == _h_T_1 ? ram_246 : _GEN_17048; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17050 = 10'hf7 == _h_T_1 ? ram_247 : _GEN_17049; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17051 = 10'hf8 == _h_T_1 ? ram_248 : _GEN_17050; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17052 = 10'hf9 == _h_T_1 ? ram_249 : _GEN_17051; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17053 = 10'hfa == _h_T_1 ? ram_250 : _GEN_17052; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17054 = 10'hfb == _h_T_1 ? ram_251 : _GEN_17053; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17055 = 10'hfc == _h_T_1 ? ram_252 : _GEN_17054; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17056 = 10'hfd == _h_T_1 ? ram_253 : _GEN_17055; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17057 = 10'hfe == _h_T_1 ? ram_254 : _GEN_17056; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17058 = 10'hff == _h_T_1 ? ram_255 : _GEN_17057; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17059 = 10'h100 == _h_T_1 ? ram_256 : _GEN_17058; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17060 = 10'h101 == _h_T_1 ? ram_257 : _GEN_17059; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17061 = 10'h102 == _h_T_1 ? ram_258 : _GEN_17060; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17062 = 10'h103 == _h_T_1 ? ram_259 : _GEN_17061; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17063 = 10'h104 == _h_T_1 ? ram_260 : _GEN_17062; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17064 = 10'h105 == _h_T_1 ? ram_261 : _GEN_17063; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17065 = 10'h106 == _h_T_1 ? ram_262 : _GEN_17064; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17066 = 10'h107 == _h_T_1 ? ram_263 : _GEN_17065; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17067 = 10'h108 == _h_T_1 ? ram_264 : _GEN_17066; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17068 = 10'h109 == _h_T_1 ? ram_265 : _GEN_17067; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17069 = 10'h10a == _h_T_1 ? ram_266 : _GEN_17068; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17070 = 10'h10b == _h_T_1 ? ram_267 : _GEN_17069; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17071 = 10'h10c == _h_T_1 ? ram_268 : _GEN_17070; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17072 = 10'h10d == _h_T_1 ? ram_269 : _GEN_17071; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17073 = 10'h10e == _h_T_1 ? ram_270 : _GEN_17072; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17074 = 10'h10f == _h_T_1 ? ram_271 : _GEN_17073; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17075 = 10'h110 == _h_T_1 ? ram_272 : _GEN_17074; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17076 = 10'h111 == _h_T_1 ? ram_273 : _GEN_17075; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17077 = 10'h112 == _h_T_1 ? ram_274 : _GEN_17076; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17078 = 10'h113 == _h_T_1 ? ram_275 : _GEN_17077; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17079 = 10'h114 == _h_T_1 ? ram_276 : _GEN_17078; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17080 = 10'h115 == _h_T_1 ? ram_277 : _GEN_17079; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17081 = 10'h116 == _h_T_1 ? ram_278 : _GEN_17080; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17082 = 10'h117 == _h_T_1 ? ram_279 : _GEN_17081; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17083 = 10'h118 == _h_T_1 ? ram_280 : _GEN_17082; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17084 = 10'h119 == _h_T_1 ? ram_281 : _GEN_17083; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17085 = 10'h11a == _h_T_1 ? ram_282 : _GEN_17084; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17086 = 10'h11b == _h_T_1 ? ram_283 : _GEN_17085; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17087 = 10'h11c == _h_T_1 ? ram_284 : _GEN_17086; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17088 = 10'h11d == _h_T_1 ? ram_285 : _GEN_17087; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17089 = 10'h11e == _h_T_1 ? ram_286 : _GEN_17088; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17090 = 10'h11f == _h_T_1 ? ram_287 : _GEN_17089; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17091 = 10'h120 == _h_T_1 ? ram_288 : _GEN_17090; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17092 = 10'h121 == _h_T_1 ? ram_289 : _GEN_17091; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17093 = 10'h122 == _h_T_1 ? ram_290 : _GEN_17092; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17094 = 10'h123 == _h_T_1 ? ram_291 : _GEN_17093; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17095 = 10'h124 == _h_T_1 ? ram_292 : _GEN_17094; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17096 = 10'h125 == _h_T_1 ? ram_293 : _GEN_17095; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17097 = 10'h126 == _h_T_1 ? ram_294 : _GEN_17096; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17098 = 10'h127 == _h_T_1 ? ram_295 : _GEN_17097; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17099 = 10'h128 == _h_T_1 ? ram_296 : _GEN_17098; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17100 = 10'h129 == _h_T_1 ? ram_297 : _GEN_17099; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17101 = 10'h12a == _h_T_1 ? ram_298 : _GEN_17100; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17102 = 10'h12b == _h_T_1 ? ram_299 : _GEN_17101; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17103 = 10'h12c == _h_T_1 ? ram_300 : _GEN_17102; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17104 = 10'h12d == _h_T_1 ? ram_301 : _GEN_17103; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17105 = 10'h12e == _h_T_1 ? ram_302 : _GEN_17104; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17106 = 10'h12f == _h_T_1 ? ram_303 : _GEN_17105; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17107 = 10'h130 == _h_T_1 ? ram_304 : _GEN_17106; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17108 = 10'h131 == _h_T_1 ? ram_305 : _GEN_17107; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17109 = 10'h132 == _h_T_1 ? ram_306 : _GEN_17108; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17110 = 10'h133 == _h_T_1 ? ram_307 : _GEN_17109; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17111 = 10'h134 == _h_T_1 ? ram_308 : _GEN_17110; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17112 = 10'h135 == _h_T_1 ? ram_309 : _GEN_17111; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17113 = 10'h136 == _h_T_1 ? ram_310 : _GEN_17112; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17114 = 10'h137 == _h_T_1 ? ram_311 : _GEN_17113; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17115 = 10'h138 == _h_T_1 ? ram_312 : _GEN_17114; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17116 = 10'h139 == _h_T_1 ? ram_313 : _GEN_17115; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17117 = 10'h13a == _h_T_1 ? ram_314 : _GEN_17116; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17118 = 10'h13b == _h_T_1 ? ram_315 : _GEN_17117; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17119 = 10'h13c == _h_T_1 ? ram_316 : _GEN_17118; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17120 = 10'h13d == _h_T_1 ? ram_317 : _GEN_17119; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17121 = 10'h13e == _h_T_1 ? ram_318 : _GEN_17120; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17122 = 10'h13f == _h_T_1 ? ram_319 : _GEN_17121; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17123 = 10'h140 == _h_T_1 ? ram_320 : _GEN_17122; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17124 = 10'h141 == _h_T_1 ? ram_321 : _GEN_17123; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17125 = 10'h142 == _h_T_1 ? ram_322 : _GEN_17124; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17126 = 10'h143 == _h_T_1 ? ram_323 : _GEN_17125; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17127 = 10'h144 == _h_T_1 ? ram_324 : _GEN_17126; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17128 = 10'h145 == _h_T_1 ? ram_325 : _GEN_17127; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17129 = 10'h146 == _h_T_1 ? ram_326 : _GEN_17128; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17130 = 10'h147 == _h_T_1 ? ram_327 : _GEN_17129; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17131 = 10'h148 == _h_T_1 ? ram_328 : _GEN_17130; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17132 = 10'h149 == _h_T_1 ? ram_329 : _GEN_17131; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17133 = 10'h14a == _h_T_1 ? ram_330 : _GEN_17132; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17134 = 10'h14b == _h_T_1 ? ram_331 : _GEN_17133; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17135 = 10'h14c == _h_T_1 ? ram_332 : _GEN_17134; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17136 = 10'h14d == _h_T_1 ? ram_333 : _GEN_17135; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17137 = 10'h14e == _h_T_1 ? ram_334 : _GEN_17136; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17138 = 10'h14f == _h_T_1 ? ram_335 : _GEN_17137; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17139 = 10'h150 == _h_T_1 ? ram_336 : _GEN_17138; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17140 = 10'h151 == _h_T_1 ? ram_337 : _GEN_17139; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17141 = 10'h152 == _h_T_1 ? ram_338 : _GEN_17140; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17142 = 10'h153 == _h_T_1 ? ram_339 : _GEN_17141; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17143 = 10'h154 == _h_T_1 ? ram_340 : _GEN_17142; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17144 = 10'h155 == _h_T_1 ? ram_341 : _GEN_17143; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17145 = 10'h156 == _h_T_1 ? ram_342 : _GEN_17144; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17146 = 10'h157 == _h_T_1 ? ram_343 : _GEN_17145; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17147 = 10'h158 == _h_T_1 ? ram_344 : _GEN_17146; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17148 = 10'h159 == _h_T_1 ? ram_345 : _GEN_17147; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17149 = 10'h15a == _h_T_1 ? ram_346 : _GEN_17148; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17150 = 10'h15b == _h_T_1 ? ram_347 : _GEN_17149; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17151 = 10'h15c == _h_T_1 ? ram_348 : _GEN_17150; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17152 = 10'h15d == _h_T_1 ? ram_349 : _GEN_17151; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17153 = 10'h15e == _h_T_1 ? ram_350 : _GEN_17152; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17154 = 10'h15f == _h_T_1 ? ram_351 : _GEN_17153; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17155 = 10'h160 == _h_T_1 ? ram_352 : _GEN_17154; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17156 = 10'h161 == _h_T_1 ? ram_353 : _GEN_17155; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17157 = 10'h162 == _h_T_1 ? ram_354 : _GEN_17156; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17158 = 10'h163 == _h_T_1 ? ram_355 : _GEN_17157; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17159 = 10'h164 == _h_T_1 ? ram_356 : _GEN_17158; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17160 = 10'h165 == _h_T_1 ? ram_357 : _GEN_17159; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17161 = 10'h166 == _h_T_1 ? ram_358 : _GEN_17160; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17162 = 10'h167 == _h_T_1 ? ram_359 : _GEN_17161; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17163 = 10'h168 == _h_T_1 ? ram_360 : _GEN_17162; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17164 = 10'h169 == _h_T_1 ? ram_361 : _GEN_17163; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17165 = 10'h16a == _h_T_1 ? ram_362 : _GEN_17164; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17166 = 10'h16b == _h_T_1 ? ram_363 : _GEN_17165; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17167 = 10'h16c == _h_T_1 ? ram_364 : _GEN_17166; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17168 = 10'h16d == _h_T_1 ? ram_365 : _GEN_17167; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17169 = 10'h16e == _h_T_1 ? ram_366 : _GEN_17168; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17170 = 10'h16f == _h_T_1 ? ram_367 : _GEN_17169; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17171 = 10'h170 == _h_T_1 ? ram_368 : _GEN_17170; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17172 = 10'h171 == _h_T_1 ? ram_369 : _GEN_17171; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17173 = 10'h172 == _h_T_1 ? ram_370 : _GEN_17172; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17174 = 10'h173 == _h_T_1 ? ram_371 : _GEN_17173; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17175 = 10'h174 == _h_T_1 ? ram_372 : _GEN_17174; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17176 = 10'h175 == _h_T_1 ? ram_373 : _GEN_17175; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17177 = 10'h176 == _h_T_1 ? ram_374 : _GEN_17176; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17178 = 10'h177 == _h_T_1 ? ram_375 : _GEN_17177; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17179 = 10'h178 == _h_T_1 ? ram_376 : _GEN_17178; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17180 = 10'h179 == _h_T_1 ? ram_377 : _GEN_17179; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17181 = 10'h17a == _h_T_1 ? ram_378 : _GEN_17180; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17182 = 10'h17b == _h_T_1 ? ram_379 : _GEN_17181; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17183 = 10'h17c == _h_T_1 ? ram_380 : _GEN_17182; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17184 = 10'h17d == _h_T_1 ? ram_381 : _GEN_17183; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17185 = 10'h17e == _h_T_1 ? ram_382 : _GEN_17184; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17186 = 10'h17f == _h_T_1 ? ram_383 : _GEN_17185; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17187 = 10'h180 == _h_T_1 ? ram_384 : _GEN_17186; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17188 = 10'h181 == _h_T_1 ? ram_385 : _GEN_17187; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17189 = 10'h182 == _h_T_1 ? ram_386 : _GEN_17188; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17190 = 10'h183 == _h_T_1 ? ram_387 : _GEN_17189; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17191 = 10'h184 == _h_T_1 ? ram_388 : _GEN_17190; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17192 = 10'h185 == _h_T_1 ? ram_389 : _GEN_17191; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17193 = 10'h186 == _h_T_1 ? ram_390 : _GEN_17192; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17194 = 10'h187 == _h_T_1 ? ram_391 : _GEN_17193; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17195 = 10'h188 == _h_T_1 ? ram_392 : _GEN_17194; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17196 = 10'h189 == _h_T_1 ? ram_393 : _GEN_17195; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17197 = 10'h18a == _h_T_1 ? ram_394 : _GEN_17196; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17198 = 10'h18b == _h_T_1 ? ram_395 : _GEN_17197; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17199 = 10'h18c == _h_T_1 ? ram_396 : _GEN_17198; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17200 = 10'h18d == _h_T_1 ? ram_397 : _GEN_17199; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17201 = 10'h18e == _h_T_1 ? ram_398 : _GEN_17200; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17202 = 10'h18f == _h_T_1 ? ram_399 : _GEN_17201; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17203 = 10'h190 == _h_T_1 ? ram_400 : _GEN_17202; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17204 = 10'h191 == _h_T_1 ? ram_401 : _GEN_17203; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17205 = 10'h192 == _h_T_1 ? ram_402 : _GEN_17204; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17206 = 10'h193 == _h_T_1 ? ram_403 : _GEN_17205; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17207 = 10'h194 == _h_T_1 ? ram_404 : _GEN_17206; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17208 = 10'h195 == _h_T_1 ? ram_405 : _GEN_17207; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17209 = 10'h196 == _h_T_1 ? ram_406 : _GEN_17208; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17210 = 10'h197 == _h_T_1 ? ram_407 : _GEN_17209; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17211 = 10'h198 == _h_T_1 ? ram_408 : _GEN_17210; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17212 = 10'h199 == _h_T_1 ? ram_409 : _GEN_17211; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17213 = 10'h19a == _h_T_1 ? ram_410 : _GEN_17212; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17214 = 10'h19b == _h_T_1 ? ram_411 : _GEN_17213; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17215 = 10'h19c == _h_T_1 ? ram_412 : _GEN_17214; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17216 = 10'h19d == _h_T_1 ? ram_413 : _GEN_17215; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17217 = 10'h19e == _h_T_1 ? ram_414 : _GEN_17216; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17218 = 10'h19f == _h_T_1 ? ram_415 : _GEN_17217; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17219 = 10'h1a0 == _h_T_1 ? ram_416 : _GEN_17218; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17220 = 10'h1a1 == _h_T_1 ? ram_417 : _GEN_17219; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17221 = 10'h1a2 == _h_T_1 ? ram_418 : _GEN_17220; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17222 = 10'h1a3 == _h_T_1 ? ram_419 : _GEN_17221; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17223 = 10'h1a4 == _h_T_1 ? ram_420 : _GEN_17222; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17224 = 10'h1a5 == _h_T_1 ? ram_421 : _GEN_17223; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17225 = 10'h1a6 == _h_T_1 ? ram_422 : _GEN_17224; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17226 = 10'h1a7 == _h_T_1 ? ram_423 : _GEN_17225; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17227 = 10'h1a8 == _h_T_1 ? ram_424 : _GEN_17226; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17228 = 10'h1a9 == _h_T_1 ? ram_425 : _GEN_17227; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17229 = 10'h1aa == _h_T_1 ? ram_426 : _GEN_17228; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17230 = 10'h1ab == _h_T_1 ? ram_427 : _GEN_17229; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17231 = 10'h1ac == _h_T_1 ? ram_428 : _GEN_17230; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17232 = 10'h1ad == _h_T_1 ? ram_429 : _GEN_17231; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17233 = 10'h1ae == _h_T_1 ? ram_430 : _GEN_17232; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17234 = 10'h1af == _h_T_1 ? ram_431 : _GEN_17233; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17235 = 10'h1b0 == _h_T_1 ? ram_432 : _GEN_17234; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17236 = 10'h1b1 == _h_T_1 ? ram_433 : _GEN_17235; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17237 = 10'h1b2 == _h_T_1 ? ram_434 : _GEN_17236; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17238 = 10'h1b3 == _h_T_1 ? ram_435 : _GEN_17237; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17239 = 10'h1b4 == _h_T_1 ? ram_436 : _GEN_17238; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17240 = 10'h1b5 == _h_T_1 ? ram_437 : _GEN_17239; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17241 = 10'h1b6 == _h_T_1 ? ram_438 : _GEN_17240; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17242 = 10'h1b7 == _h_T_1 ? ram_439 : _GEN_17241; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17243 = 10'h1b8 == _h_T_1 ? ram_440 : _GEN_17242; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17244 = 10'h1b9 == _h_T_1 ? ram_441 : _GEN_17243; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17245 = 10'h1ba == _h_T_1 ? ram_442 : _GEN_17244; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17246 = 10'h1bb == _h_T_1 ? ram_443 : _GEN_17245; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17247 = 10'h1bc == _h_T_1 ? ram_444 : _GEN_17246; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17248 = 10'h1bd == _h_T_1 ? ram_445 : _GEN_17247; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17249 = 10'h1be == _h_T_1 ? ram_446 : _GEN_17248; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17250 = 10'h1bf == _h_T_1 ? ram_447 : _GEN_17249; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17251 = 10'h1c0 == _h_T_1 ? ram_448 : _GEN_17250; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17252 = 10'h1c1 == _h_T_1 ? ram_449 : _GEN_17251; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17253 = 10'h1c2 == _h_T_1 ? ram_450 : _GEN_17252; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17254 = 10'h1c3 == _h_T_1 ? ram_451 : _GEN_17253; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17255 = 10'h1c4 == _h_T_1 ? ram_452 : _GEN_17254; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17256 = 10'h1c5 == _h_T_1 ? ram_453 : _GEN_17255; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17257 = 10'h1c6 == _h_T_1 ? ram_454 : _GEN_17256; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17258 = 10'h1c7 == _h_T_1 ? ram_455 : _GEN_17257; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17259 = 10'h1c8 == _h_T_1 ? ram_456 : _GEN_17258; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17260 = 10'h1c9 == _h_T_1 ? ram_457 : _GEN_17259; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17261 = 10'h1ca == _h_T_1 ? ram_458 : _GEN_17260; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17262 = 10'h1cb == _h_T_1 ? ram_459 : _GEN_17261; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17263 = 10'h1cc == _h_T_1 ? ram_460 : _GEN_17262; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17264 = 10'h1cd == _h_T_1 ? ram_461 : _GEN_17263; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17265 = 10'h1ce == _h_T_1 ? ram_462 : _GEN_17264; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17266 = 10'h1cf == _h_T_1 ? ram_463 : _GEN_17265; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17267 = 10'h1d0 == _h_T_1 ? ram_464 : _GEN_17266; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17268 = 10'h1d1 == _h_T_1 ? ram_465 : _GEN_17267; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17269 = 10'h1d2 == _h_T_1 ? ram_466 : _GEN_17268; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17270 = 10'h1d3 == _h_T_1 ? ram_467 : _GEN_17269; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17271 = 10'h1d4 == _h_T_1 ? ram_468 : _GEN_17270; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17272 = 10'h1d5 == _h_T_1 ? ram_469 : _GEN_17271; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17273 = 10'h1d6 == _h_T_1 ? ram_470 : _GEN_17272; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17274 = 10'h1d7 == _h_T_1 ? ram_471 : _GEN_17273; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17275 = 10'h1d8 == _h_T_1 ? ram_472 : _GEN_17274; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17276 = 10'h1d9 == _h_T_1 ? ram_473 : _GEN_17275; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17277 = 10'h1da == _h_T_1 ? ram_474 : _GEN_17276; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17278 = 10'h1db == _h_T_1 ? ram_475 : _GEN_17277; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17279 = 10'h1dc == _h_T_1 ? ram_476 : _GEN_17278; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17280 = 10'h1dd == _h_T_1 ? ram_477 : _GEN_17279; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17281 = 10'h1de == _h_T_1 ? ram_478 : _GEN_17280; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17282 = 10'h1df == _h_T_1 ? ram_479 : _GEN_17281; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17283 = 10'h1e0 == _h_T_1 ? ram_480 : _GEN_17282; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17284 = 10'h1e1 == _h_T_1 ? ram_481 : _GEN_17283; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17285 = 10'h1e2 == _h_T_1 ? ram_482 : _GEN_17284; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17286 = 10'h1e3 == _h_T_1 ? ram_483 : _GEN_17285; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17287 = 10'h1e4 == _h_T_1 ? ram_484 : _GEN_17286; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17288 = 10'h1e5 == _h_T_1 ? ram_485 : _GEN_17287; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17289 = 10'h1e6 == _h_T_1 ? ram_486 : _GEN_17288; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17290 = 10'h1e7 == _h_T_1 ? ram_487 : _GEN_17289; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17291 = 10'h1e8 == _h_T_1 ? ram_488 : _GEN_17290; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17292 = 10'h1e9 == _h_T_1 ? ram_489 : _GEN_17291; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17293 = 10'h1ea == _h_T_1 ? ram_490 : _GEN_17292; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17294 = 10'h1eb == _h_T_1 ? ram_491 : _GEN_17293; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17295 = 10'h1ec == _h_T_1 ? ram_492 : _GEN_17294; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17296 = 10'h1ed == _h_T_1 ? ram_493 : _GEN_17295; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17297 = 10'h1ee == _h_T_1 ? ram_494 : _GEN_17296; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17298 = 10'h1ef == _h_T_1 ? ram_495 : _GEN_17297; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17299 = 10'h1f0 == _h_T_1 ? ram_496 : _GEN_17298; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17300 = 10'h1f1 == _h_T_1 ? ram_497 : _GEN_17299; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17301 = 10'h1f2 == _h_T_1 ? ram_498 : _GEN_17300; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17302 = 10'h1f3 == _h_T_1 ? ram_499 : _GEN_17301; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17303 = 10'h1f4 == _h_T_1 ? ram_500 : _GEN_17302; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17304 = 10'h1f5 == _h_T_1 ? ram_501 : _GEN_17303; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17305 = 10'h1f6 == _h_T_1 ? ram_502 : _GEN_17304; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17306 = 10'h1f7 == _h_T_1 ? ram_503 : _GEN_17305; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17307 = 10'h1f8 == _h_T_1 ? ram_504 : _GEN_17306; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17308 = 10'h1f9 == _h_T_1 ? ram_505 : _GEN_17307; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17309 = 10'h1fa == _h_T_1 ? ram_506 : _GEN_17308; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17310 = 10'h1fb == _h_T_1 ? ram_507 : _GEN_17309; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17311 = 10'h1fc == _h_T_1 ? ram_508 : _GEN_17310; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17312 = 10'h1fd == _h_T_1 ? ram_509 : _GEN_17311; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17313 = 10'h1fe == _h_T_1 ? ram_510 : _GEN_17312; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17314 = 10'h1ff == _h_T_1 ? ram_511 : _GEN_17313; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17315 = 10'h200 == _h_T_1 ? ram_512 : _GEN_17314; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17316 = 10'h201 == _h_T_1 ? ram_513 : _GEN_17315; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17317 = 10'h202 == _h_T_1 ? ram_514 : _GEN_17316; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17318 = 10'h203 == _h_T_1 ? ram_515 : _GEN_17317; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17319 = 10'h204 == _h_T_1 ? ram_516 : _GEN_17318; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17320 = 10'h205 == _h_T_1 ? ram_517 : _GEN_17319; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17321 = 10'h206 == _h_T_1 ? ram_518 : _GEN_17320; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17322 = 10'h207 == _h_T_1 ? ram_519 : _GEN_17321; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17323 = 10'h208 == _h_T_1 ? ram_520 : _GEN_17322; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17324 = 10'h209 == _h_T_1 ? ram_521 : _GEN_17323; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17325 = 10'h20a == _h_T_1 ? ram_522 : _GEN_17324; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17326 = 10'h20b == _h_T_1 ? ram_523 : _GEN_17325; // @[vga.scala 64:41 vga.scala 64:41]
  wire [287:0] _GEN_17327 = 10'h20c == _h_T_1 ? ram_524 : _GEN_17326; // @[vga.scala 64:41 vga.scala 64:41]
  wire [8477:0] _GEN_19093 = {{8190'd0}, _GEN_17327}; // @[vga.scala 64:41]
  wire [8477:0] _ram_T_441 = _GEN_19093 ^ _ram_T_440; // @[vga.scala 64:41]
  wire [8:0] _v_T_1 = v + 9'h9; // @[vga.scala 66:13]
  reg [23:0] rdwrPort; // @[vga.scala 68:23]
  wire [287:0] _GEN_18535 = 10'h1 == io_h_addr ? ram_1 : ram_0; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18536 = 10'h2 == io_h_addr ? ram_2 : _GEN_18535; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18537 = 10'h3 == io_h_addr ? ram_3 : _GEN_18536; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18538 = 10'h4 == io_h_addr ? ram_4 : _GEN_18537; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18539 = 10'h5 == io_h_addr ? ram_5 : _GEN_18538; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18540 = 10'h6 == io_h_addr ? ram_6 : _GEN_18539; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18541 = 10'h7 == io_h_addr ? ram_7 : _GEN_18540; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18542 = 10'h8 == io_h_addr ? ram_8 : _GEN_18541; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18543 = 10'h9 == io_h_addr ? ram_9 : _GEN_18542; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18544 = 10'ha == io_h_addr ? ram_10 : _GEN_18543; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18545 = 10'hb == io_h_addr ? ram_11 : _GEN_18544; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18546 = 10'hc == io_h_addr ? ram_12 : _GEN_18545; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18547 = 10'hd == io_h_addr ? ram_13 : _GEN_18546; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18548 = 10'he == io_h_addr ? ram_14 : _GEN_18547; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18549 = 10'hf == io_h_addr ? ram_15 : _GEN_18548; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18550 = 10'h10 == io_h_addr ? ram_16 : _GEN_18549; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18551 = 10'h11 == io_h_addr ? ram_17 : _GEN_18550; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18552 = 10'h12 == io_h_addr ? ram_18 : _GEN_18551; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18553 = 10'h13 == io_h_addr ? ram_19 : _GEN_18552; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18554 = 10'h14 == io_h_addr ? ram_20 : _GEN_18553; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18555 = 10'h15 == io_h_addr ? ram_21 : _GEN_18554; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18556 = 10'h16 == io_h_addr ? ram_22 : _GEN_18555; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18557 = 10'h17 == io_h_addr ? ram_23 : _GEN_18556; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18558 = 10'h18 == io_h_addr ? ram_24 : _GEN_18557; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18559 = 10'h19 == io_h_addr ? ram_25 : _GEN_18558; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18560 = 10'h1a == io_h_addr ? ram_26 : _GEN_18559; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18561 = 10'h1b == io_h_addr ? ram_27 : _GEN_18560; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18562 = 10'h1c == io_h_addr ? ram_28 : _GEN_18561; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18563 = 10'h1d == io_h_addr ? ram_29 : _GEN_18562; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18564 = 10'h1e == io_h_addr ? ram_30 : _GEN_18563; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18565 = 10'h1f == io_h_addr ? ram_31 : _GEN_18564; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18566 = 10'h20 == io_h_addr ? ram_32 : _GEN_18565; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18567 = 10'h21 == io_h_addr ? ram_33 : _GEN_18566; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18568 = 10'h22 == io_h_addr ? ram_34 : _GEN_18567; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18569 = 10'h23 == io_h_addr ? ram_35 : _GEN_18568; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18570 = 10'h24 == io_h_addr ? ram_36 : _GEN_18569; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18571 = 10'h25 == io_h_addr ? ram_37 : _GEN_18570; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18572 = 10'h26 == io_h_addr ? ram_38 : _GEN_18571; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18573 = 10'h27 == io_h_addr ? ram_39 : _GEN_18572; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18574 = 10'h28 == io_h_addr ? ram_40 : _GEN_18573; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18575 = 10'h29 == io_h_addr ? ram_41 : _GEN_18574; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18576 = 10'h2a == io_h_addr ? ram_42 : _GEN_18575; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18577 = 10'h2b == io_h_addr ? ram_43 : _GEN_18576; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18578 = 10'h2c == io_h_addr ? ram_44 : _GEN_18577; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18579 = 10'h2d == io_h_addr ? ram_45 : _GEN_18578; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18580 = 10'h2e == io_h_addr ? ram_46 : _GEN_18579; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18581 = 10'h2f == io_h_addr ? ram_47 : _GEN_18580; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18582 = 10'h30 == io_h_addr ? ram_48 : _GEN_18581; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18583 = 10'h31 == io_h_addr ? ram_49 : _GEN_18582; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18584 = 10'h32 == io_h_addr ? ram_50 : _GEN_18583; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18585 = 10'h33 == io_h_addr ? ram_51 : _GEN_18584; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18586 = 10'h34 == io_h_addr ? ram_52 : _GEN_18585; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18587 = 10'h35 == io_h_addr ? ram_53 : _GEN_18586; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18588 = 10'h36 == io_h_addr ? ram_54 : _GEN_18587; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18589 = 10'h37 == io_h_addr ? ram_55 : _GEN_18588; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18590 = 10'h38 == io_h_addr ? ram_56 : _GEN_18589; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18591 = 10'h39 == io_h_addr ? ram_57 : _GEN_18590; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18592 = 10'h3a == io_h_addr ? ram_58 : _GEN_18591; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18593 = 10'h3b == io_h_addr ? ram_59 : _GEN_18592; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18594 = 10'h3c == io_h_addr ? ram_60 : _GEN_18593; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18595 = 10'h3d == io_h_addr ? ram_61 : _GEN_18594; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18596 = 10'h3e == io_h_addr ? ram_62 : _GEN_18595; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18597 = 10'h3f == io_h_addr ? ram_63 : _GEN_18596; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18598 = 10'h40 == io_h_addr ? ram_64 : _GEN_18597; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18599 = 10'h41 == io_h_addr ? ram_65 : _GEN_18598; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18600 = 10'h42 == io_h_addr ? ram_66 : _GEN_18599; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18601 = 10'h43 == io_h_addr ? ram_67 : _GEN_18600; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18602 = 10'h44 == io_h_addr ? ram_68 : _GEN_18601; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18603 = 10'h45 == io_h_addr ? ram_69 : _GEN_18602; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18604 = 10'h46 == io_h_addr ? ram_70 : _GEN_18603; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18605 = 10'h47 == io_h_addr ? ram_71 : _GEN_18604; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18606 = 10'h48 == io_h_addr ? ram_72 : _GEN_18605; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18607 = 10'h49 == io_h_addr ? ram_73 : _GEN_18606; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18608 = 10'h4a == io_h_addr ? ram_74 : _GEN_18607; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18609 = 10'h4b == io_h_addr ? ram_75 : _GEN_18608; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18610 = 10'h4c == io_h_addr ? ram_76 : _GEN_18609; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18611 = 10'h4d == io_h_addr ? ram_77 : _GEN_18610; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18612 = 10'h4e == io_h_addr ? ram_78 : _GEN_18611; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18613 = 10'h4f == io_h_addr ? ram_79 : _GEN_18612; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18614 = 10'h50 == io_h_addr ? ram_80 : _GEN_18613; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18615 = 10'h51 == io_h_addr ? ram_81 : _GEN_18614; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18616 = 10'h52 == io_h_addr ? ram_82 : _GEN_18615; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18617 = 10'h53 == io_h_addr ? ram_83 : _GEN_18616; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18618 = 10'h54 == io_h_addr ? ram_84 : _GEN_18617; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18619 = 10'h55 == io_h_addr ? ram_85 : _GEN_18618; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18620 = 10'h56 == io_h_addr ? ram_86 : _GEN_18619; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18621 = 10'h57 == io_h_addr ? ram_87 : _GEN_18620; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18622 = 10'h58 == io_h_addr ? ram_88 : _GEN_18621; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18623 = 10'h59 == io_h_addr ? ram_89 : _GEN_18622; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18624 = 10'h5a == io_h_addr ? ram_90 : _GEN_18623; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18625 = 10'h5b == io_h_addr ? ram_91 : _GEN_18624; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18626 = 10'h5c == io_h_addr ? ram_92 : _GEN_18625; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18627 = 10'h5d == io_h_addr ? ram_93 : _GEN_18626; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18628 = 10'h5e == io_h_addr ? ram_94 : _GEN_18627; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18629 = 10'h5f == io_h_addr ? ram_95 : _GEN_18628; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18630 = 10'h60 == io_h_addr ? ram_96 : _GEN_18629; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18631 = 10'h61 == io_h_addr ? ram_97 : _GEN_18630; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18632 = 10'h62 == io_h_addr ? ram_98 : _GEN_18631; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18633 = 10'h63 == io_h_addr ? ram_99 : _GEN_18632; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18634 = 10'h64 == io_h_addr ? ram_100 : _GEN_18633; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18635 = 10'h65 == io_h_addr ? ram_101 : _GEN_18634; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18636 = 10'h66 == io_h_addr ? ram_102 : _GEN_18635; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18637 = 10'h67 == io_h_addr ? ram_103 : _GEN_18636; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18638 = 10'h68 == io_h_addr ? ram_104 : _GEN_18637; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18639 = 10'h69 == io_h_addr ? ram_105 : _GEN_18638; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18640 = 10'h6a == io_h_addr ? ram_106 : _GEN_18639; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18641 = 10'h6b == io_h_addr ? ram_107 : _GEN_18640; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18642 = 10'h6c == io_h_addr ? ram_108 : _GEN_18641; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18643 = 10'h6d == io_h_addr ? ram_109 : _GEN_18642; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18644 = 10'h6e == io_h_addr ? ram_110 : _GEN_18643; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18645 = 10'h6f == io_h_addr ? ram_111 : _GEN_18644; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18646 = 10'h70 == io_h_addr ? ram_112 : _GEN_18645; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18647 = 10'h71 == io_h_addr ? ram_113 : _GEN_18646; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18648 = 10'h72 == io_h_addr ? ram_114 : _GEN_18647; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18649 = 10'h73 == io_h_addr ? ram_115 : _GEN_18648; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18650 = 10'h74 == io_h_addr ? ram_116 : _GEN_18649; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18651 = 10'h75 == io_h_addr ? ram_117 : _GEN_18650; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18652 = 10'h76 == io_h_addr ? ram_118 : _GEN_18651; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18653 = 10'h77 == io_h_addr ? ram_119 : _GEN_18652; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18654 = 10'h78 == io_h_addr ? ram_120 : _GEN_18653; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18655 = 10'h79 == io_h_addr ? ram_121 : _GEN_18654; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18656 = 10'h7a == io_h_addr ? ram_122 : _GEN_18655; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18657 = 10'h7b == io_h_addr ? ram_123 : _GEN_18656; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18658 = 10'h7c == io_h_addr ? ram_124 : _GEN_18657; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18659 = 10'h7d == io_h_addr ? ram_125 : _GEN_18658; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18660 = 10'h7e == io_h_addr ? ram_126 : _GEN_18659; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18661 = 10'h7f == io_h_addr ? ram_127 : _GEN_18660; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18662 = 10'h80 == io_h_addr ? ram_128 : _GEN_18661; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18663 = 10'h81 == io_h_addr ? ram_129 : _GEN_18662; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18664 = 10'h82 == io_h_addr ? ram_130 : _GEN_18663; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18665 = 10'h83 == io_h_addr ? ram_131 : _GEN_18664; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18666 = 10'h84 == io_h_addr ? ram_132 : _GEN_18665; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18667 = 10'h85 == io_h_addr ? ram_133 : _GEN_18666; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18668 = 10'h86 == io_h_addr ? ram_134 : _GEN_18667; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18669 = 10'h87 == io_h_addr ? ram_135 : _GEN_18668; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18670 = 10'h88 == io_h_addr ? ram_136 : _GEN_18669; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18671 = 10'h89 == io_h_addr ? ram_137 : _GEN_18670; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18672 = 10'h8a == io_h_addr ? ram_138 : _GEN_18671; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18673 = 10'h8b == io_h_addr ? ram_139 : _GEN_18672; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18674 = 10'h8c == io_h_addr ? ram_140 : _GEN_18673; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18675 = 10'h8d == io_h_addr ? ram_141 : _GEN_18674; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18676 = 10'h8e == io_h_addr ? ram_142 : _GEN_18675; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18677 = 10'h8f == io_h_addr ? ram_143 : _GEN_18676; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18678 = 10'h90 == io_h_addr ? ram_144 : _GEN_18677; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18679 = 10'h91 == io_h_addr ? ram_145 : _GEN_18678; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18680 = 10'h92 == io_h_addr ? ram_146 : _GEN_18679; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18681 = 10'h93 == io_h_addr ? ram_147 : _GEN_18680; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18682 = 10'h94 == io_h_addr ? ram_148 : _GEN_18681; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18683 = 10'h95 == io_h_addr ? ram_149 : _GEN_18682; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18684 = 10'h96 == io_h_addr ? ram_150 : _GEN_18683; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18685 = 10'h97 == io_h_addr ? ram_151 : _GEN_18684; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18686 = 10'h98 == io_h_addr ? ram_152 : _GEN_18685; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18687 = 10'h99 == io_h_addr ? ram_153 : _GEN_18686; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18688 = 10'h9a == io_h_addr ? ram_154 : _GEN_18687; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18689 = 10'h9b == io_h_addr ? ram_155 : _GEN_18688; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18690 = 10'h9c == io_h_addr ? ram_156 : _GEN_18689; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18691 = 10'h9d == io_h_addr ? ram_157 : _GEN_18690; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18692 = 10'h9e == io_h_addr ? ram_158 : _GEN_18691; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18693 = 10'h9f == io_h_addr ? ram_159 : _GEN_18692; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18694 = 10'ha0 == io_h_addr ? ram_160 : _GEN_18693; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18695 = 10'ha1 == io_h_addr ? ram_161 : _GEN_18694; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18696 = 10'ha2 == io_h_addr ? ram_162 : _GEN_18695; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18697 = 10'ha3 == io_h_addr ? ram_163 : _GEN_18696; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18698 = 10'ha4 == io_h_addr ? ram_164 : _GEN_18697; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18699 = 10'ha5 == io_h_addr ? ram_165 : _GEN_18698; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18700 = 10'ha6 == io_h_addr ? ram_166 : _GEN_18699; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18701 = 10'ha7 == io_h_addr ? ram_167 : _GEN_18700; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18702 = 10'ha8 == io_h_addr ? ram_168 : _GEN_18701; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18703 = 10'ha9 == io_h_addr ? ram_169 : _GEN_18702; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18704 = 10'haa == io_h_addr ? ram_170 : _GEN_18703; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18705 = 10'hab == io_h_addr ? ram_171 : _GEN_18704; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18706 = 10'hac == io_h_addr ? ram_172 : _GEN_18705; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18707 = 10'had == io_h_addr ? ram_173 : _GEN_18706; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18708 = 10'hae == io_h_addr ? ram_174 : _GEN_18707; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18709 = 10'haf == io_h_addr ? ram_175 : _GEN_18708; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18710 = 10'hb0 == io_h_addr ? ram_176 : _GEN_18709; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18711 = 10'hb1 == io_h_addr ? ram_177 : _GEN_18710; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18712 = 10'hb2 == io_h_addr ? ram_178 : _GEN_18711; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18713 = 10'hb3 == io_h_addr ? ram_179 : _GEN_18712; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18714 = 10'hb4 == io_h_addr ? ram_180 : _GEN_18713; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18715 = 10'hb5 == io_h_addr ? ram_181 : _GEN_18714; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18716 = 10'hb6 == io_h_addr ? ram_182 : _GEN_18715; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18717 = 10'hb7 == io_h_addr ? ram_183 : _GEN_18716; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18718 = 10'hb8 == io_h_addr ? ram_184 : _GEN_18717; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18719 = 10'hb9 == io_h_addr ? ram_185 : _GEN_18718; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18720 = 10'hba == io_h_addr ? ram_186 : _GEN_18719; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18721 = 10'hbb == io_h_addr ? ram_187 : _GEN_18720; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18722 = 10'hbc == io_h_addr ? ram_188 : _GEN_18721; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18723 = 10'hbd == io_h_addr ? ram_189 : _GEN_18722; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18724 = 10'hbe == io_h_addr ? ram_190 : _GEN_18723; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18725 = 10'hbf == io_h_addr ? ram_191 : _GEN_18724; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18726 = 10'hc0 == io_h_addr ? ram_192 : _GEN_18725; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18727 = 10'hc1 == io_h_addr ? ram_193 : _GEN_18726; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18728 = 10'hc2 == io_h_addr ? ram_194 : _GEN_18727; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18729 = 10'hc3 == io_h_addr ? ram_195 : _GEN_18728; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18730 = 10'hc4 == io_h_addr ? ram_196 : _GEN_18729; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18731 = 10'hc5 == io_h_addr ? ram_197 : _GEN_18730; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18732 = 10'hc6 == io_h_addr ? ram_198 : _GEN_18731; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18733 = 10'hc7 == io_h_addr ? ram_199 : _GEN_18732; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18734 = 10'hc8 == io_h_addr ? ram_200 : _GEN_18733; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18735 = 10'hc9 == io_h_addr ? ram_201 : _GEN_18734; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18736 = 10'hca == io_h_addr ? ram_202 : _GEN_18735; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18737 = 10'hcb == io_h_addr ? ram_203 : _GEN_18736; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18738 = 10'hcc == io_h_addr ? ram_204 : _GEN_18737; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18739 = 10'hcd == io_h_addr ? ram_205 : _GEN_18738; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18740 = 10'hce == io_h_addr ? ram_206 : _GEN_18739; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18741 = 10'hcf == io_h_addr ? ram_207 : _GEN_18740; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18742 = 10'hd0 == io_h_addr ? ram_208 : _GEN_18741; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18743 = 10'hd1 == io_h_addr ? ram_209 : _GEN_18742; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18744 = 10'hd2 == io_h_addr ? ram_210 : _GEN_18743; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18745 = 10'hd3 == io_h_addr ? ram_211 : _GEN_18744; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18746 = 10'hd4 == io_h_addr ? ram_212 : _GEN_18745; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18747 = 10'hd5 == io_h_addr ? ram_213 : _GEN_18746; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18748 = 10'hd6 == io_h_addr ? ram_214 : _GEN_18747; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18749 = 10'hd7 == io_h_addr ? ram_215 : _GEN_18748; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18750 = 10'hd8 == io_h_addr ? ram_216 : _GEN_18749; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18751 = 10'hd9 == io_h_addr ? ram_217 : _GEN_18750; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18752 = 10'hda == io_h_addr ? ram_218 : _GEN_18751; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18753 = 10'hdb == io_h_addr ? ram_219 : _GEN_18752; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18754 = 10'hdc == io_h_addr ? ram_220 : _GEN_18753; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18755 = 10'hdd == io_h_addr ? ram_221 : _GEN_18754; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18756 = 10'hde == io_h_addr ? ram_222 : _GEN_18755; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18757 = 10'hdf == io_h_addr ? ram_223 : _GEN_18756; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18758 = 10'he0 == io_h_addr ? ram_224 : _GEN_18757; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18759 = 10'he1 == io_h_addr ? ram_225 : _GEN_18758; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18760 = 10'he2 == io_h_addr ? ram_226 : _GEN_18759; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18761 = 10'he3 == io_h_addr ? ram_227 : _GEN_18760; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18762 = 10'he4 == io_h_addr ? ram_228 : _GEN_18761; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18763 = 10'he5 == io_h_addr ? ram_229 : _GEN_18762; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18764 = 10'he6 == io_h_addr ? ram_230 : _GEN_18763; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18765 = 10'he7 == io_h_addr ? ram_231 : _GEN_18764; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18766 = 10'he8 == io_h_addr ? ram_232 : _GEN_18765; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18767 = 10'he9 == io_h_addr ? ram_233 : _GEN_18766; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18768 = 10'hea == io_h_addr ? ram_234 : _GEN_18767; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18769 = 10'heb == io_h_addr ? ram_235 : _GEN_18768; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18770 = 10'hec == io_h_addr ? ram_236 : _GEN_18769; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18771 = 10'hed == io_h_addr ? ram_237 : _GEN_18770; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18772 = 10'hee == io_h_addr ? ram_238 : _GEN_18771; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18773 = 10'hef == io_h_addr ? ram_239 : _GEN_18772; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18774 = 10'hf0 == io_h_addr ? ram_240 : _GEN_18773; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18775 = 10'hf1 == io_h_addr ? ram_241 : _GEN_18774; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18776 = 10'hf2 == io_h_addr ? ram_242 : _GEN_18775; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18777 = 10'hf3 == io_h_addr ? ram_243 : _GEN_18776; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18778 = 10'hf4 == io_h_addr ? ram_244 : _GEN_18777; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18779 = 10'hf5 == io_h_addr ? ram_245 : _GEN_18778; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18780 = 10'hf6 == io_h_addr ? ram_246 : _GEN_18779; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18781 = 10'hf7 == io_h_addr ? ram_247 : _GEN_18780; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18782 = 10'hf8 == io_h_addr ? ram_248 : _GEN_18781; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18783 = 10'hf9 == io_h_addr ? ram_249 : _GEN_18782; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18784 = 10'hfa == io_h_addr ? ram_250 : _GEN_18783; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18785 = 10'hfb == io_h_addr ? ram_251 : _GEN_18784; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18786 = 10'hfc == io_h_addr ? ram_252 : _GEN_18785; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18787 = 10'hfd == io_h_addr ? ram_253 : _GEN_18786; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18788 = 10'hfe == io_h_addr ? ram_254 : _GEN_18787; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18789 = 10'hff == io_h_addr ? ram_255 : _GEN_18788; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18790 = 10'h100 == io_h_addr ? ram_256 : _GEN_18789; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18791 = 10'h101 == io_h_addr ? ram_257 : _GEN_18790; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18792 = 10'h102 == io_h_addr ? ram_258 : _GEN_18791; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18793 = 10'h103 == io_h_addr ? ram_259 : _GEN_18792; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18794 = 10'h104 == io_h_addr ? ram_260 : _GEN_18793; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18795 = 10'h105 == io_h_addr ? ram_261 : _GEN_18794; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18796 = 10'h106 == io_h_addr ? ram_262 : _GEN_18795; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18797 = 10'h107 == io_h_addr ? ram_263 : _GEN_18796; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18798 = 10'h108 == io_h_addr ? ram_264 : _GEN_18797; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18799 = 10'h109 == io_h_addr ? ram_265 : _GEN_18798; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18800 = 10'h10a == io_h_addr ? ram_266 : _GEN_18799; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18801 = 10'h10b == io_h_addr ? ram_267 : _GEN_18800; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18802 = 10'h10c == io_h_addr ? ram_268 : _GEN_18801; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18803 = 10'h10d == io_h_addr ? ram_269 : _GEN_18802; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18804 = 10'h10e == io_h_addr ? ram_270 : _GEN_18803; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18805 = 10'h10f == io_h_addr ? ram_271 : _GEN_18804; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18806 = 10'h110 == io_h_addr ? ram_272 : _GEN_18805; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18807 = 10'h111 == io_h_addr ? ram_273 : _GEN_18806; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18808 = 10'h112 == io_h_addr ? ram_274 : _GEN_18807; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18809 = 10'h113 == io_h_addr ? ram_275 : _GEN_18808; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18810 = 10'h114 == io_h_addr ? ram_276 : _GEN_18809; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18811 = 10'h115 == io_h_addr ? ram_277 : _GEN_18810; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18812 = 10'h116 == io_h_addr ? ram_278 : _GEN_18811; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18813 = 10'h117 == io_h_addr ? ram_279 : _GEN_18812; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18814 = 10'h118 == io_h_addr ? ram_280 : _GEN_18813; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18815 = 10'h119 == io_h_addr ? ram_281 : _GEN_18814; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18816 = 10'h11a == io_h_addr ? ram_282 : _GEN_18815; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18817 = 10'h11b == io_h_addr ? ram_283 : _GEN_18816; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18818 = 10'h11c == io_h_addr ? ram_284 : _GEN_18817; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18819 = 10'h11d == io_h_addr ? ram_285 : _GEN_18818; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18820 = 10'h11e == io_h_addr ? ram_286 : _GEN_18819; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18821 = 10'h11f == io_h_addr ? ram_287 : _GEN_18820; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18822 = 10'h120 == io_h_addr ? ram_288 : _GEN_18821; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18823 = 10'h121 == io_h_addr ? ram_289 : _GEN_18822; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18824 = 10'h122 == io_h_addr ? ram_290 : _GEN_18823; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18825 = 10'h123 == io_h_addr ? ram_291 : _GEN_18824; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18826 = 10'h124 == io_h_addr ? ram_292 : _GEN_18825; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18827 = 10'h125 == io_h_addr ? ram_293 : _GEN_18826; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18828 = 10'h126 == io_h_addr ? ram_294 : _GEN_18827; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18829 = 10'h127 == io_h_addr ? ram_295 : _GEN_18828; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18830 = 10'h128 == io_h_addr ? ram_296 : _GEN_18829; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18831 = 10'h129 == io_h_addr ? ram_297 : _GEN_18830; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18832 = 10'h12a == io_h_addr ? ram_298 : _GEN_18831; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18833 = 10'h12b == io_h_addr ? ram_299 : _GEN_18832; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18834 = 10'h12c == io_h_addr ? ram_300 : _GEN_18833; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18835 = 10'h12d == io_h_addr ? ram_301 : _GEN_18834; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18836 = 10'h12e == io_h_addr ? ram_302 : _GEN_18835; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18837 = 10'h12f == io_h_addr ? ram_303 : _GEN_18836; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18838 = 10'h130 == io_h_addr ? ram_304 : _GEN_18837; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18839 = 10'h131 == io_h_addr ? ram_305 : _GEN_18838; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18840 = 10'h132 == io_h_addr ? ram_306 : _GEN_18839; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18841 = 10'h133 == io_h_addr ? ram_307 : _GEN_18840; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18842 = 10'h134 == io_h_addr ? ram_308 : _GEN_18841; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18843 = 10'h135 == io_h_addr ? ram_309 : _GEN_18842; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18844 = 10'h136 == io_h_addr ? ram_310 : _GEN_18843; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18845 = 10'h137 == io_h_addr ? ram_311 : _GEN_18844; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18846 = 10'h138 == io_h_addr ? ram_312 : _GEN_18845; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18847 = 10'h139 == io_h_addr ? ram_313 : _GEN_18846; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18848 = 10'h13a == io_h_addr ? ram_314 : _GEN_18847; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18849 = 10'h13b == io_h_addr ? ram_315 : _GEN_18848; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18850 = 10'h13c == io_h_addr ? ram_316 : _GEN_18849; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18851 = 10'h13d == io_h_addr ? ram_317 : _GEN_18850; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18852 = 10'h13e == io_h_addr ? ram_318 : _GEN_18851; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18853 = 10'h13f == io_h_addr ? ram_319 : _GEN_18852; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18854 = 10'h140 == io_h_addr ? ram_320 : _GEN_18853; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18855 = 10'h141 == io_h_addr ? ram_321 : _GEN_18854; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18856 = 10'h142 == io_h_addr ? ram_322 : _GEN_18855; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18857 = 10'h143 == io_h_addr ? ram_323 : _GEN_18856; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18858 = 10'h144 == io_h_addr ? ram_324 : _GEN_18857; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18859 = 10'h145 == io_h_addr ? ram_325 : _GEN_18858; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18860 = 10'h146 == io_h_addr ? ram_326 : _GEN_18859; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18861 = 10'h147 == io_h_addr ? ram_327 : _GEN_18860; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18862 = 10'h148 == io_h_addr ? ram_328 : _GEN_18861; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18863 = 10'h149 == io_h_addr ? ram_329 : _GEN_18862; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18864 = 10'h14a == io_h_addr ? ram_330 : _GEN_18863; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18865 = 10'h14b == io_h_addr ? ram_331 : _GEN_18864; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18866 = 10'h14c == io_h_addr ? ram_332 : _GEN_18865; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18867 = 10'h14d == io_h_addr ? ram_333 : _GEN_18866; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18868 = 10'h14e == io_h_addr ? ram_334 : _GEN_18867; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18869 = 10'h14f == io_h_addr ? ram_335 : _GEN_18868; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18870 = 10'h150 == io_h_addr ? ram_336 : _GEN_18869; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18871 = 10'h151 == io_h_addr ? ram_337 : _GEN_18870; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18872 = 10'h152 == io_h_addr ? ram_338 : _GEN_18871; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18873 = 10'h153 == io_h_addr ? ram_339 : _GEN_18872; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18874 = 10'h154 == io_h_addr ? ram_340 : _GEN_18873; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18875 = 10'h155 == io_h_addr ? ram_341 : _GEN_18874; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18876 = 10'h156 == io_h_addr ? ram_342 : _GEN_18875; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18877 = 10'h157 == io_h_addr ? ram_343 : _GEN_18876; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18878 = 10'h158 == io_h_addr ? ram_344 : _GEN_18877; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18879 = 10'h159 == io_h_addr ? ram_345 : _GEN_18878; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18880 = 10'h15a == io_h_addr ? ram_346 : _GEN_18879; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18881 = 10'h15b == io_h_addr ? ram_347 : _GEN_18880; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18882 = 10'h15c == io_h_addr ? ram_348 : _GEN_18881; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18883 = 10'h15d == io_h_addr ? ram_349 : _GEN_18882; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18884 = 10'h15e == io_h_addr ? ram_350 : _GEN_18883; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18885 = 10'h15f == io_h_addr ? ram_351 : _GEN_18884; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18886 = 10'h160 == io_h_addr ? ram_352 : _GEN_18885; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18887 = 10'h161 == io_h_addr ? ram_353 : _GEN_18886; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18888 = 10'h162 == io_h_addr ? ram_354 : _GEN_18887; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18889 = 10'h163 == io_h_addr ? ram_355 : _GEN_18888; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18890 = 10'h164 == io_h_addr ? ram_356 : _GEN_18889; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18891 = 10'h165 == io_h_addr ? ram_357 : _GEN_18890; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18892 = 10'h166 == io_h_addr ? ram_358 : _GEN_18891; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18893 = 10'h167 == io_h_addr ? ram_359 : _GEN_18892; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18894 = 10'h168 == io_h_addr ? ram_360 : _GEN_18893; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18895 = 10'h169 == io_h_addr ? ram_361 : _GEN_18894; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18896 = 10'h16a == io_h_addr ? ram_362 : _GEN_18895; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18897 = 10'h16b == io_h_addr ? ram_363 : _GEN_18896; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18898 = 10'h16c == io_h_addr ? ram_364 : _GEN_18897; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18899 = 10'h16d == io_h_addr ? ram_365 : _GEN_18898; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18900 = 10'h16e == io_h_addr ? ram_366 : _GEN_18899; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18901 = 10'h16f == io_h_addr ? ram_367 : _GEN_18900; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18902 = 10'h170 == io_h_addr ? ram_368 : _GEN_18901; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18903 = 10'h171 == io_h_addr ? ram_369 : _GEN_18902; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18904 = 10'h172 == io_h_addr ? ram_370 : _GEN_18903; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18905 = 10'h173 == io_h_addr ? ram_371 : _GEN_18904; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18906 = 10'h174 == io_h_addr ? ram_372 : _GEN_18905; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18907 = 10'h175 == io_h_addr ? ram_373 : _GEN_18906; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18908 = 10'h176 == io_h_addr ? ram_374 : _GEN_18907; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18909 = 10'h177 == io_h_addr ? ram_375 : _GEN_18908; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18910 = 10'h178 == io_h_addr ? ram_376 : _GEN_18909; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18911 = 10'h179 == io_h_addr ? ram_377 : _GEN_18910; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18912 = 10'h17a == io_h_addr ? ram_378 : _GEN_18911; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18913 = 10'h17b == io_h_addr ? ram_379 : _GEN_18912; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18914 = 10'h17c == io_h_addr ? ram_380 : _GEN_18913; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18915 = 10'h17d == io_h_addr ? ram_381 : _GEN_18914; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18916 = 10'h17e == io_h_addr ? ram_382 : _GEN_18915; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18917 = 10'h17f == io_h_addr ? ram_383 : _GEN_18916; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18918 = 10'h180 == io_h_addr ? ram_384 : _GEN_18917; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18919 = 10'h181 == io_h_addr ? ram_385 : _GEN_18918; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18920 = 10'h182 == io_h_addr ? ram_386 : _GEN_18919; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18921 = 10'h183 == io_h_addr ? ram_387 : _GEN_18920; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18922 = 10'h184 == io_h_addr ? ram_388 : _GEN_18921; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18923 = 10'h185 == io_h_addr ? ram_389 : _GEN_18922; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18924 = 10'h186 == io_h_addr ? ram_390 : _GEN_18923; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18925 = 10'h187 == io_h_addr ? ram_391 : _GEN_18924; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18926 = 10'h188 == io_h_addr ? ram_392 : _GEN_18925; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18927 = 10'h189 == io_h_addr ? ram_393 : _GEN_18926; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18928 = 10'h18a == io_h_addr ? ram_394 : _GEN_18927; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18929 = 10'h18b == io_h_addr ? ram_395 : _GEN_18928; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18930 = 10'h18c == io_h_addr ? ram_396 : _GEN_18929; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18931 = 10'h18d == io_h_addr ? ram_397 : _GEN_18930; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18932 = 10'h18e == io_h_addr ? ram_398 : _GEN_18931; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18933 = 10'h18f == io_h_addr ? ram_399 : _GEN_18932; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18934 = 10'h190 == io_h_addr ? ram_400 : _GEN_18933; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18935 = 10'h191 == io_h_addr ? ram_401 : _GEN_18934; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18936 = 10'h192 == io_h_addr ? ram_402 : _GEN_18935; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18937 = 10'h193 == io_h_addr ? ram_403 : _GEN_18936; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18938 = 10'h194 == io_h_addr ? ram_404 : _GEN_18937; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18939 = 10'h195 == io_h_addr ? ram_405 : _GEN_18938; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18940 = 10'h196 == io_h_addr ? ram_406 : _GEN_18939; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18941 = 10'h197 == io_h_addr ? ram_407 : _GEN_18940; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18942 = 10'h198 == io_h_addr ? ram_408 : _GEN_18941; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18943 = 10'h199 == io_h_addr ? ram_409 : _GEN_18942; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18944 = 10'h19a == io_h_addr ? ram_410 : _GEN_18943; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18945 = 10'h19b == io_h_addr ? ram_411 : _GEN_18944; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18946 = 10'h19c == io_h_addr ? ram_412 : _GEN_18945; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18947 = 10'h19d == io_h_addr ? ram_413 : _GEN_18946; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18948 = 10'h19e == io_h_addr ? ram_414 : _GEN_18947; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18949 = 10'h19f == io_h_addr ? ram_415 : _GEN_18948; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18950 = 10'h1a0 == io_h_addr ? ram_416 : _GEN_18949; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18951 = 10'h1a1 == io_h_addr ? ram_417 : _GEN_18950; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18952 = 10'h1a2 == io_h_addr ? ram_418 : _GEN_18951; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18953 = 10'h1a3 == io_h_addr ? ram_419 : _GEN_18952; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18954 = 10'h1a4 == io_h_addr ? ram_420 : _GEN_18953; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18955 = 10'h1a5 == io_h_addr ? ram_421 : _GEN_18954; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18956 = 10'h1a6 == io_h_addr ? ram_422 : _GEN_18955; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18957 = 10'h1a7 == io_h_addr ? ram_423 : _GEN_18956; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18958 = 10'h1a8 == io_h_addr ? ram_424 : _GEN_18957; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18959 = 10'h1a9 == io_h_addr ? ram_425 : _GEN_18958; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18960 = 10'h1aa == io_h_addr ? ram_426 : _GEN_18959; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18961 = 10'h1ab == io_h_addr ? ram_427 : _GEN_18960; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18962 = 10'h1ac == io_h_addr ? ram_428 : _GEN_18961; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18963 = 10'h1ad == io_h_addr ? ram_429 : _GEN_18962; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18964 = 10'h1ae == io_h_addr ? ram_430 : _GEN_18963; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18965 = 10'h1af == io_h_addr ? ram_431 : _GEN_18964; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18966 = 10'h1b0 == io_h_addr ? ram_432 : _GEN_18965; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18967 = 10'h1b1 == io_h_addr ? ram_433 : _GEN_18966; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18968 = 10'h1b2 == io_h_addr ? ram_434 : _GEN_18967; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18969 = 10'h1b3 == io_h_addr ? ram_435 : _GEN_18968; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18970 = 10'h1b4 == io_h_addr ? ram_436 : _GEN_18969; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18971 = 10'h1b5 == io_h_addr ? ram_437 : _GEN_18970; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18972 = 10'h1b6 == io_h_addr ? ram_438 : _GEN_18971; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18973 = 10'h1b7 == io_h_addr ? ram_439 : _GEN_18972; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18974 = 10'h1b8 == io_h_addr ? ram_440 : _GEN_18973; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18975 = 10'h1b9 == io_h_addr ? ram_441 : _GEN_18974; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18976 = 10'h1ba == io_h_addr ? ram_442 : _GEN_18975; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18977 = 10'h1bb == io_h_addr ? ram_443 : _GEN_18976; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18978 = 10'h1bc == io_h_addr ? ram_444 : _GEN_18977; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18979 = 10'h1bd == io_h_addr ? ram_445 : _GEN_18978; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18980 = 10'h1be == io_h_addr ? ram_446 : _GEN_18979; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18981 = 10'h1bf == io_h_addr ? ram_447 : _GEN_18980; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18982 = 10'h1c0 == io_h_addr ? ram_448 : _GEN_18981; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18983 = 10'h1c1 == io_h_addr ? ram_449 : _GEN_18982; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18984 = 10'h1c2 == io_h_addr ? ram_450 : _GEN_18983; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18985 = 10'h1c3 == io_h_addr ? ram_451 : _GEN_18984; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18986 = 10'h1c4 == io_h_addr ? ram_452 : _GEN_18985; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18987 = 10'h1c5 == io_h_addr ? ram_453 : _GEN_18986; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18988 = 10'h1c6 == io_h_addr ? ram_454 : _GEN_18987; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18989 = 10'h1c7 == io_h_addr ? ram_455 : _GEN_18988; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18990 = 10'h1c8 == io_h_addr ? ram_456 : _GEN_18989; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18991 = 10'h1c9 == io_h_addr ? ram_457 : _GEN_18990; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18992 = 10'h1ca == io_h_addr ? ram_458 : _GEN_18991; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18993 = 10'h1cb == io_h_addr ? ram_459 : _GEN_18992; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18994 = 10'h1cc == io_h_addr ? ram_460 : _GEN_18993; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18995 = 10'h1cd == io_h_addr ? ram_461 : _GEN_18994; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18996 = 10'h1ce == io_h_addr ? ram_462 : _GEN_18995; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18997 = 10'h1cf == io_h_addr ? ram_463 : _GEN_18996; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18998 = 10'h1d0 == io_h_addr ? ram_464 : _GEN_18997; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_18999 = 10'h1d1 == io_h_addr ? ram_465 : _GEN_18998; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19000 = 10'h1d2 == io_h_addr ? ram_466 : _GEN_18999; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19001 = 10'h1d3 == io_h_addr ? ram_467 : _GEN_19000; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19002 = 10'h1d4 == io_h_addr ? ram_468 : _GEN_19001; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19003 = 10'h1d5 == io_h_addr ? ram_469 : _GEN_19002; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19004 = 10'h1d6 == io_h_addr ? ram_470 : _GEN_19003; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19005 = 10'h1d7 == io_h_addr ? ram_471 : _GEN_19004; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19006 = 10'h1d8 == io_h_addr ? ram_472 : _GEN_19005; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19007 = 10'h1d9 == io_h_addr ? ram_473 : _GEN_19006; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19008 = 10'h1da == io_h_addr ? ram_474 : _GEN_19007; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19009 = 10'h1db == io_h_addr ? ram_475 : _GEN_19008; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19010 = 10'h1dc == io_h_addr ? ram_476 : _GEN_19009; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19011 = 10'h1dd == io_h_addr ? ram_477 : _GEN_19010; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19012 = 10'h1de == io_h_addr ? ram_478 : _GEN_19011; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19013 = 10'h1df == io_h_addr ? ram_479 : _GEN_19012; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19014 = 10'h1e0 == io_h_addr ? ram_480 : _GEN_19013; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19015 = 10'h1e1 == io_h_addr ? ram_481 : _GEN_19014; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19016 = 10'h1e2 == io_h_addr ? ram_482 : _GEN_19015; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19017 = 10'h1e3 == io_h_addr ? ram_483 : _GEN_19016; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19018 = 10'h1e4 == io_h_addr ? ram_484 : _GEN_19017; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19019 = 10'h1e5 == io_h_addr ? ram_485 : _GEN_19018; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19020 = 10'h1e6 == io_h_addr ? ram_486 : _GEN_19019; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19021 = 10'h1e7 == io_h_addr ? ram_487 : _GEN_19020; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19022 = 10'h1e8 == io_h_addr ? ram_488 : _GEN_19021; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19023 = 10'h1e9 == io_h_addr ? ram_489 : _GEN_19022; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19024 = 10'h1ea == io_h_addr ? ram_490 : _GEN_19023; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19025 = 10'h1eb == io_h_addr ? ram_491 : _GEN_19024; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19026 = 10'h1ec == io_h_addr ? ram_492 : _GEN_19025; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19027 = 10'h1ed == io_h_addr ? ram_493 : _GEN_19026; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19028 = 10'h1ee == io_h_addr ? ram_494 : _GEN_19027; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19029 = 10'h1ef == io_h_addr ? ram_495 : _GEN_19028; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19030 = 10'h1f0 == io_h_addr ? ram_496 : _GEN_19029; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19031 = 10'h1f1 == io_h_addr ? ram_497 : _GEN_19030; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19032 = 10'h1f2 == io_h_addr ? ram_498 : _GEN_19031; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19033 = 10'h1f3 == io_h_addr ? ram_499 : _GEN_19032; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19034 = 10'h1f4 == io_h_addr ? ram_500 : _GEN_19033; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19035 = 10'h1f5 == io_h_addr ? ram_501 : _GEN_19034; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19036 = 10'h1f6 == io_h_addr ? ram_502 : _GEN_19035; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19037 = 10'h1f7 == io_h_addr ? ram_503 : _GEN_19036; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19038 = 10'h1f8 == io_h_addr ? ram_504 : _GEN_19037; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19039 = 10'h1f9 == io_h_addr ? ram_505 : _GEN_19038; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19040 = 10'h1fa == io_h_addr ? ram_506 : _GEN_19039; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19041 = 10'h1fb == io_h_addr ? ram_507 : _GEN_19040; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19042 = 10'h1fc == io_h_addr ? ram_508 : _GEN_19041; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19043 = 10'h1fd == io_h_addr ? ram_509 : _GEN_19042; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19044 = 10'h1fe == io_h_addr ? ram_510 : _GEN_19043; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19045 = 10'h1ff == io_h_addr ? ram_511 : _GEN_19044; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19046 = 10'h200 == io_h_addr ? ram_512 : _GEN_19045; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19047 = 10'h201 == io_h_addr ? ram_513 : _GEN_19046; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19048 = 10'h202 == io_h_addr ? ram_514 : _GEN_19047; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19049 = 10'h203 == io_h_addr ? ram_515 : _GEN_19048; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19050 = 10'h204 == io_h_addr ? ram_516 : _GEN_19049; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19051 = 10'h205 == io_h_addr ? ram_517 : _GEN_19050; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19052 = 10'h206 == io_h_addr ? ram_518 : _GEN_19051; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19053 = 10'h207 == io_h_addr ? ram_519 : _GEN_19052; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19054 = 10'h208 == io_h_addr ? ram_520 : _GEN_19053; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19055 = 10'h209 == io_h_addr ? ram_521 : _GEN_19054; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19056 = 10'h20a == io_h_addr ? ram_522 : _GEN_19055; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19057 = 10'h20b == io_h_addr ? ram_523 : _GEN_19056; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _GEN_19058 = 10'h20c == io_h_addr ? ram_524 : _GEN_19057; // @[vga.scala 69:24 vga.scala 69:24]
  wire [287:0] _T_40 = _GEN_19058 >> io_v_addr; // @[vga.scala 69:24]
  assign vga_mem_ram_MPORT_addr = vga_mem_ram_MPORT_addr_pipe_0;
  assign vga_mem_ram_MPORT_data = vga_mem[vga_mem_ram_MPORT_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_1_addr = vga_mem_ram_MPORT_1_addr_pipe_0;
  assign vga_mem_ram_MPORT_1_data = vga_mem[vga_mem_ram_MPORT_1_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_2_addr = vga_mem_ram_MPORT_2_addr_pipe_0;
  assign vga_mem_ram_MPORT_2_data = vga_mem[vga_mem_ram_MPORT_2_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_3_addr = vga_mem_ram_MPORT_3_addr_pipe_0;
  assign vga_mem_ram_MPORT_3_data = vga_mem[vga_mem_ram_MPORT_3_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_4_addr = vga_mem_ram_MPORT_4_addr_pipe_0;
  assign vga_mem_ram_MPORT_4_data = vga_mem[vga_mem_ram_MPORT_4_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_5_addr = vga_mem_ram_MPORT_5_addr_pipe_0;
  assign vga_mem_ram_MPORT_5_data = vga_mem[vga_mem_ram_MPORT_5_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_6_addr = vga_mem_ram_MPORT_6_addr_pipe_0;
  assign vga_mem_ram_MPORT_6_data = vga_mem[vga_mem_ram_MPORT_6_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_7_addr = vga_mem_ram_MPORT_7_addr_pipe_0;
  assign vga_mem_ram_MPORT_7_data = vga_mem[vga_mem_ram_MPORT_7_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_8_addr = vga_mem_ram_MPORT_8_addr_pipe_0;
  assign vga_mem_ram_MPORT_8_data = vga_mem[vga_mem_ram_MPORT_8_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_9_addr = vga_mem_ram_MPORT_9_addr_pipe_0;
  assign vga_mem_ram_MPORT_9_data = vga_mem[vga_mem_ram_MPORT_9_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_10_addr = vga_mem_ram_MPORT_10_addr_pipe_0;
  assign vga_mem_ram_MPORT_10_data = vga_mem[vga_mem_ram_MPORT_10_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_11_addr = vga_mem_ram_MPORT_11_addr_pipe_0;
  assign vga_mem_ram_MPORT_11_data = vga_mem[vga_mem_ram_MPORT_11_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_12_addr = vga_mem_ram_MPORT_12_addr_pipe_0;
  assign vga_mem_ram_MPORT_12_data = vga_mem[vga_mem_ram_MPORT_12_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_13_addr = vga_mem_ram_MPORT_13_addr_pipe_0;
  assign vga_mem_ram_MPORT_13_data = vga_mem[vga_mem_ram_MPORT_13_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_14_addr = vga_mem_ram_MPORT_14_addr_pipe_0;
  assign vga_mem_ram_MPORT_14_data = vga_mem[vga_mem_ram_MPORT_14_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_15_addr = vga_mem_ram_MPORT_15_addr_pipe_0;
  assign vga_mem_ram_MPORT_15_data = vga_mem[vga_mem_ram_MPORT_15_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_16_addr = vga_mem_ram_MPORT_16_addr_pipe_0;
  assign vga_mem_ram_MPORT_16_data = vga_mem[vga_mem_ram_MPORT_16_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_17_addr = vga_mem_ram_MPORT_17_addr_pipe_0;
  assign vga_mem_ram_MPORT_17_data = vga_mem[vga_mem_ram_MPORT_17_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_18_addr = vga_mem_ram_MPORT_18_addr_pipe_0;
  assign vga_mem_ram_MPORT_18_data = vga_mem[vga_mem_ram_MPORT_18_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_19_addr = vga_mem_ram_MPORT_19_addr_pipe_0;
  assign vga_mem_ram_MPORT_19_data = vga_mem[vga_mem_ram_MPORT_19_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_20_addr = vga_mem_ram_MPORT_20_addr_pipe_0;
  assign vga_mem_ram_MPORT_20_data = vga_mem[vga_mem_ram_MPORT_20_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_21_addr = vga_mem_ram_MPORT_21_addr_pipe_0;
  assign vga_mem_ram_MPORT_21_data = vga_mem[vga_mem_ram_MPORT_21_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_22_addr = vga_mem_ram_MPORT_22_addr_pipe_0;
  assign vga_mem_ram_MPORT_22_data = vga_mem[vga_mem_ram_MPORT_22_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_23_addr = vga_mem_ram_MPORT_23_addr_pipe_0;
  assign vga_mem_ram_MPORT_23_data = vga_mem[vga_mem_ram_MPORT_23_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_24_addr = vga_mem_ram_MPORT_24_addr_pipe_0;
  assign vga_mem_ram_MPORT_24_data = vga_mem[vga_mem_ram_MPORT_24_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_25_addr = vga_mem_ram_MPORT_25_addr_pipe_0;
  assign vga_mem_ram_MPORT_25_data = vga_mem[vga_mem_ram_MPORT_25_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_26_addr = vga_mem_ram_MPORT_26_addr_pipe_0;
  assign vga_mem_ram_MPORT_26_data = vga_mem[vga_mem_ram_MPORT_26_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_27_addr = vga_mem_ram_MPORT_27_addr_pipe_0;
  assign vga_mem_ram_MPORT_27_data = vga_mem[vga_mem_ram_MPORT_27_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_28_addr = vga_mem_ram_MPORT_28_addr_pipe_0;
  assign vga_mem_ram_MPORT_28_data = vga_mem[vga_mem_ram_MPORT_28_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_29_addr = vga_mem_ram_MPORT_29_addr_pipe_0;
  assign vga_mem_ram_MPORT_29_data = vga_mem[vga_mem_ram_MPORT_29_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_30_addr = vga_mem_ram_MPORT_30_addr_pipe_0;
  assign vga_mem_ram_MPORT_30_data = vga_mem[vga_mem_ram_MPORT_30_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_31_addr = vga_mem_ram_MPORT_31_addr_pipe_0;
  assign vga_mem_ram_MPORT_31_data = vga_mem[vga_mem_ram_MPORT_31_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_32_addr = vga_mem_ram_MPORT_32_addr_pipe_0;
  assign vga_mem_ram_MPORT_32_data = vga_mem[vga_mem_ram_MPORT_32_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_33_addr = vga_mem_ram_MPORT_33_addr_pipe_0;
  assign vga_mem_ram_MPORT_33_data = vga_mem[vga_mem_ram_MPORT_33_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_34_addr = vga_mem_ram_MPORT_34_addr_pipe_0;
  assign vga_mem_ram_MPORT_34_data = vga_mem[vga_mem_ram_MPORT_34_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_35_addr = vga_mem_ram_MPORT_35_addr_pipe_0;
  assign vga_mem_ram_MPORT_35_data = vga_mem[vga_mem_ram_MPORT_35_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_36_addr = vga_mem_ram_MPORT_36_addr_pipe_0;
  assign vga_mem_ram_MPORT_36_data = vga_mem[vga_mem_ram_MPORT_36_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_37_addr = vga_mem_ram_MPORT_37_addr_pipe_0;
  assign vga_mem_ram_MPORT_37_data = vga_mem[vga_mem_ram_MPORT_37_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_38_addr = vga_mem_ram_MPORT_38_addr_pipe_0;
  assign vga_mem_ram_MPORT_38_data = vga_mem[vga_mem_ram_MPORT_38_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_39_addr = vga_mem_ram_MPORT_39_addr_pipe_0;
  assign vga_mem_ram_MPORT_39_data = vga_mem[vga_mem_ram_MPORT_39_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_40_addr = vga_mem_ram_MPORT_40_addr_pipe_0;
  assign vga_mem_ram_MPORT_40_data = vga_mem[vga_mem_ram_MPORT_40_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_41_addr = vga_mem_ram_MPORT_41_addr_pipe_0;
  assign vga_mem_ram_MPORT_41_data = vga_mem[vga_mem_ram_MPORT_41_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_42_addr = vga_mem_ram_MPORT_42_addr_pipe_0;
  assign vga_mem_ram_MPORT_42_data = vga_mem[vga_mem_ram_MPORT_42_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_43_addr = vga_mem_ram_MPORT_43_addr_pipe_0;
  assign vga_mem_ram_MPORT_43_data = vga_mem[vga_mem_ram_MPORT_43_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_44_addr = vga_mem_ram_MPORT_44_addr_pipe_0;
  assign vga_mem_ram_MPORT_44_data = vga_mem[vga_mem_ram_MPORT_44_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_45_addr = vga_mem_ram_MPORT_45_addr_pipe_0;
  assign vga_mem_ram_MPORT_45_data = vga_mem[vga_mem_ram_MPORT_45_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_46_addr = vga_mem_ram_MPORT_46_addr_pipe_0;
  assign vga_mem_ram_MPORT_46_data = vga_mem[vga_mem_ram_MPORT_46_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_47_addr = vga_mem_ram_MPORT_47_addr_pipe_0;
  assign vga_mem_ram_MPORT_47_data = vga_mem[vga_mem_ram_MPORT_47_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_48_addr = vga_mem_ram_MPORT_48_addr_pipe_0;
  assign vga_mem_ram_MPORT_48_data = vga_mem[vga_mem_ram_MPORT_48_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_49_addr = vga_mem_ram_MPORT_49_addr_pipe_0;
  assign vga_mem_ram_MPORT_49_data = vga_mem[vga_mem_ram_MPORT_49_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_50_addr = vga_mem_ram_MPORT_50_addr_pipe_0;
  assign vga_mem_ram_MPORT_50_data = vga_mem[vga_mem_ram_MPORT_50_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_51_addr = vga_mem_ram_MPORT_51_addr_pipe_0;
  assign vga_mem_ram_MPORT_51_data = vga_mem[vga_mem_ram_MPORT_51_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_52_addr = vga_mem_ram_MPORT_52_addr_pipe_0;
  assign vga_mem_ram_MPORT_52_data = vga_mem[vga_mem_ram_MPORT_52_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_53_addr = vga_mem_ram_MPORT_53_addr_pipe_0;
  assign vga_mem_ram_MPORT_53_data = vga_mem[vga_mem_ram_MPORT_53_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_54_addr = vga_mem_ram_MPORT_54_addr_pipe_0;
  assign vga_mem_ram_MPORT_54_data = vga_mem[vga_mem_ram_MPORT_54_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_55_addr = vga_mem_ram_MPORT_55_addr_pipe_0;
  assign vga_mem_ram_MPORT_55_data = vga_mem[vga_mem_ram_MPORT_55_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_56_addr = vga_mem_ram_MPORT_56_addr_pipe_0;
  assign vga_mem_ram_MPORT_56_data = vga_mem[vga_mem_ram_MPORT_56_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_57_addr = vga_mem_ram_MPORT_57_addr_pipe_0;
  assign vga_mem_ram_MPORT_57_data = vga_mem[vga_mem_ram_MPORT_57_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_58_addr = vga_mem_ram_MPORT_58_addr_pipe_0;
  assign vga_mem_ram_MPORT_58_data = vga_mem[vga_mem_ram_MPORT_58_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_59_addr = vga_mem_ram_MPORT_59_addr_pipe_0;
  assign vga_mem_ram_MPORT_59_data = vga_mem[vga_mem_ram_MPORT_59_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_60_addr = vga_mem_ram_MPORT_60_addr_pipe_0;
  assign vga_mem_ram_MPORT_60_data = vga_mem[vga_mem_ram_MPORT_60_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_61_addr = vga_mem_ram_MPORT_61_addr_pipe_0;
  assign vga_mem_ram_MPORT_61_data = vga_mem[vga_mem_ram_MPORT_61_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_62_addr = vga_mem_ram_MPORT_62_addr_pipe_0;
  assign vga_mem_ram_MPORT_62_data = vga_mem[vga_mem_ram_MPORT_62_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_63_addr = vga_mem_ram_MPORT_63_addr_pipe_0;
  assign vga_mem_ram_MPORT_63_data = vga_mem[vga_mem_ram_MPORT_63_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_64_addr = vga_mem_ram_MPORT_64_addr_pipe_0;
  assign vga_mem_ram_MPORT_64_data = vga_mem[vga_mem_ram_MPORT_64_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_65_addr = vga_mem_ram_MPORT_65_addr_pipe_0;
  assign vga_mem_ram_MPORT_65_data = vga_mem[vga_mem_ram_MPORT_65_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_66_addr = vga_mem_ram_MPORT_66_addr_pipe_0;
  assign vga_mem_ram_MPORT_66_data = vga_mem[vga_mem_ram_MPORT_66_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_67_addr = vga_mem_ram_MPORT_67_addr_pipe_0;
  assign vga_mem_ram_MPORT_67_data = vga_mem[vga_mem_ram_MPORT_67_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_68_addr = vga_mem_ram_MPORT_68_addr_pipe_0;
  assign vga_mem_ram_MPORT_68_data = vga_mem[vga_mem_ram_MPORT_68_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_69_addr = vga_mem_ram_MPORT_69_addr_pipe_0;
  assign vga_mem_ram_MPORT_69_data = vga_mem[vga_mem_ram_MPORT_69_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_70_addr = vga_mem_ram_MPORT_70_addr_pipe_0;
  assign vga_mem_ram_MPORT_70_data = vga_mem[vga_mem_ram_MPORT_70_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_71_addr = vga_mem_ram_MPORT_71_addr_pipe_0;
  assign vga_mem_ram_MPORT_71_data = vga_mem[vga_mem_ram_MPORT_71_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_72_addr = vga_mem_ram_MPORT_72_addr_pipe_0;
  assign vga_mem_ram_MPORT_72_data = vga_mem[vga_mem_ram_MPORT_72_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_73_addr = vga_mem_ram_MPORT_73_addr_pipe_0;
  assign vga_mem_ram_MPORT_73_data = vga_mem[vga_mem_ram_MPORT_73_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_74_addr = vga_mem_ram_MPORT_74_addr_pipe_0;
  assign vga_mem_ram_MPORT_74_data = vga_mem[vga_mem_ram_MPORT_74_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_75_addr = vga_mem_ram_MPORT_75_addr_pipe_0;
  assign vga_mem_ram_MPORT_75_data = vga_mem[vga_mem_ram_MPORT_75_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_76_addr = vga_mem_ram_MPORT_76_addr_pipe_0;
  assign vga_mem_ram_MPORT_76_data = vga_mem[vga_mem_ram_MPORT_76_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_77_addr = vga_mem_ram_MPORT_77_addr_pipe_0;
  assign vga_mem_ram_MPORT_77_data = vga_mem[vga_mem_ram_MPORT_77_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_78_addr = vga_mem_ram_MPORT_78_addr_pipe_0;
  assign vga_mem_ram_MPORT_78_data = vga_mem[vga_mem_ram_MPORT_78_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_79_addr = vga_mem_ram_MPORT_79_addr_pipe_0;
  assign vga_mem_ram_MPORT_79_data = vga_mem[vga_mem_ram_MPORT_79_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_80_addr = vga_mem_ram_MPORT_80_addr_pipe_0;
  assign vga_mem_ram_MPORT_80_data = vga_mem[vga_mem_ram_MPORT_80_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_81_addr = vga_mem_ram_MPORT_81_addr_pipe_0;
  assign vga_mem_ram_MPORT_81_data = vga_mem[vga_mem_ram_MPORT_81_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_82_addr = vga_mem_ram_MPORT_82_addr_pipe_0;
  assign vga_mem_ram_MPORT_82_data = vga_mem[vga_mem_ram_MPORT_82_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_83_addr = vga_mem_ram_MPORT_83_addr_pipe_0;
  assign vga_mem_ram_MPORT_83_data = vga_mem[vga_mem_ram_MPORT_83_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_84_addr = vga_mem_ram_MPORT_84_addr_pipe_0;
  assign vga_mem_ram_MPORT_84_data = vga_mem[vga_mem_ram_MPORT_84_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_85_addr = vga_mem_ram_MPORT_85_addr_pipe_0;
  assign vga_mem_ram_MPORT_85_data = vga_mem[vga_mem_ram_MPORT_85_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_86_addr = vga_mem_ram_MPORT_86_addr_pipe_0;
  assign vga_mem_ram_MPORT_86_data = vga_mem[vga_mem_ram_MPORT_86_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_87_addr = vga_mem_ram_MPORT_87_addr_pipe_0;
  assign vga_mem_ram_MPORT_87_data = vga_mem[vga_mem_ram_MPORT_87_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_88_addr = vga_mem_ram_MPORT_88_addr_pipe_0;
  assign vga_mem_ram_MPORT_88_data = vga_mem[vga_mem_ram_MPORT_88_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_89_addr = vga_mem_ram_MPORT_89_addr_pipe_0;
  assign vga_mem_ram_MPORT_89_data = vga_mem[vga_mem_ram_MPORT_89_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_90_addr = vga_mem_ram_MPORT_90_addr_pipe_0;
  assign vga_mem_ram_MPORT_90_data = vga_mem[vga_mem_ram_MPORT_90_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_91_addr = vga_mem_ram_MPORT_91_addr_pipe_0;
  assign vga_mem_ram_MPORT_91_data = vga_mem[vga_mem_ram_MPORT_91_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_92_addr = vga_mem_ram_MPORT_92_addr_pipe_0;
  assign vga_mem_ram_MPORT_92_data = vga_mem[vga_mem_ram_MPORT_92_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_93_addr = vga_mem_ram_MPORT_93_addr_pipe_0;
  assign vga_mem_ram_MPORT_93_data = vga_mem[vga_mem_ram_MPORT_93_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_94_addr = vga_mem_ram_MPORT_94_addr_pipe_0;
  assign vga_mem_ram_MPORT_94_data = vga_mem[vga_mem_ram_MPORT_94_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_95_addr = vga_mem_ram_MPORT_95_addr_pipe_0;
  assign vga_mem_ram_MPORT_95_data = vga_mem[vga_mem_ram_MPORT_95_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_96_addr = vga_mem_ram_MPORT_96_addr_pipe_0;
  assign vga_mem_ram_MPORT_96_data = vga_mem[vga_mem_ram_MPORT_96_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_97_addr = vga_mem_ram_MPORT_97_addr_pipe_0;
  assign vga_mem_ram_MPORT_97_data = vga_mem[vga_mem_ram_MPORT_97_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_98_addr = vga_mem_ram_MPORT_98_addr_pipe_0;
  assign vga_mem_ram_MPORT_98_data = vga_mem[vga_mem_ram_MPORT_98_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_99_addr = vga_mem_ram_MPORT_99_addr_pipe_0;
  assign vga_mem_ram_MPORT_99_data = vga_mem[vga_mem_ram_MPORT_99_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_100_addr = vga_mem_ram_MPORT_100_addr_pipe_0;
  assign vga_mem_ram_MPORT_100_data = vga_mem[vga_mem_ram_MPORT_100_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_101_addr = vga_mem_ram_MPORT_101_addr_pipe_0;
  assign vga_mem_ram_MPORT_101_data = vga_mem[vga_mem_ram_MPORT_101_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_102_addr = vga_mem_ram_MPORT_102_addr_pipe_0;
  assign vga_mem_ram_MPORT_102_data = vga_mem[vga_mem_ram_MPORT_102_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_103_addr = vga_mem_ram_MPORT_103_addr_pipe_0;
  assign vga_mem_ram_MPORT_103_data = vga_mem[vga_mem_ram_MPORT_103_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_104_addr = vga_mem_ram_MPORT_104_addr_pipe_0;
  assign vga_mem_ram_MPORT_104_data = vga_mem[vga_mem_ram_MPORT_104_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_105_addr = vga_mem_ram_MPORT_105_addr_pipe_0;
  assign vga_mem_ram_MPORT_105_data = vga_mem[vga_mem_ram_MPORT_105_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_106_addr = vga_mem_ram_MPORT_106_addr_pipe_0;
  assign vga_mem_ram_MPORT_106_data = vga_mem[vga_mem_ram_MPORT_106_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_107_addr = vga_mem_ram_MPORT_107_addr_pipe_0;
  assign vga_mem_ram_MPORT_107_data = vga_mem[vga_mem_ram_MPORT_107_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_108_addr = vga_mem_ram_MPORT_108_addr_pipe_0;
  assign vga_mem_ram_MPORT_108_data = vga_mem[vga_mem_ram_MPORT_108_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_109_addr = vga_mem_ram_MPORT_109_addr_pipe_0;
  assign vga_mem_ram_MPORT_109_data = vga_mem[vga_mem_ram_MPORT_109_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_110_addr = vga_mem_ram_MPORT_110_addr_pipe_0;
  assign vga_mem_ram_MPORT_110_data = vga_mem[vga_mem_ram_MPORT_110_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_111_addr = vga_mem_ram_MPORT_111_addr_pipe_0;
  assign vga_mem_ram_MPORT_111_data = vga_mem[vga_mem_ram_MPORT_111_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_112_addr = vga_mem_ram_MPORT_112_addr_pipe_0;
  assign vga_mem_ram_MPORT_112_data = vga_mem[vga_mem_ram_MPORT_112_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_113_addr = vga_mem_ram_MPORT_113_addr_pipe_0;
  assign vga_mem_ram_MPORT_113_data = vga_mem[vga_mem_ram_MPORT_113_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_114_addr = vga_mem_ram_MPORT_114_addr_pipe_0;
  assign vga_mem_ram_MPORT_114_data = vga_mem[vga_mem_ram_MPORT_114_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_115_addr = vga_mem_ram_MPORT_115_addr_pipe_0;
  assign vga_mem_ram_MPORT_115_data = vga_mem[vga_mem_ram_MPORT_115_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_116_addr = vga_mem_ram_MPORT_116_addr_pipe_0;
  assign vga_mem_ram_MPORT_116_data = vga_mem[vga_mem_ram_MPORT_116_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_117_addr = vga_mem_ram_MPORT_117_addr_pipe_0;
  assign vga_mem_ram_MPORT_117_data = vga_mem[vga_mem_ram_MPORT_117_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_118_addr = vga_mem_ram_MPORT_118_addr_pipe_0;
  assign vga_mem_ram_MPORT_118_data = vga_mem[vga_mem_ram_MPORT_118_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_119_addr = vga_mem_ram_MPORT_119_addr_pipe_0;
  assign vga_mem_ram_MPORT_119_data = vga_mem[vga_mem_ram_MPORT_119_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_120_addr = vga_mem_ram_MPORT_120_addr_pipe_0;
  assign vga_mem_ram_MPORT_120_data = vga_mem[vga_mem_ram_MPORT_120_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_121_addr = vga_mem_ram_MPORT_121_addr_pipe_0;
  assign vga_mem_ram_MPORT_121_data = vga_mem[vga_mem_ram_MPORT_121_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_122_addr = vga_mem_ram_MPORT_122_addr_pipe_0;
  assign vga_mem_ram_MPORT_122_data = vga_mem[vga_mem_ram_MPORT_122_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_123_addr = vga_mem_ram_MPORT_123_addr_pipe_0;
  assign vga_mem_ram_MPORT_123_data = vga_mem[vga_mem_ram_MPORT_123_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_124_addr = vga_mem_ram_MPORT_124_addr_pipe_0;
  assign vga_mem_ram_MPORT_124_data = vga_mem[vga_mem_ram_MPORT_124_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_125_addr = vga_mem_ram_MPORT_125_addr_pipe_0;
  assign vga_mem_ram_MPORT_125_data = vga_mem[vga_mem_ram_MPORT_125_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_126_addr = vga_mem_ram_MPORT_126_addr_pipe_0;
  assign vga_mem_ram_MPORT_126_data = vga_mem[vga_mem_ram_MPORT_126_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_127_addr = vga_mem_ram_MPORT_127_addr_pipe_0;
  assign vga_mem_ram_MPORT_127_data = vga_mem[vga_mem_ram_MPORT_127_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_128_addr = vga_mem_ram_MPORT_128_addr_pipe_0;
  assign vga_mem_ram_MPORT_128_data = vga_mem[vga_mem_ram_MPORT_128_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_129_addr = vga_mem_ram_MPORT_129_addr_pipe_0;
  assign vga_mem_ram_MPORT_129_data = vga_mem[vga_mem_ram_MPORT_129_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_130_addr = vga_mem_ram_MPORT_130_addr_pipe_0;
  assign vga_mem_ram_MPORT_130_data = vga_mem[vga_mem_ram_MPORT_130_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_131_addr = vga_mem_ram_MPORT_131_addr_pipe_0;
  assign vga_mem_ram_MPORT_131_data = vga_mem[vga_mem_ram_MPORT_131_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_132_addr = vga_mem_ram_MPORT_132_addr_pipe_0;
  assign vga_mem_ram_MPORT_132_data = vga_mem[vga_mem_ram_MPORT_132_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_133_addr = vga_mem_ram_MPORT_133_addr_pipe_0;
  assign vga_mem_ram_MPORT_133_data = vga_mem[vga_mem_ram_MPORT_133_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_134_addr = vga_mem_ram_MPORT_134_addr_pipe_0;
  assign vga_mem_ram_MPORT_134_data = vga_mem[vga_mem_ram_MPORT_134_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_135_addr = vga_mem_ram_MPORT_135_addr_pipe_0;
  assign vga_mem_ram_MPORT_135_data = vga_mem[vga_mem_ram_MPORT_135_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_136_addr = vga_mem_ram_MPORT_136_addr_pipe_0;
  assign vga_mem_ram_MPORT_136_data = vga_mem[vga_mem_ram_MPORT_136_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_137_addr = vga_mem_ram_MPORT_137_addr_pipe_0;
  assign vga_mem_ram_MPORT_137_data = vga_mem[vga_mem_ram_MPORT_137_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_138_addr = vga_mem_ram_MPORT_138_addr_pipe_0;
  assign vga_mem_ram_MPORT_138_data = vga_mem[vga_mem_ram_MPORT_138_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_139_addr = vga_mem_ram_MPORT_139_addr_pipe_0;
  assign vga_mem_ram_MPORT_139_data = vga_mem[vga_mem_ram_MPORT_139_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_140_addr = vga_mem_ram_MPORT_140_addr_pipe_0;
  assign vga_mem_ram_MPORT_140_data = vga_mem[vga_mem_ram_MPORT_140_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_141_addr = vga_mem_ram_MPORT_141_addr_pipe_0;
  assign vga_mem_ram_MPORT_141_data = vga_mem[vga_mem_ram_MPORT_141_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_142_addr = vga_mem_ram_MPORT_142_addr_pipe_0;
  assign vga_mem_ram_MPORT_142_data = vga_mem[vga_mem_ram_MPORT_142_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_143_addr = vga_mem_ram_MPORT_143_addr_pipe_0;
  assign vga_mem_ram_MPORT_143_data = vga_mem[vga_mem_ram_MPORT_143_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_144_addr = vga_mem_ram_MPORT_144_addr_pipe_0;
  assign vga_mem_ram_MPORT_144_data = vga_mem[vga_mem_ram_MPORT_144_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_145_addr = vga_mem_ram_MPORT_145_addr_pipe_0;
  assign vga_mem_ram_MPORT_145_data = vga_mem[vga_mem_ram_MPORT_145_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_146_addr = vga_mem_ram_MPORT_146_addr_pipe_0;
  assign vga_mem_ram_MPORT_146_data = vga_mem[vga_mem_ram_MPORT_146_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_147_addr = vga_mem_ram_MPORT_147_addr_pipe_0;
  assign vga_mem_ram_MPORT_147_data = vga_mem[vga_mem_ram_MPORT_147_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_148_addr = vga_mem_ram_MPORT_148_addr_pipe_0;
  assign vga_mem_ram_MPORT_148_data = vga_mem[vga_mem_ram_MPORT_148_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_149_addr = vga_mem_ram_MPORT_149_addr_pipe_0;
  assign vga_mem_ram_MPORT_149_data = vga_mem[vga_mem_ram_MPORT_149_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_150_addr = vga_mem_ram_MPORT_150_addr_pipe_0;
  assign vga_mem_ram_MPORT_150_data = vga_mem[vga_mem_ram_MPORT_150_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_151_addr = vga_mem_ram_MPORT_151_addr_pipe_0;
  assign vga_mem_ram_MPORT_151_data = vga_mem[vga_mem_ram_MPORT_151_addr]; // @[vga.scala 50:30]
  assign vga_mem_ram_MPORT_152_addr = vga_mem_ram_MPORT_152_addr_pipe_0;
  assign vga_mem_ram_MPORT_152_data = vga_mem[vga_mem_ram_MPORT_152_addr]; // @[vga.scala 50:30]
  assign io_vga_data = rdwrPort; // @[vga.scala 74:16]
  always @(posedge clock) begin
    vga_mem_ram_MPORT_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_1_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_1_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_2_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_2_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_3_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_3_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_4_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_4_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_5_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_5_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_6_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_6_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_7_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_7_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_8_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_8_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_9_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_9_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_10_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_10_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_11_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_11_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_12_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_12_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_13_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_13_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_14_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_14_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_15_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_15_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_16_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_16_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_17_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_17_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_18_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_18_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_19_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_19_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_20_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_20_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_21_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_21_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_22_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_22_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_23_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_23_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_24_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_24_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_25_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_25_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_26_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_26_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_27_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_27_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_28_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_28_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_29_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_29_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_30_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_30_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_31_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_31_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_32_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_32_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_33_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_33_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_34_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_34_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_35_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_35_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_36_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_36_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_37_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_37_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_38_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_38_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_39_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_39_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_40_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_40_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_41_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_41_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_42_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_42_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_43_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_43_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_44_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_44_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_45_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_45_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_46_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_46_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_47_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_47_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_48_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_48_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_49_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_49_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_50_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_50_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_51_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_51_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_52_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_52_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_53_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_53_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_54_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_54_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_55_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_55_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_56_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_56_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_57_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_57_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_58_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_58_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_59_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_59_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_60_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_60_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_61_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_61_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_62_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_62_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_63_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_63_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_64_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_64_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_65_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_65_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_66_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_66_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_67_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_67_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_68_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_68_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_69_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_69_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_70_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_70_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_71_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_71_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_72_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_72_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_73_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_73_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_74_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_74_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_75_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_75_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_76_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_76_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_77_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_77_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_78_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_78_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_79_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_79_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_80_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_80_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_81_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_81_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_82_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_82_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_83_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_83_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_84_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_84_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_85_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_85_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_86_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_86_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_87_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_87_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_88_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_88_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_89_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_89_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_90_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_90_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_91_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_91_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_92_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_92_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_93_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_93_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_94_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_94_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_95_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_95_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_96_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_96_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_97_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_97_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_98_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_98_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_99_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_99_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_100_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_100_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_101_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_101_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_102_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_102_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_103_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_103_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_104_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_104_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_105_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_105_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_106_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_106_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_107_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_107_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_108_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_108_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_109_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_109_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_110_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_110_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_111_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_111_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_112_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_112_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_113_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_113_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_114_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_114_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_115_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_115_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_116_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_116_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_117_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_117_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_118_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_118_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_119_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_119_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_120_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_120_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_121_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_121_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_122_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_122_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_123_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_123_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_124_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_124_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_125_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_125_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_126_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_126_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_127_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_127_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_128_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_128_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_129_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_129_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_130_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_130_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_131_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_131_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_132_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_132_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_133_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_133_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_134_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_134_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_135_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_135_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_136_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_136_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_137_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_137_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_138_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_138_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_139_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_139_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_140_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_140_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_141_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_141_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_142_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_142_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_143_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_143_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_144_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_144_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_145_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_145_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_146_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_146_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_147_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_147_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_148_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_148_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_149_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_149_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_150_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_150_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_151_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_151_addr_pipe_0 <= _ram_T_2[11:0];
    end
    vga_mem_ram_MPORT_152_en_pipe_0 <= io_now != 2'h0;
    if (io_now != 2'h0) begin
      vga_mem_ram_MPORT_152_addr_pipe_0 <= _ram_T_2[11:0];
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_0 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_0 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h0 == _T_37) begin // @[vga.scala 64:24]
        ram_0 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_0 <= _GEN_15228;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_1 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_1 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1 == _T_37) begin // @[vga.scala 64:24]
        ram_1 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_1 <= _GEN_15229;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_2 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_2 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2 == _T_37) begin // @[vga.scala 64:24]
        ram_2 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_2 <= _GEN_15230;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_3 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_3 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3 == _T_37) begin // @[vga.scala 64:24]
        ram_3 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_3 <= _GEN_15231;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_4 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_4 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4 == _T_37) begin // @[vga.scala 64:24]
        ram_4 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_4 <= _GEN_15232;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_5 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_5 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5 == _T_37) begin // @[vga.scala 64:24]
        ram_5 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_5 <= _GEN_15233;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_6 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_6 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6 == _T_37) begin // @[vga.scala 64:24]
        ram_6 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_6 <= _GEN_15234;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_7 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_7 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7 == _T_37) begin // @[vga.scala 64:24]
        ram_7 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_7 <= _GEN_15235;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_8 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_8 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8 == _T_37) begin // @[vga.scala 64:24]
        ram_8 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_8 <= _GEN_15236;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_9 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_9 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9 == _T_37) begin // @[vga.scala 64:24]
        ram_9 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_9 <= _GEN_15237;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_10 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha == _h_T_1) begin // @[vga.scala 64:24]
        ram_10 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha == _T_37) begin // @[vga.scala 64:24]
        ram_10 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_10 <= _GEN_15238;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_11 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb == _h_T_1) begin // @[vga.scala 64:24]
        ram_11 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb == _T_37) begin // @[vga.scala 64:24]
        ram_11 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_11 <= _GEN_15239;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_12 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc == _h_T_1) begin // @[vga.scala 64:24]
        ram_12 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc == _T_37) begin // @[vga.scala 64:24]
        ram_12 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_12 <= _GEN_15240;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_13 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd == _h_T_1) begin // @[vga.scala 64:24]
        ram_13 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd == _T_37) begin // @[vga.scala 64:24]
        ram_13 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_13 <= _GEN_15241;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_14 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he == _h_T_1) begin // @[vga.scala 64:24]
        ram_14 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he == _T_37) begin // @[vga.scala 64:24]
        ram_14 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_14 <= _GEN_15242;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_15 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf == _h_T_1) begin // @[vga.scala 64:24]
        ram_15 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf == _T_37) begin // @[vga.scala 64:24]
        ram_15 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_15 <= _GEN_15243;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_16 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10 == _h_T_1) begin // @[vga.scala 64:24]
        ram_16 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10 == _T_37) begin // @[vga.scala 64:24]
        ram_16 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_16 <= _GEN_15244;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_17 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11 == _h_T_1) begin // @[vga.scala 64:24]
        ram_17 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11 == _T_37) begin // @[vga.scala 64:24]
        ram_17 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_17 <= _GEN_15245;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_18 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12 == _h_T_1) begin // @[vga.scala 64:24]
        ram_18 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12 == _T_37) begin // @[vga.scala 64:24]
        ram_18 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_18 <= _GEN_15246;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_19 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13 == _h_T_1) begin // @[vga.scala 64:24]
        ram_19 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13 == _T_37) begin // @[vga.scala 64:24]
        ram_19 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_19 <= _GEN_15247;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_20 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14 == _h_T_1) begin // @[vga.scala 64:24]
        ram_20 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14 == _T_37) begin // @[vga.scala 64:24]
        ram_20 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_20 <= _GEN_15248;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_21 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15 == _h_T_1) begin // @[vga.scala 64:24]
        ram_21 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15 == _T_37) begin // @[vga.scala 64:24]
        ram_21 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_21 <= _GEN_15249;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_22 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16 == _h_T_1) begin // @[vga.scala 64:24]
        ram_22 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16 == _T_37) begin // @[vga.scala 64:24]
        ram_22 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_22 <= _GEN_15250;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_23 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17 == _h_T_1) begin // @[vga.scala 64:24]
        ram_23 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17 == _T_37) begin // @[vga.scala 64:24]
        ram_23 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_23 <= _GEN_15251;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_24 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18 == _h_T_1) begin // @[vga.scala 64:24]
        ram_24 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18 == _T_37) begin // @[vga.scala 64:24]
        ram_24 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_24 <= _GEN_15252;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_25 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19 == _h_T_1) begin // @[vga.scala 64:24]
        ram_25 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19 == _T_37) begin // @[vga.scala 64:24]
        ram_25 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_25 <= _GEN_15253;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_26 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a == _h_T_1) begin // @[vga.scala 64:24]
        ram_26 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a == _T_37) begin // @[vga.scala 64:24]
        ram_26 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_26 <= _GEN_15254;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_27 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b == _h_T_1) begin // @[vga.scala 64:24]
        ram_27 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b == _T_37) begin // @[vga.scala 64:24]
        ram_27 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_27 <= _GEN_15255;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_28 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c == _h_T_1) begin // @[vga.scala 64:24]
        ram_28 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c == _T_37) begin // @[vga.scala 64:24]
        ram_28 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_28 <= _GEN_15256;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_29 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d == _h_T_1) begin // @[vga.scala 64:24]
        ram_29 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d == _T_37) begin // @[vga.scala 64:24]
        ram_29 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_29 <= _GEN_15257;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_30 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e == _h_T_1) begin // @[vga.scala 64:24]
        ram_30 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e == _T_37) begin // @[vga.scala 64:24]
        ram_30 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_30 <= _GEN_15258;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_31 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f == _h_T_1) begin // @[vga.scala 64:24]
        ram_31 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f == _T_37) begin // @[vga.scala 64:24]
        ram_31 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_31 <= _GEN_15259;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_32 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h20 == _h_T_1) begin // @[vga.scala 64:24]
        ram_32 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h20 == _T_37) begin // @[vga.scala 64:24]
        ram_32 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_32 <= _GEN_15260;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_33 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h21 == _h_T_1) begin // @[vga.scala 64:24]
        ram_33 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h21 == _T_37) begin // @[vga.scala 64:24]
        ram_33 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_33 <= _GEN_15261;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_34 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h22 == _h_T_1) begin // @[vga.scala 64:24]
        ram_34 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h22 == _T_37) begin // @[vga.scala 64:24]
        ram_34 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_34 <= _GEN_15262;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_35 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h23 == _h_T_1) begin // @[vga.scala 64:24]
        ram_35 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h23 == _T_37) begin // @[vga.scala 64:24]
        ram_35 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_35 <= _GEN_15263;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_36 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h24 == _h_T_1) begin // @[vga.scala 64:24]
        ram_36 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h24 == _T_37) begin // @[vga.scala 64:24]
        ram_36 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_36 <= _GEN_15264;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_37 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h25 == _h_T_1) begin // @[vga.scala 64:24]
        ram_37 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h25 == _T_37) begin // @[vga.scala 64:24]
        ram_37 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_37 <= _GEN_15265;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_38 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h26 == _h_T_1) begin // @[vga.scala 64:24]
        ram_38 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h26 == _T_37) begin // @[vga.scala 64:24]
        ram_38 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_38 <= _GEN_15266;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_39 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h27 == _h_T_1) begin // @[vga.scala 64:24]
        ram_39 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h27 == _T_37) begin // @[vga.scala 64:24]
        ram_39 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_39 <= _GEN_15267;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_40 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h28 == _h_T_1) begin // @[vga.scala 64:24]
        ram_40 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h28 == _T_37) begin // @[vga.scala 64:24]
        ram_40 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_40 <= _GEN_15268;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_41 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h29 == _h_T_1) begin // @[vga.scala 64:24]
        ram_41 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h29 == _T_37) begin // @[vga.scala 64:24]
        ram_41 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_41 <= _GEN_15269;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_42 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2a == _h_T_1) begin // @[vga.scala 64:24]
        ram_42 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2a == _T_37) begin // @[vga.scala 64:24]
        ram_42 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_42 <= _GEN_15270;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_43 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2b == _h_T_1) begin // @[vga.scala 64:24]
        ram_43 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2b == _T_37) begin // @[vga.scala 64:24]
        ram_43 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_43 <= _GEN_15271;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_44 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2c == _h_T_1) begin // @[vga.scala 64:24]
        ram_44 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2c == _T_37) begin // @[vga.scala 64:24]
        ram_44 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_44 <= _GEN_15272;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_45 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2d == _h_T_1) begin // @[vga.scala 64:24]
        ram_45 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2d == _T_37) begin // @[vga.scala 64:24]
        ram_45 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_45 <= _GEN_15273;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_46 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2e == _h_T_1) begin // @[vga.scala 64:24]
        ram_46 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2e == _T_37) begin // @[vga.scala 64:24]
        ram_46 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_46 <= _GEN_15274;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_47 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h2f == _h_T_1) begin // @[vga.scala 64:24]
        ram_47 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h2f == _T_37) begin // @[vga.scala 64:24]
        ram_47 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_47 <= _GEN_15275;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_48 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h30 == _h_T_1) begin // @[vga.scala 64:24]
        ram_48 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h30 == _T_37) begin // @[vga.scala 64:24]
        ram_48 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_48 <= _GEN_15276;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_49 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h31 == _h_T_1) begin // @[vga.scala 64:24]
        ram_49 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h31 == _T_37) begin // @[vga.scala 64:24]
        ram_49 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_49 <= _GEN_15277;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_50 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h32 == _h_T_1) begin // @[vga.scala 64:24]
        ram_50 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h32 == _T_37) begin // @[vga.scala 64:24]
        ram_50 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_50 <= _GEN_15278;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_51 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h33 == _h_T_1) begin // @[vga.scala 64:24]
        ram_51 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h33 == _T_37) begin // @[vga.scala 64:24]
        ram_51 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_51 <= _GEN_15279;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_52 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h34 == _h_T_1) begin // @[vga.scala 64:24]
        ram_52 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h34 == _T_37) begin // @[vga.scala 64:24]
        ram_52 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_52 <= _GEN_15280;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_53 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h35 == _h_T_1) begin // @[vga.scala 64:24]
        ram_53 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h35 == _T_37) begin // @[vga.scala 64:24]
        ram_53 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_53 <= _GEN_15281;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_54 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h36 == _h_T_1) begin // @[vga.scala 64:24]
        ram_54 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h36 == _T_37) begin // @[vga.scala 64:24]
        ram_54 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_54 <= _GEN_15282;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_55 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h37 == _h_T_1) begin // @[vga.scala 64:24]
        ram_55 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h37 == _T_37) begin // @[vga.scala 64:24]
        ram_55 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_55 <= _GEN_15283;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_56 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h38 == _h_T_1) begin // @[vga.scala 64:24]
        ram_56 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h38 == _T_37) begin // @[vga.scala 64:24]
        ram_56 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_56 <= _GEN_15284;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_57 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h39 == _h_T_1) begin // @[vga.scala 64:24]
        ram_57 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h39 == _T_37) begin // @[vga.scala 64:24]
        ram_57 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_57 <= _GEN_15285;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_58 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3a == _h_T_1) begin // @[vga.scala 64:24]
        ram_58 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3a == _T_37) begin // @[vga.scala 64:24]
        ram_58 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_58 <= _GEN_15286;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_59 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3b == _h_T_1) begin // @[vga.scala 64:24]
        ram_59 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3b == _T_37) begin // @[vga.scala 64:24]
        ram_59 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_59 <= _GEN_15287;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_60 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3c == _h_T_1) begin // @[vga.scala 64:24]
        ram_60 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3c == _T_37) begin // @[vga.scala 64:24]
        ram_60 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_60 <= _GEN_15288;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_61 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3d == _h_T_1) begin // @[vga.scala 64:24]
        ram_61 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3d == _T_37) begin // @[vga.scala 64:24]
        ram_61 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_61 <= _GEN_15289;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_62 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3e == _h_T_1) begin // @[vga.scala 64:24]
        ram_62 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3e == _T_37) begin // @[vga.scala 64:24]
        ram_62 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_62 <= _GEN_15290;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_63 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h3f == _h_T_1) begin // @[vga.scala 64:24]
        ram_63 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h3f == _T_37) begin // @[vga.scala 64:24]
        ram_63 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_63 <= _GEN_15291;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_64 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h40 == _h_T_1) begin // @[vga.scala 64:24]
        ram_64 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h40 == _T_37) begin // @[vga.scala 64:24]
        ram_64 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_64 <= _GEN_15292;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_65 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h41 == _h_T_1) begin // @[vga.scala 64:24]
        ram_65 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h41 == _T_37) begin // @[vga.scala 64:24]
        ram_65 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_65 <= _GEN_15293;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_66 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h42 == _h_T_1) begin // @[vga.scala 64:24]
        ram_66 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h42 == _T_37) begin // @[vga.scala 64:24]
        ram_66 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_66 <= _GEN_15294;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_67 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h43 == _h_T_1) begin // @[vga.scala 64:24]
        ram_67 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h43 == _T_37) begin // @[vga.scala 64:24]
        ram_67 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_67 <= _GEN_15295;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_68 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h44 == _h_T_1) begin // @[vga.scala 64:24]
        ram_68 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h44 == _T_37) begin // @[vga.scala 64:24]
        ram_68 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_68 <= _GEN_15296;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_69 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h45 == _h_T_1) begin // @[vga.scala 64:24]
        ram_69 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h45 == _T_37) begin // @[vga.scala 64:24]
        ram_69 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_69 <= _GEN_15297;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_70 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h46 == _h_T_1) begin // @[vga.scala 64:24]
        ram_70 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h46 == _T_37) begin // @[vga.scala 64:24]
        ram_70 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_70 <= _GEN_15298;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_71 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h47 == _h_T_1) begin // @[vga.scala 64:24]
        ram_71 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h47 == _T_37) begin // @[vga.scala 64:24]
        ram_71 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_71 <= _GEN_15299;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_72 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h48 == _h_T_1) begin // @[vga.scala 64:24]
        ram_72 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h48 == _T_37) begin // @[vga.scala 64:24]
        ram_72 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_72 <= _GEN_15300;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_73 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h49 == _h_T_1) begin // @[vga.scala 64:24]
        ram_73 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h49 == _T_37) begin // @[vga.scala 64:24]
        ram_73 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_73 <= _GEN_15301;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_74 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4a == _h_T_1) begin // @[vga.scala 64:24]
        ram_74 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4a == _T_37) begin // @[vga.scala 64:24]
        ram_74 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_74 <= _GEN_15302;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_75 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4b == _h_T_1) begin // @[vga.scala 64:24]
        ram_75 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4b == _T_37) begin // @[vga.scala 64:24]
        ram_75 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_75 <= _GEN_15303;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_76 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4c == _h_T_1) begin // @[vga.scala 64:24]
        ram_76 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4c == _T_37) begin // @[vga.scala 64:24]
        ram_76 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_76 <= _GEN_15304;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_77 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4d == _h_T_1) begin // @[vga.scala 64:24]
        ram_77 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4d == _T_37) begin // @[vga.scala 64:24]
        ram_77 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_77 <= _GEN_15305;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_78 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4e == _h_T_1) begin // @[vga.scala 64:24]
        ram_78 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4e == _T_37) begin // @[vga.scala 64:24]
        ram_78 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_78 <= _GEN_15306;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_79 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h4f == _h_T_1) begin // @[vga.scala 64:24]
        ram_79 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h4f == _T_37) begin // @[vga.scala 64:24]
        ram_79 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_79 <= _GEN_15307;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_80 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h50 == _h_T_1) begin // @[vga.scala 64:24]
        ram_80 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h50 == _T_37) begin // @[vga.scala 64:24]
        ram_80 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_80 <= _GEN_15308;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_81 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h51 == _h_T_1) begin // @[vga.scala 64:24]
        ram_81 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h51 == _T_37) begin // @[vga.scala 64:24]
        ram_81 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_81 <= _GEN_15309;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_82 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h52 == _h_T_1) begin // @[vga.scala 64:24]
        ram_82 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h52 == _T_37) begin // @[vga.scala 64:24]
        ram_82 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_82 <= _GEN_15310;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_83 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h53 == _h_T_1) begin // @[vga.scala 64:24]
        ram_83 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h53 == _T_37) begin // @[vga.scala 64:24]
        ram_83 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_83 <= _GEN_15311;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_84 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h54 == _h_T_1) begin // @[vga.scala 64:24]
        ram_84 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h54 == _T_37) begin // @[vga.scala 64:24]
        ram_84 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_84 <= _GEN_15312;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_85 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h55 == _h_T_1) begin // @[vga.scala 64:24]
        ram_85 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h55 == _T_37) begin // @[vga.scala 64:24]
        ram_85 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_85 <= _GEN_15313;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_86 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h56 == _h_T_1) begin // @[vga.scala 64:24]
        ram_86 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h56 == _T_37) begin // @[vga.scala 64:24]
        ram_86 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_86 <= _GEN_15314;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_87 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h57 == _h_T_1) begin // @[vga.scala 64:24]
        ram_87 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h57 == _T_37) begin // @[vga.scala 64:24]
        ram_87 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_87 <= _GEN_15315;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_88 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h58 == _h_T_1) begin // @[vga.scala 64:24]
        ram_88 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h58 == _T_37) begin // @[vga.scala 64:24]
        ram_88 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_88 <= _GEN_15316;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_89 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h59 == _h_T_1) begin // @[vga.scala 64:24]
        ram_89 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h59 == _T_37) begin // @[vga.scala 64:24]
        ram_89 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_89 <= _GEN_15317;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_90 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5a == _h_T_1) begin // @[vga.scala 64:24]
        ram_90 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5a == _T_37) begin // @[vga.scala 64:24]
        ram_90 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_90 <= _GEN_15318;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_91 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5b == _h_T_1) begin // @[vga.scala 64:24]
        ram_91 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5b == _T_37) begin // @[vga.scala 64:24]
        ram_91 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_91 <= _GEN_15319;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_92 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5c == _h_T_1) begin // @[vga.scala 64:24]
        ram_92 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5c == _T_37) begin // @[vga.scala 64:24]
        ram_92 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_92 <= _GEN_15320;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_93 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5d == _h_T_1) begin // @[vga.scala 64:24]
        ram_93 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5d == _T_37) begin // @[vga.scala 64:24]
        ram_93 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_93 <= _GEN_15321;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_94 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5e == _h_T_1) begin // @[vga.scala 64:24]
        ram_94 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5e == _T_37) begin // @[vga.scala 64:24]
        ram_94 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_94 <= _GEN_15322;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_95 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h5f == _h_T_1) begin // @[vga.scala 64:24]
        ram_95 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h5f == _T_37) begin // @[vga.scala 64:24]
        ram_95 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_95 <= _GEN_15323;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_96 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h60 == _h_T_1) begin // @[vga.scala 64:24]
        ram_96 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h60 == _T_37) begin // @[vga.scala 64:24]
        ram_96 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_96 <= _GEN_15324;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_97 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h61 == _h_T_1) begin // @[vga.scala 64:24]
        ram_97 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h61 == _T_37) begin // @[vga.scala 64:24]
        ram_97 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_97 <= _GEN_15325;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_98 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h62 == _h_T_1) begin // @[vga.scala 64:24]
        ram_98 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h62 == _T_37) begin // @[vga.scala 64:24]
        ram_98 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_98 <= _GEN_15326;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_99 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h63 == _h_T_1) begin // @[vga.scala 64:24]
        ram_99 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h63 == _T_37) begin // @[vga.scala 64:24]
        ram_99 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_99 <= _GEN_15327;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_100 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h64 == _h_T_1) begin // @[vga.scala 64:24]
        ram_100 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h64 == _T_37) begin // @[vga.scala 64:24]
        ram_100 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_100 <= _GEN_15328;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_101 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h65 == _h_T_1) begin // @[vga.scala 64:24]
        ram_101 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h65 == _T_37) begin // @[vga.scala 64:24]
        ram_101 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_101 <= _GEN_15329;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_102 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h66 == _h_T_1) begin // @[vga.scala 64:24]
        ram_102 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h66 == _T_37) begin // @[vga.scala 64:24]
        ram_102 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_102 <= _GEN_15330;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_103 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h67 == _h_T_1) begin // @[vga.scala 64:24]
        ram_103 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h67 == _T_37) begin // @[vga.scala 64:24]
        ram_103 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_103 <= _GEN_15331;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_104 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h68 == _h_T_1) begin // @[vga.scala 64:24]
        ram_104 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h68 == _T_37) begin // @[vga.scala 64:24]
        ram_104 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_104 <= _GEN_15332;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_105 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h69 == _h_T_1) begin // @[vga.scala 64:24]
        ram_105 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h69 == _T_37) begin // @[vga.scala 64:24]
        ram_105 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_105 <= _GEN_15333;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_106 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6a == _h_T_1) begin // @[vga.scala 64:24]
        ram_106 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6a == _T_37) begin // @[vga.scala 64:24]
        ram_106 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_106 <= _GEN_15334;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_107 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6b == _h_T_1) begin // @[vga.scala 64:24]
        ram_107 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6b == _T_37) begin // @[vga.scala 64:24]
        ram_107 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_107 <= _GEN_15335;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_108 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6c == _h_T_1) begin // @[vga.scala 64:24]
        ram_108 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6c == _T_37) begin // @[vga.scala 64:24]
        ram_108 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_108 <= _GEN_15336;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_109 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6d == _h_T_1) begin // @[vga.scala 64:24]
        ram_109 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6d == _T_37) begin // @[vga.scala 64:24]
        ram_109 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_109 <= _GEN_15337;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_110 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6e == _h_T_1) begin // @[vga.scala 64:24]
        ram_110 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6e == _T_37) begin // @[vga.scala 64:24]
        ram_110 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_110 <= _GEN_15338;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_111 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h6f == _h_T_1) begin // @[vga.scala 64:24]
        ram_111 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h6f == _T_37) begin // @[vga.scala 64:24]
        ram_111 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_111 <= _GEN_15339;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_112 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h70 == _h_T_1) begin // @[vga.scala 64:24]
        ram_112 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h70 == _T_37) begin // @[vga.scala 64:24]
        ram_112 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_112 <= _GEN_15340;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_113 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h71 == _h_T_1) begin // @[vga.scala 64:24]
        ram_113 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h71 == _T_37) begin // @[vga.scala 64:24]
        ram_113 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_113 <= _GEN_15341;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_114 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h72 == _h_T_1) begin // @[vga.scala 64:24]
        ram_114 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h72 == _T_37) begin // @[vga.scala 64:24]
        ram_114 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_114 <= _GEN_15342;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_115 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h73 == _h_T_1) begin // @[vga.scala 64:24]
        ram_115 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h73 == _T_37) begin // @[vga.scala 64:24]
        ram_115 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_115 <= _GEN_15343;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_116 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h74 == _h_T_1) begin // @[vga.scala 64:24]
        ram_116 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h74 == _T_37) begin // @[vga.scala 64:24]
        ram_116 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_116 <= _GEN_15344;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_117 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h75 == _h_T_1) begin // @[vga.scala 64:24]
        ram_117 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h75 == _T_37) begin // @[vga.scala 64:24]
        ram_117 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_117 <= _GEN_15345;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_118 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h76 == _h_T_1) begin // @[vga.scala 64:24]
        ram_118 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h76 == _T_37) begin // @[vga.scala 64:24]
        ram_118 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_118 <= _GEN_15346;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_119 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h77 == _h_T_1) begin // @[vga.scala 64:24]
        ram_119 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h77 == _T_37) begin // @[vga.scala 64:24]
        ram_119 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_119 <= _GEN_15347;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_120 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h78 == _h_T_1) begin // @[vga.scala 64:24]
        ram_120 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h78 == _T_37) begin // @[vga.scala 64:24]
        ram_120 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_120 <= _GEN_15348;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_121 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h79 == _h_T_1) begin // @[vga.scala 64:24]
        ram_121 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h79 == _T_37) begin // @[vga.scala 64:24]
        ram_121 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_121 <= _GEN_15349;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_122 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7a == _h_T_1) begin // @[vga.scala 64:24]
        ram_122 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7a == _T_37) begin // @[vga.scala 64:24]
        ram_122 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_122 <= _GEN_15350;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_123 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7b == _h_T_1) begin // @[vga.scala 64:24]
        ram_123 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7b == _T_37) begin // @[vga.scala 64:24]
        ram_123 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_123 <= _GEN_15351;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_124 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7c == _h_T_1) begin // @[vga.scala 64:24]
        ram_124 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7c == _T_37) begin // @[vga.scala 64:24]
        ram_124 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_124 <= _GEN_15352;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_125 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7d == _h_T_1) begin // @[vga.scala 64:24]
        ram_125 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7d == _T_37) begin // @[vga.scala 64:24]
        ram_125 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_125 <= _GEN_15353;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_126 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7e == _h_T_1) begin // @[vga.scala 64:24]
        ram_126 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7e == _T_37) begin // @[vga.scala 64:24]
        ram_126 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_126 <= _GEN_15354;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_127 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h7f == _h_T_1) begin // @[vga.scala 64:24]
        ram_127 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h7f == _T_37) begin // @[vga.scala 64:24]
        ram_127 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_127 <= _GEN_15355;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_128 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h80 == _h_T_1) begin // @[vga.scala 64:24]
        ram_128 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h80 == _T_37) begin // @[vga.scala 64:24]
        ram_128 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_128 <= _GEN_15356;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_129 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h81 == _h_T_1) begin // @[vga.scala 64:24]
        ram_129 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h81 == _T_37) begin // @[vga.scala 64:24]
        ram_129 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_129 <= _GEN_15357;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_130 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h82 == _h_T_1) begin // @[vga.scala 64:24]
        ram_130 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h82 == _T_37) begin // @[vga.scala 64:24]
        ram_130 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_130 <= _GEN_15358;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_131 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h83 == _h_T_1) begin // @[vga.scala 64:24]
        ram_131 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h83 == _T_37) begin // @[vga.scala 64:24]
        ram_131 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_131 <= _GEN_15359;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_132 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h84 == _h_T_1) begin // @[vga.scala 64:24]
        ram_132 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h84 == _T_37) begin // @[vga.scala 64:24]
        ram_132 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_132 <= _GEN_15360;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_133 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h85 == _h_T_1) begin // @[vga.scala 64:24]
        ram_133 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h85 == _T_37) begin // @[vga.scala 64:24]
        ram_133 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_133 <= _GEN_15361;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_134 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h86 == _h_T_1) begin // @[vga.scala 64:24]
        ram_134 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h86 == _T_37) begin // @[vga.scala 64:24]
        ram_134 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_134 <= _GEN_15362;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_135 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h87 == _h_T_1) begin // @[vga.scala 64:24]
        ram_135 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h87 == _T_37) begin // @[vga.scala 64:24]
        ram_135 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_135 <= _GEN_15363;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_136 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h88 == _h_T_1) begin // @[vga.scala 64:24]
        ram_136 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h88 == _T_37) begin // @[vga.scala 64:24]
        ram_136 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_136 <= _GEN_15364;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_137 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h89 == _h_T_1) begin // @[vga.scala 64:24]
        ram_137 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h89 == _T_37) begin // @[vga.scala 64:24]
        ram_137 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_137 <= _GEN_15365;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_138 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8a == _h_T_1) begin // @[vga.scala 64:24]
        ram_138 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8a == _T_37) begin // @[vga.scala 64:24]
        ram_138 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_138 <= _GEN_15366;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_139 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8b == _h_T_1) begin // @[vga.scala 64:24]
        ram_139 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8b == _T_37) begin // @[vga.scala 64:24]
        ram_139 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_139 <= _GEN_15367;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_140 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8c == _h_T_1) begin // @[vga.scala 64:24]
        ram_140 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8c == _T_37) begin // @[vga.scala 64:24]
        ram_140 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_140 <= _GEN_15368;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_141 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8d == _h_T_1) begin // @[vga.scala 64:24]
        ram_141 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8d == _T_37) begin // @[vga.scala 64:24]
        ram_141 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_141 <= _GEN_15369;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_142 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8e == _h_T_1) begin // @[vga.scala 64:24]
        ram_142 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8e == _T_37) begin // @[vga.scala 64:24]
        ram_142 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_142 <= _GEN_15370;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_143 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h8f == _h_T_1) begin // @[vga.scala 64:24]
        ram_143 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h8f == _T_37) begin // @[vga.scala 64:24]
        ram_143 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_143 <= _GEN_15371;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_144 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h90 == _h_T_1) begin // @[vga.scala 64:24]
        ram_144 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h90 == _T_37) begin // @[vga.scala 64:24]
        ram_144 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_144 <= _GEN_15372;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_145 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h91 == _h_T_1) begin // @[vga.scala 64:24]
        ram_145 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h91 == _T_37) begin // @[vga.scala 64:24]
        ram_145 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_145 <= _GEN_15373;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_146 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h92 == _h_T_1) begin // @[vga.scala 64:24]
        ram_146 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h92 == _T_37) begin // @[vga.scala 64:24]
        ram_146 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_146 <= _GEN_15374;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_147 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h93 == _h_T_1) begin // @[vga.scala 64:24]
        ram_147 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h93 == _T_37) begin // @[vga.scala 64:24]
        ram_147 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_147 <= _GEN_15375;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_148 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h94 == _h_T_1) begin // @[vga.scala 64:24]
        ram_148 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h94 == _T_37) begin // @[vga.scala 64:24]
        ram_148 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_148 <= _GEN_15376;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_149 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h95 == _h_T_1) begin // @[vga.scala 64:24]
        ram_149 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h95 == _T_37) begin // @[vga.scala 64:24]
        ram_149 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_149 <= _GEN_15377;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_150 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h96 == _h_T_1) begin // @[vga.scala 64:24]
        ram_150 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h96 == _T_37) begin // @[vga.scala 64:24]
        ram_150 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_150 <= _GEN_15378;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_151 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h97 == _h_T_1) begin // @[vga.scala 64:24]
        ram_151 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h97 == _T_37) begin // @[vga.scala 64:24]
        ram_151 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_151 <= _GEN_15379;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_152 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h98 == _h_T_1) begin // @[vga.scala 64:24]
        ram_152 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h98 == _T_37) begin // @[vga.scala 64:24]
        ram_152 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_152 <= _GEN_15380;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_153 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h99 == _h_T_1) begin // @[vga.scala 64:24]
        ram_153 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h99 == _T_37) begin // @[vga.scala 64:24]
        ram_153 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_153 <= _GEN_15381;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_154 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9a == _h_T_1) begin // @[vga.scala 64:24]
        ram_154 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9a == _T_37) begin // @[vga.scala 64:24]
        ram_154 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_154 <= _GEN_15382;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_155 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9b == _h_T_1) begin // @[vga.scala 64:24]
        ram_155 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9b == _T_37) begin // @[vga.scala 64:24]
        ram_155 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_155 <= _GEN_15383;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_156 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9c == _h_T_1) begin // @[vga.scala 64:24]
        ram_156 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9c == _T_37) begin // @[vga.scala 64:24]
        ram_156 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_156 <= _GEN_15384;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_157 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9d == _h_T_1) begin // @[vga.scala 64:24]
        ram_157 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9d == _T_37) begin // @[vga.scala 64:24]
        ram_157 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_157 <= _GEN_15385;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_158 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9e == _h_T_1) begin // @[vga.scala 64:24]
        ram_158 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9e == _T_37) begin // @[vga.scala 64:24]
        ram_158 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_158 <= _GEN_15386;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_159 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h9f == _h_T_1) begin // @[vga.scala 64:24]
        ram_159 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h9f == _T_37) begin // @[vga.scala 64:24]
        ram_159 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_159 <= _GEN_15387;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_160 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_160 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha0 == _T_37) begin // @[vga.scala 64:24]
        ram_160 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_160 <= _GEN_15388;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_161 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_161 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha1 == _T_37) begin // @[vga.scala 64:24]
        ram_161 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_161 <= _GEN_15389;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_162 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_162 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha2 == _T_37) begin // @[vga.scala 64:24]
        ram_162 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_162 <= _GEN_15390;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_163 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_163 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha3 == _T_37) begin // @[vga.scala 64:24]
        ram_163 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_163 <= _GEN_15391;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_164 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_164 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha4 == _T_37) begin // @[vga.scala 64:24]
        ram_164 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_164 <= _GEN_15392;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_165 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_165 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha5 == _T_37) begin // @[vga.scala 64:24]
        ram_165 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_165 <= _GEN_15393;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_166 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_166 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha6 == _T_37) begin // @[vga.scala 64:24]
        ram_166 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_166 <= _GEN_15394;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_167 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_167 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha7 == _T_37) begin // @[vga.scala 64:24]
        ram_167 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_167 <= _GEN_15395;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_168 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_168 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha8 == _T_37) begin // @[vga.scala 64:24]
        ram_168 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_168 <= _GEN_15396;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_169 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'ha9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_169 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'ha9 == _T_37) begin // @[vga.scala 64:24]
        ram_169 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_169 <= _GEN_15397;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_170 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'haa == _h_T_1) begin // @[vga.scala 64:24]
        ram_170 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'haa == _T_37) begin // @[vga.scala 64:24]
        ram_170 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_170 <= _GEN_15398;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_171 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hab == _h_T_1) begin // @[vga.scala 64:24]
        ram_171 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hab == _T_37) begin // @[vga.scala 64:24]
        ram_171 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_171 <= _GEN_15399;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_172 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hac == _h_T_1) begin // @[vga.scala 64:24]
        ram_172 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hac == _T_37) begin // @[vga.scala 64:24]
        ram_172 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_172 <= _GEN_15400;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_173 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'had == _h_T_1) begin // @[vga.scala 64:24]
        ram_173 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'had == _T_37) begin // @[vga.scala 64:24]
        ram_173 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_173 <= _GEN_15401;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_174 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hae == _h_T_1) begin // @[vga.scala 64:24]
        ram_174 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hae == _T_37) begin // @[vga.scala 64:24]
        ram_174 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_174 <= _GEN_15402;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_175 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'haf == _h_T_1) begin // @[vga.scala 64:24]
        ram_175 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'haf == _T_37) begin // @[vga.scala 64:24]
        ram_175 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_175 <= _GEN_15403;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_176 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_176 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb0 == _T_37) begin // @[vga.scala 64:24]
        ram_176 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_176 <= _GEN_15404;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_177 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_177 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb1 == _T_37) begin // @[vga.scala 64:24]
        ram_177 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_177 <= _GEN_15405;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_178 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_178 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb2 == _T_37) begin // @[vga.scala 64:24]
        ram_178 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_178 <= _GEN_15406;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_179 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_179 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb3 == _T_37) begin // @[vga.scala 64:24]
        ram_179 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_179 <= _GEN_15407;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_180 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_180 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb4 == _T_37) begin // @[vga.scala 64:24]
        ram_180 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_180 <= _GEN_15408;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_181 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_181 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb5 == _T_37) begin // @[vga.scala 64:24]
        ram_181 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_181 <= _GEN_15409;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_182 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_182 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb6 == _T_37) begin // @[vga.scala 64:24]
        ram_182 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_182 <= _GEN_15410;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_183 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_183 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb7 == _T_37) begin // @[vga.scala 64:24]
        ram_183 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_183 <= _GEN_15411;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_184 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_184 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb8 == _T_37) begin // @[vga.scala 64:24]
        ram_184 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_184 <= _GEN_15412;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_185 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hb9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_185 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hb9 == _T_37) begin // @[vga.scala 64:24]
        ram_185 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_185 <= _GEN_15413;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_186 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hba == _h_T_1) begin // @[vga.scala 64:24]
        ram_186 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hba == _T_37) begin // @[vga.scala 64:24]
        ram_186 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_186 <= _GEN_15414;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_187 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hbb == _h_T_1) begin // @[vga.scala 64:24]
        ram_187 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hbb == _T_37) begin // @[vga.scala 64:24]
        ram_187 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_187 <= _GEN_15415;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_188 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hbc == _h_T_1) begin // @[vga.scala 64:24]
        ram_188 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hbc == _T_37) begin // @[vga.scala 64:24]
        ram_188 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_188 <= _GEN_15416;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_189 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hbd == _h_T_1) begin // @[vga.scala 64:24]
        ram_189 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hbd == _T_37) begin // @[vga.scala 64:24]
        ram_189 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_189 <= _GEN_15417;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_190 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hbe == _h_T_1) begin // @[vga.scala 64:24]
        ram_190 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hbe == _T_37) begin // @[vga.scala 64:24]
        ram_190 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_190 <= _GEN_15418;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_191 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hbf == _h_T_1) begin // @[vga.scala 64:24]
        ram_191 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hbf == _T_37) begin // @[vga.scala 64:24]
        ram_191 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_191 <= _GEN_15419;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_192 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_192 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc0 == _T_37) begin // @[vga.scala 64:24]
        ram_192 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_192 <= _GEN_15420;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_193 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_193 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc1 == _T_37) begin // @[vga.scala 64:24]
        ram_193 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_193 <= _GEN_15421;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_194 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_194 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc2 == _T_37) begin // @[vga.scala 64:24]
        ram_194 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_194 <= _GEN_15422;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_195 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_195 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc3 == _T_37) begin // @[vga.scala 64:24]
        ram_195 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_195 <= _GEN_15423;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_196 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_196 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc4 == _T_37) begin // @[vga.scala 64:24]
        ram_196 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_196 <= _GEN_15424;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_197 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_197 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc5 == _T_37) begin // @[vga.scala 64:24]
        ram_197 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_197 <= _GEN_15425;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_198 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_198 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc6 == _T_37) begin // @[vga.scala 64:24]
        ram_198 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_198 <= _GEN_15426;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_199 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_199 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc7 == _T_37) begin // @[vga.scala 64:24]
        ram_199 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_199 <= _GEN_15427;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_200 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_200 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc8 == _T_37) begin // @[vga.scala 64:24]
        ram_200 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_200 <= _GEN_15428;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_201 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hc9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_201 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hc9 == _T_37) begin // @[vga.scala 64:24]
        ram_201 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_201 <= _GEN_15429;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_202 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hca == _h_T_1) begin // @[vga.scala 64:24]
        ram_202 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hca == _T_37) begin // @[vga.scala 64:24]
        ram_202 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_202 <= _GEN_15430;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_203 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hcb == _h_T_1) begin // @[vga.scala 64:24]
        ram_203 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hcb == _T_37) begin // @[vga.scala 64:24]
        ram_203 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_203 <= _GEN_15431;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_204 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hcc == _h_T_1) begin // @[vga.scala 64:24]
        ram_204 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hcc == _T_37) begin // @[vga.scala 64:24]
        ram_204 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_204 <= _GEN_15432;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_205 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hcd == _h_T_1) begin // @[vga.scala 64:24]
        ram_205 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hcd == _T_37) begin // @[vga.scala 64:24]
        ram_205 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_205 <= _GEN_15433;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_206 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hce == _h_T_1) begin // @[vga.scala 64:24]
        ram_206 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hce == _T_37) begin // @[vga.scala 64:24]
        ram_206 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_206 <= _GEN_15434;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_207 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hcf == _h_T_1) begin // @[vga.scala 64:24]
        ram_207 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hcf == _T_37) begin // @[vga.scala 64:24]
        ram_207 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_207 <= _GEN_15435;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_208 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_208 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd0 == _T_37) begin // @[vga.scala 64:24]
        ram_208 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_208 <= _GEN_15436;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_209 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_209 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd1 == _T_37) begin // @[vga.scala 64:24]
        ram_209 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_209 <= _GEN_15437;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_210 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_210 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd2 == _T_37) begin // @[vga.scala 64:24]
        ram_210 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_210 <= _GEN_15438;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_211 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_211 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd3 == _T_37) begin // @[vga.scala 64:24]
        ram_211 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_211 <= _GEN_15439;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_212 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_212 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd4 == _T_37) begin // @[vga.scala 64:24]
        ram_212 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_212 <= _GEN_15440;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_213 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_213 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd5 == _T_37) begin // @[vga.scala 64:24]
        ram_213 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_213 <= _GEN_15441;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_214 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_214 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd6 == _T_37) begin // @[vga.scala 64:24]
        ram_214 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_214 <= _GEN_15442;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_215 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_215 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd7 == _T_37) begin // @[vga.scala 64:24]
        ram_215 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_215 <= _GEN_15443;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_216 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_216 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd8 == _T_37) begin // @[vga.scala 64:24]
        ram_216 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_216 <= _GEN_15444;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_217 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hd9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_217 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hd9 == _T_37) begin // @[vga.scala 64:24]
        ram_217 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_217 <= _GEN_15445;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_218 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hda == _h_T_1) begin // @[vga.scala 64:24]
        ram_218 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hda == _T_37) begin // @[vga.scala 64:24]
        ram_218 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_218 <= _GEN_15446;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_219 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hdb == _h_T_1) begin // @[vga.scala 64:24]
        ram_219 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hdb == _T_37) begin // @[vga.scala 64:24]
        ram_219 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_219 <= _GEN_15447;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_220 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hdc == _h_T_1) begin // @[vga.scala 64:24]
        ram_220 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hdc == _T_37) begin // @[vga.scala 64:24]
        ram_220 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_220 <= _GEN_15448;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_221 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hdd == _h_T_1) begin // @[vga.scala 64:24]
        ram_221 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hdd == _T_37) begin // @[vga.scala 64:24]
        ram_221 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_221 <= _GEN_15449;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_222 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hde == _h_T_1) begin // @[vga.scala 64:24]
        ram_222 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hde == _T_37) begin // @[vga.scala 64:24]
        ram_222 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_222 <= _GEN_15450;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_223 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hdf == _h_T_1) begin // @[vga.scala 64:24]
        ram_223 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hdf == _T_37) begin // @[vga.scala 64:24]
        ram_223 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_223 <= _GEN_15451;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_224 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_224 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he0 == _T_37) begin // @[vga.scala 64:24]
        ram_224 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_224 <= _GEN_15452;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_225 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_225 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he1 == _T_37) begin // @[vga.scala 64:24]
        ram_225 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_225 <= _GEN_15453;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_226 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_226 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he2 == _T_37) begin // @[vga.scala 64:24]
        ram_226 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_226 <= _GEN_15454;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_227 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_227 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he3 == _T_37) begin // @[vga.scala 64:24]
        ram_227 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_227 <= _GEN_15455;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_228 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_228 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he4 == _T_37) begin // @[vga.scala 64:24]
        ram_228 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_228 <= _GEN_15456;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_229 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_229 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he5 == _T_37) begin // @[vga.scala 64:24]
        ram_229 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_229 <= _GEN_15457;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_230 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_230 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he6 == _T_37) begin // @[vga.scala 64:24]
        ram_230 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_230 <= _GEN_15458;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_231 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_231 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he7 == _T_37) begin // @[vga.scala 64:24]
        ram_231 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_231 <= _GEN_15459;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_232 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_232 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he8 == _T_37) begin // @[vga.scala 64:24]
        ram_232 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_232 <= _GEN_15460;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_233 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'he9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_233 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'he9 == _T_37) begin // @[vga.scala 64:24]
        ram_233 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_233 <= _GEN_15461;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_234 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hea == _h_T_1) begin // @[vga.scala 64:24]
        ram_234 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hea == _T_37) begin // @[vga.scala 64:24]
        ram_234 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_234 <= _GEN_15462;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_235 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'heb == _h_T_1) begin // @[vga.scala 64:24]
        ram_235 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'heb == _T_37) begin // @[vga.scala 64:24]
        ram_235 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_235 <= _GEN_15463;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_236 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hec == _h_T_1) begin // @[vga.scala 64:24]
        ram_236 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hec == _T_37) begin // @[vga.scala 64:24]
        ram_236 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_236 <= _GEN_15464;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_237 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hed == _h_T_1) begin // @[vga.scala 64:24]
        ram_237 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hed == _T_37) begin // @[vga.scala 64:24]
        ram_237 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_237 <= _GEN_15465;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_238 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hee == _h_T_1) begin // @[vga.scala 64:24]
        ram_238 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hee == _T_37) begin // @[vga.scala 64:24]
        ram_238 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_238 <= _GEN_15466;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_239 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hef == _h_T_1) begin // @[vga.scala 64:24]
        ram_239 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hef == _T_37) begin // @[vga.scala 64:24]
        ram_239 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_239 <= _GEN_15467;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_240 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_240 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf0 == _T_37) begin // @[vga.scala 64:24]
        ram_240 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_240 <= _GEN_15468;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_241 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_241 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf1 == _T_37) begin // @[vga.scala 64:24]
        ram_241 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_241 <= _GEN_15469;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_242 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_242 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf2 == _T_37) begin // @[vga.scala 64:24]
        ram_242 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_242 <= _GEN_15470;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_243 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_243 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf3 == _T_37) begin // @[vga.scala 64:24]
        ram_243 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_243 <= _GEN_15471;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_244 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_244 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf4 == _T_37) begin // @[vga.scala 64:24]
        ram_244 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_244 <= _GEN_15472;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_245 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_245 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf5 == _T_37) begin // @[vga.scala 64:24]
        ram_245 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_245 <= _GEN_15473;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_246 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_246 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf6 == _T_37) begin // @[vga.scala 64:24]
        ram_246 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_246 <= _GEN_15474;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_247 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_247 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf7 == _T_37) begin // @[vga.scala 64:24]
        ram_247 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_247 <= _GEN_15475;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_248 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_248 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf8 == _T_37) begin // @[vga.scala 64:24]
        ram_248 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_248 <= _GEN_15476;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_249 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hf9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_249 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hf9 == _T_37) begin // @[vga.scala 64:24]
        ram_249 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_249 <= _GEN_15477;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_250 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hfa == _h_T_1) begin // @[vga.scala 64:24]
        ram_250 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hfa == _T_37) begin // @[vga.scala 64:24]
        ram_250 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_250 <= _GEN_15478;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_251 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hfb == _h_T_1) begin // @[vga.scala 64:24]
        ram_251 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hfb == _T_37) begin // @[vga.scala 64:24]
        ram_251 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_251 <= _GEN_15479;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_252 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hfc == _h_T_1) begin // @[vga.scala 64:24]
        ram_252 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hfc == _T_37) begin // @[vga.scala 64:24]
        ram_252 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_252 <= _GEN_15480;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_253 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hfd == _h_T_1) begin // @[vga.scala 64:24]
        ram_253 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hfd == _T_37) begin // @[vga.scala 64:24]
        ram_253 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_253 <= _GEN_15481;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_254 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hfe == _h_T_1) begin // @[vga.scala 64:24]
        ram_254 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hfe == _T_37) begin // @[vga.scala 64:24]
        ram_254 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_254 <= _GEN_15482;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_255 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'hff == _h_T_1) begin // @[vga.scala 64:24]
        ram_255 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'hff == _T_37) begin // @[vga.scala 64:24]
        ram_255 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_255 <= _GEN_15483;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_256 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h100 == _h_T_1) begin // @[vga.scala 64:24]
        ram_256 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h100 == _T_37) begin // @[vga.scala 64:24]
        ram_256 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_256 <= _GEN_15484;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_257 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h101 == _h_T_1) begin // @[vga.scala 64:24]
        ram_257 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h101 == _T_37) begin // @[vga.scala 64:24]
        ram_257 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_257 <= _GEN_15485;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_258 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h102 == _h_T_1) begin // @[vga.scala 64:24]
        ram_258 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h102 == _T_37) begin // @[vga.scala 64:24]
        ram_258 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_258 <= _GEN_15486;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_259 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h103 == _h_T_1) begin // @[vga.scala 64:24]
        ram_259 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h103 == _T_37) begin // @[vga.scala 64:24]
        ram_259 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_259 <= _GEN_15487;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_260 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h104 == _h_T_1) begin // @[vga.scala 64:24]
        ram_260 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h104 == _T_37) begin // @[vga.scala 64:24]
        ram_260 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_260 <= _GEN_15488;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_261 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h105 == _h_T_1) begin // @[vga.scala 64:24]
        ram_261 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h105 == _T_37) begin // @[vga.scala 64:24]
        ram_261 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_261 <= _GEN_15489;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_262 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h106 == _h_T_1) begin // @[vga.scala 64:24]
        ram_262 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h106 == _T_37) begin // @[vga.scala 64:24]
        ram_262 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_262 <= _GEN_15490;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_263 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h107 == _h_T_1) begin // @[vga.scala 64:24]
        ram_263 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h107 == _T_37) begin // @[vga.scala 64:24]
        ram_263 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_263 <= _GEN_15491;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_264 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h108 == _h_T_1) begin // @[vga.scala 64:24]
        ram_264 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h108 == _T_37) begin // @[vga.scala 64:24]
        ram_264 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_264 <= _GEN_15492;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_265 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h109 == _h_T_1) begin // @[vga.scala 64:24]
        ram_265 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h109 == _T_37) begin // @[vga.scala 64:24]
        ram_265 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_265 <= _GEN_15493;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_266 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10a == _h_T_1) begin // @[vga.scala 64:24]
        ram_266 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10a == _T_37) begin // @[vga.scala 64:24]
        ram_266 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_266 <= _GEN_15494;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_267 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10b == _h_T_1) begin // @[vga.scala 64:24]
        ram_267 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10b == _T_37) begin // @[vga.scala 64:24]
        ram_267 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_267 <= _GEN_15495;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_268 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10c == _h_T_1) begin // @[vga.scala 64:24]
        ram_268 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10c == _T_37) begin // @[vga.scala 64:24]
        ram_268 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_268 <= _GEN_15496;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_269 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10d == _h_T_1) begin // @[vga.scala 64:24]
        ram_269 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10d == _T_37) begin // @[vga.scala 64:24]
        ram_269 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_269 <= _GEN_15497;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_270 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10e == _h_T_1) begin // @[vga.scala 64:24]
        ram_270 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10e == _T_37) begin // @[vga.scala 64:24]
        ram_270 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_270 <= _GEN_15498;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_271 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h10f == _h_T_1) begin // @[vga.scala 64:24]
        ram_271 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h10f == _T_37) begin // @[vga.scala 64:24]
        ram_271 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_271 <= _GEN_15499;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_272 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h110 == _h_T_1) begin // @[vga.scala 64:24]
        ram_272 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h110 == _T_37) begin // @[vga.scala 64:24]
        ram_272 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_272 <= _GEN_15500;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_273 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h111 == _h_T_1) begin // @[vga.scala 64:24]
        ram_273 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h111 == _T_37) begin // @[vga.scala 64:24]
        ram_273 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_273 <= _GEN_15501;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_274 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h112 == _h_T_1) begin // @[vga.scala 64:24]
        ram_274 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h112 == _T_37) begin // @[vga.scala 64:24]
        ram_274 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_274 <= _GEN_15502;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_275 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h113 == _h_T_1) begin // @[vga.scala 64:24]
        ram_275 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h113 == _T_37) begin // @[vga.scala 64:24]
        ram_275 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_275 <= _GEN_15503;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_276 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h114 == _h_T_1) begin // @[vga.scala 64:24]
        ram_276 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h114 == _T_37) begin // @[vga.scala 64:24]
        ram_276 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_276 <= _GEN_15504;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_277 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h115 == _h_T_1) begin // @[vga.scala 64:24]
        ram_277 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h115 == _T_37) begin // @[vga.scala 64:24]
        ram_277 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_277 <= _GEN_15505;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_278 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h116 == _h_T_1) begin // @[vga.scala 64:24]
        ram_278 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h116 == _T_37) begin // @[vga.scala 64:24]
        ram_278 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_278 <= _GEN_15506;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_279 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h117 == _h_T_1) begin // @[vga.scala 64:24]
        ram_279 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h117 == _T_37) begin // @[vga.scala 64:24]
        ram_279 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_279 <= _GEN_15507;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_280 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h118 == _h_T_1) begin // @[vga.scala 64:24]
        ram_280 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h118 == _T_37) begin // @[vga.scala 64:24]
        ram_280 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_280 <= _GEN_15508;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_281 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h119 == _h_T_1) begin // @[vga.scala 64:24]
        ram_281 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h119 == _T_37) begin // @[vga.scala 64:24]
        ram_281 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_281 <= _GEN_15509;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_282 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11a == _h_T_1) begin // @[vga.scala 64:24]
        ram_282 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11a == _T_37) begin // @[vga.scala 64:24]
        ram_282 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_282 <= _GEN_15510;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_283 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11b == _h_T_1) begin // @[vga.scala 64:24]
        ram_283 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11b == _T_37) begin // @[vga.scala 64:24]
        ram_283 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_283 <= _GEN_15511;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_284 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11c == _h_T_1) begin // @[vga.scala 64:24]
        ram_284 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11c == _T_37) begin // @[vga.scala 64:24]
        ram_284 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_284 <= _GEN_15512;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_285 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11d == _h_T_1) begin // @[vga.scala 64:24]
        ram_285 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11d == _T_37) begin // @[vga.scala 64:24]
        ram_285 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_285 <= _GEN_15513;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_286 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11e == _h_T_1) begin // @[vga.scala 64:24]
        ram_286 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11e == _T_37) begin // @[vga.scala 64:24]
        ram_286 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_286 <= _GEN_15514;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_287 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h11f == _h_T_1) begin // @[vga.scala 64:24]
        ram_287 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h11f == _T_37) begin // @[vga.scala 64:24]
        ram_287 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_287 <= _GEN_15515;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_288 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h120 == _h_T_1) begin // @[vga.scala 64:24]
        ram_288 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h120 == _T_37) begin // @[vga.scala 64:24]
        ram_288 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_288 <= _GEN_15516;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_289 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h121 == _h_T_1) begin // @[vga.scala 64:24]
        ram_289 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h121 == _T_37) begin // @[vga.scala 64:24]
        ram_289 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_289 <= _GEN_15517;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_290 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h122 == _h_T_1) begin // @[vga.scala 64:24]
        ram_290 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h122 == _T_37) begin // @[vga.scala 64:24]
        ram_290 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_290 <= _GEN_15518;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_291 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h123 == _h_T_1) begin // @[vga.scala 64:24]
        ram_291 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h123 == _T_37) begin // @[vga.scala 64:24]
        ram_291 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_291 <= _GEN_15519;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_292 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h124 == _h_T_1) begin // @[vga.scala 64:24]
        ram_292 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h124 == _T_37) begin // @[vga.scala 64:24]
        ram_292 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_292 <= _GEN_15520;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_293 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h125 == _h_T_1) begin // @[vga.scala 64:24]
        ram_293 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h125 == _T_37) begin // @[vga.scala 64:24]
        ram_293 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_293 <= _GEN_15521;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_294 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h126 == _h_T_1) begin // @[vga.scala 64:24]
        ram_294 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h126 == _T_37) begin // @[vga.scala 64:24]
        ram_294 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_294 <= _GEN_15522;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_295 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h127 == _h_T_1) begin // @[vga.scala 64:24]
        ram_295 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h127 == _T_37) begin // @[vga.scala 64:24]
        ram_295 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_295 <= _GEN_15523;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_296 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h128 == _h_T_1) begin // @[vga.scala 64:24]
        ram_296 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h128 == _T_37) begin // @[vga.scala 64:24]
        ram_296 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_296 <= _GEN_15524;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_297 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h129 == _h_T_1) begin // @[vga.scala 64:24]
        ram_297 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h129 == _T_37) begin // @[vga.scala 64:24]
        ram_297 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_297 <= _GEN_15525;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_298 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12a == _h_T_1) begin // @[vga.scala 64:24]
        ram_298 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12a == _T_37) begin // @[vga.scala 64:24]
        ram_298 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_298 <= _GEN_15526;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_299 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12b == _h_T_1) begin // @[vga.scala 64:24]
        ram_299 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12b == _T_37) begin // @[vga.scala 64:24]
        ram_299 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_299 <= _GEN_15527;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_300 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12c == _h_T_1) begin // @[vga.scala 64:24]
        ram_300 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12c == _T_37) begin // @[vga.scala 64:24]
        ram_300 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_300 <= _GEN_15528;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_301 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12d == _h_T_1) begin // @[vga.scala 64:24]
        ram_301 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12d == _T_37) begin // @[vga.scala 64:24]
        ram_301 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_301 <= _GEN_15529;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_302 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12e == _h_T_1) begin // @[vga.scala 64:24]
        ram_302 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12e == _T_37) begin // @[vga.scala 64:24]
        ram_302 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_302 <= _GEN_15530;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_303 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h12f == _h_T_1) begin // @[vga.scala 64:24]
        ram_303 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h12f == _T_37) begin // @[vga.scala 64:24]
        ram_303 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_303 <= _GEN_15531;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_304 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h130 == _h_T_1) begin // @[vga.scala 64:24]
        ram_304 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h130 == _T_37) begin // @[vga.scala 64:24]
        ram_304 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_304 <= _GEN_15532;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_305 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h131 == _h_T_1) begin // @[vga.scala 64:24]
        ram_305 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h131 == _T_37) begin // @[vga.scala 64:24]
        ram_305 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_305 <= _GEN_15533;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_306 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h132 == _h_T_1) begin // @[vga.scala 64:24]
        ram_306 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h132 == _T_37) begin // @[vga.scala 64:24]
        ram_306 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_306 <= _GEN_15534;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_307 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h133 == _h_T_1) begin // @[vga.scala 64:24]
        ram_307 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h133 == _T_37) begin // @[vga.scala 64:24]
        ram_307 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_307 <= _GEN_15535;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_308 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h134 == _h_T_1) begin // @[vga.scala 64:24]
        ram_308 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h134 == _T_37) begin // @[vga.scala 64:24]
        ram_308 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_308 <= _GEN_15536;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_309 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h135 == _h_T_1) begin // @[vga.scala 64:24]
        ram_309 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h135 == _T_37) begin // @[vga.scala 64:24]
        ram_309 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_309 <= _GEN_15537;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_310 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h136 == _h_T_1) begin // @[vga.scala 64:24]
        ram_310 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h136 == _T_37) begin // @[vga.scala 64:24]
        ram_310 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_310 <= _GEN_15538;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_311 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h137 == _h_T_1) begin // @[vga.scala 64:24]
        ram_311 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h137 == _T_37) begin // @[vga.scala 64:24]
        ram_311 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_311 <= _GEN_15539;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_312 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h138 == _h_T_1) begin // @[vga.scala 64:24]
        ram_312 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h138 == _T_37) begin // @[vga.scala 64:24]
        ram_312 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_312 <= _GEN_15540;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_313 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h139 == _h_T_1) begin // @[vga.scala 64:24]
        ram_313 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h139 == _T_37) begin // @[vga.scala 64:24]
        ram_313 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_313 <= _GEN_15541;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_314 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13a == _h_T_1) begin // @[vga.scala 64:24]
        ram_314 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13a == _T_37) begin // @[vga.scala 64:24]
        ram_314 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_314 <= _GEN_15542;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_315 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13b == _h_T_1) begin // @[vga.scala 64:24]
        ram_315 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13b == _T_37) begin // @[vga.scala 64:24]
        ram_315 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_315 <= _GEN_15543;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_316 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13c == _h_T_1) begin // @[vga.scala 64:24]
        ram_316 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13c == _T_37) begin // @[vga.scala 64:24]
        ram_316 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_316 <= _GEN_15544;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_317 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13d == _h_T_1) begin // @[vga.scala 64:24]
        ram_317 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13d == _T_37) begin // @[vga.scala 64:24]
        ram_317 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_317 <= _GEN_15545;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_318 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13e == _h_T_1) begin // @[vga.scala 64:24]
        ram_318 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13e == _T_37) begin // @[vga.scala 64:24]
        ram_318 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_318 <= _GEN_15546;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_319 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h13f == _h_T_1) begin // @[vga.scala 64:24]
        ram_319 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h13f == _T_37) begin // @[vga.scala 64:24]
        ram_319 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_319 <= _GEN_15547;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_320 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h140 == _h_T_1) begin // @[vga.scala 64:24]
        ram_320 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h140 == _T_37) begin // @[vga.scala 64:24]
        ram_320 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_320 <= _GEN_15548;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_321 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h141 == _h_T_1) begin // @[vga.scala 64:24]
        ram_321 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h141 == _T_37) begin // @[vga.scala 64:24]
        ram_321 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_321 <= _GEN_15549;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_322 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h142 == _h_T_1) begin // @[vga.scala 64:24]
        ram_322 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h142 == _T_37) begin // @[vga.scala 64:24]
        ram_322 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_322 <= _GEN_15550;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_323 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h143 == _h_T_1) begin // @[vga.scala 64:24]
        ram_323 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h143 == _T_37) begin // @[vga.scala 64:24]
        ram_323 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_323 <= _GEN_15551;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_324 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h144 == _h_T_1) begin // @[vga.scala 64:24]
        ram_324 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h144 == _T_37) begin // @[vga.scala 64:24]
        ram_324 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_324 <= _GEN_15552;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_325 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h145 == _h_T_1) begin // @[vga.scala 64:24]
        ram_325 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h145 == _T_37) begin // @[vga.scala 64:24]
        ram_325 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_325 <= _GEN_15553;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_326 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h146 == _h_T_1) begin // @[vga.scala 64:24]
        ram_326 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h146 == _T_37) begin // @[vga.scala 64:24]
        ram_326 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_326 <= _GEN_15554;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_327 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h147 == _h_T_1) begin // @[vga.scala 64:24]
        ram_327 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h147 == _T_37) begin // @[vga.scala 64:24]
        ram_327 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_327 <= _GEN_15555;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_328 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h148 == _h_T_1) begin // @[vga.scala 64:24]
        ram_328 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h148 == _T_37) begin // @[vga.scala 64:24]
        ram_328 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_328 <= _GEN_15556;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_329 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h149 == _h_T_1) begin // @[vga.scala 64:24]
        ram_329 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h149 == _T_37) begin // @[vga.scala 64:24]
        ram_329 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_329 <= _GEN_15557;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_330 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14a == _h_T_1) begin // @[vga.scala 64:24]
        ram_330 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14a == _T_37) begin // @[vga.scala 64:24]
        ram_330 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_330 <= _GEN_15558;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_331 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14b == _h_T_1) begin // @[vga.scala 64:24]
        ram_331 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14b == _T_37) begin // @[vga.scala 64:24]
        ram_331 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_331 <= _GEN_15559;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_332 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14c == _h_T_1) begin // @[vga.scala 64:24]
        ram_332 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14c == _T_37) begin // @[vga.scala 64:24]
        ram_332 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_332 <= _GEN_15560;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_333 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14d == _h_T_1) begin // @[vga.scala 64:24]
        ram_333 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14d == _T_37) begin // @[vga.scala 64:24]
        ram_333 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_333 <= _GEN_15561;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_334 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14e == _h_T_1) begin // @[vga.scala 64:24]
        ram_334 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14e == _T_37) begin // @[vga.scala 64:24]
        ram_334 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_334 <= _GEN_15562;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_335 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h14f == _h_T_1) begin // @[vga.scala 64:24]
        ram_335 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h14f == _T_37) begin // @[vga.scala 64:24]
        ram_335 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_335 <= _GEN_15563;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_336 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h150 == _h_T_1) begin // @[vga.scala 64:24]
        ram_336 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h150 == _T_37) begin // @[vga.scala 64:24]
        ram_336 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_336 <= _GEN_15564;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_337 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h151 == _h_T_1) begin // @[vga.scala 64:24]
        ram_337 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h151 == _T_37) begin // @[vga.scala 64:24]
        ram_337 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_337 <= _GEN_15565;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_338 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h152 == _h_T_1) begin // @[vga.scala 64:24]
        ram_338 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h152 == _T_37) begin // @[vga.scala 64:24]
        ram_338 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_338 <= _GEN_15566;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_339 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h153 == _h_T_1) begin // @[vga.scala 64:24]
        ram_339 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h153 == _T_37) begin // @[vga.scala 64:24]
        ram_339 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_339 <= _GEN_15567;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_340 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h154 == _h_T_1) begin // @[vga.scala 64:24]
        ram_340 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h154 == _T_37) begin // @[vga.scala 64:24]
        ram_340 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_340 <= _GEN_15568;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_341 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h155 == _h_T_1) begin // @[vga.scala 64:24]
        ram_341 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h155 == _T_37) begin // @[vga.scala 64:24]
        ram_341 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_341 <= _GEN_15569;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_342 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h156 == _h_T_1) begin // @[vga.scala 64:24]
        ram_342 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h156 == _T_37) begin // @[vga.scala 64:24]
        ram_342 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_342 <= _GEN_15570;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_343 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h157 == _h_T_1) begin // @[vga.scala 64:24]
        ram_343 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h157 == _T_37) begin // @[vga.scala 64:24]
        ram_343 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_343 <= _GEN_15571;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_344 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h158 == _h_T_1) begin // @[vga.scala 64:24]
        ram_344 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h158 == _T_37) begin // @[vga.scala 64:24]
        ram_344 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_344 <= _GEN_15572;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_345 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h159 == _h_T_1) begin // @[vga.scala 64:24]
        ram_345 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h159 == _T_37) begin // @[vga.scala 64:24]
        ram_345 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_345 <= _GEN_15573;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_346 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15a == _h_T_1) begin // @[vga.scala 64:24]
        ram_346 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15a == _T_37) begin // @[vga.scala 64:24]
        ram_346 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_346 <= _GEN_15574;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_347 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15b == _h_T_1) begin // @[vga.scala 64:24]
        ram_347 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15b == _T_37) begin // @[vga.scala 64:24]
        ram_347 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_347 <= _GEN_15575;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_348 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15c == _h_T_1) begin // @[vga.scala 64:24]
        ram_348 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15c == _T_37) begin // @[vga.scala 64:24]
        ram_348 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_348 <= _GEN_15576;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_349 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15d == _h_T_1) begin // @[vga.scala 64:24]
        ram_349 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15d == _T_37) begin // @[vga.scala 64:24]
        ram_349 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_349 <= _GEN_15577;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_350 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15e == _h_T_1) begin // @[vga.scala 64:24]
        ram_350 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15e == _T_37) begin // @[vga.scala 64:24]
        ram_350 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_350 <= _GEN_15578;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_351 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h15f == _h_T_1) begin // @[vga.scala 64:24]
        ram_351 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h15f == _T_37) begin // @[vga.scala 64:24]
        ram_351 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_351 <= _GEN_15579;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_352 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h160 == _h_T_1) begin // @[vga.scala 64:24]
        ram_352 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h160 == _T_37) begin // @[vga.scala 64:24]
        ram_352 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_352 <= _GEN_15580;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_353 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h161 == _h_T_1) begin // @[vga.scala 64:24]
        ram_353 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h161 == _T_37) begin // @[vga.scala 64:24]
        ram_353 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_353 <= _GEN_15581;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_354 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h162 == _h_T_1) begin // @[vga.scala 64:24]
        ram_354 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h162 == _T_37) begin // @[vga.scala 64:24]
        ram_354 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_354 <= _GEN_15582;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_355 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h163 == _h_T_1) begin // @[vga.scala 64:24]
        ram_355 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h163 == _T_37) begin // @[vga.scala 64:24]
        ram_355 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_355 <= _GEN_15583;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_356 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h164 == _h_T_1) begin // @[vga.scala 64:24]
        ram_356 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h164 == _T_37) begin // @[vga.scala 64:24]
        ram_356 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_356 <= _GEN_15584;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_357 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h165 == _h_T_1) begin // @[vga.scala 64:24]
        ram_357 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h165 == _T_37) begin // @[vga.scala 64:24]
        ram_357 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_357 <= _GEN_15585;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_358 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h166 == _h_T_1) begin // @[vga.scala 64:24]
        ram_358 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h166 == _T_37) begin // @[vga.scala 64:24]
        ram_358 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_358 <= _GEN_15586;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_359 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h167 == _h_T_1) begin // @[vga.scala 64:24]
        ram_359 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h167 == _T_37) begin // @[vga.scala 64:24]
        ram_359 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_359 <= _GEN_15587;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_360 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h168 == _h_T_1) begin // @[vga.scala 64:24]
        ram_360 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h168 == _T_37) begin // @[vga.scala 64:24]
        ram_360 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_360 <= _GEN_15588;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_361 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h169 == _h_T_1) begin // @[vga.scala 64:24]
        ram_361 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h169 == _T_37) begin // @[vga.scala 64:24]
        ram_361 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_361 <= _GEN_15589;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_362 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16a == _h_T_1) begin // @[vga.scala 64:24]
        ram_362 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16a == _T_37) begin // @[vga.scala 64:24]
        ram_362 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_362 <= _GEN_15590;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_363 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16b == _h_T_1) begin // @[vga.scala 64:24]
        ram_363 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16b == _T_37) begin // @[vga.scala 64:24]
        ram_363 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_363 <= _GEN_15591;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_364 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16c == _h_T_1) begin // @[vga.scala 64:24]
        ram_364 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16c == _T_37) begin // @[vga.scala 64:24]
        ram_364 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_364 <= _GEN_15592;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_365 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16d == _h_T_1) begin // @[vga.scala 64:24]
        ram_365 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16d == _T_37) begin // @[vga.scala 64:24]
        ram_365 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_365 <= _GEN_15593;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_366 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16e == _h_T_1) begin // @[vga.scala 64:24]
        ram_366 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16e == _T_37) begin // @[vga.scala 64:24]
        ram_366 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_366 <= _GEN_15594;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_367 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h16f == _h_T_1) begin // @[vga.scala 64:24]
        ram_367 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h16f == _T_37) begin // @[vga.scala 64:24]
        ram_367 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_367 <= _GEN_15595;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_368 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h170 == _h_T_1) begin // @[vga.scala 64:24]
        ram_368 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h170 == _T_37) begin // @[vga.scala 64:24]
        ram_368 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_368 <= _GEN_15596;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_369 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h171 == _h_T_1) begin // @[vga.scala 64:24]
        ram_369 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h171 == _T_37) begin // @[vga.scala 64:24]
        ram_369 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_369 <= _GEN_15597;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_370 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h172 == _h_T_1) begin // @[vga.scala 64:24]
        ram_370 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h172 == _T_37) begin // @[vga.scala 64:24]
        ram_370 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_370 <= _GEN_15598;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_371 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h173 == _h_T_1) begin // @[vga.scala 64:24]
        ram_371 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h173 == _T_37) begin // @[vga.scala 64:24]
        ram_371 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_371 <= _GEN_15599;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_372 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h174 == _h_T_1) begin // @[vga.scala 64:24]
        ram_372 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h174 == _T_37) begin // @[vga.scala 64:24]
        ram_372 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_372 <= _GEN_15600;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_373 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h175 == _h_T_1) begin // @[vga.scala 64:24]
        ram_373 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h175 == _T_37) begin // @[vga.scala 64:24]
        ram_373 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_373 <= _GEN_15601;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_374 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h176 == _h_T_1) begin // @[vga.scala 64:24]
        ram_374 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h176 == _T_37) begin // @[vga.scala 64:24]
        ram_374 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_374 <= _GEN_15602;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_375 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h177 == _h_T_1) begin // @[vga.scala 64:24]
        ram_375 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h177 == _T_37) begin // @[vga.scala 64:24]
        ram_375 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_375 <= _GEN_15603;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_376 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h178 == _h_T_1) begin // @[vga.scala 64:24]
        ram_376 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h178 == _T_37) begin // @[vga.scala 64:24]
        ram_376 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_376 <= _GEN_15604;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_377 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h179 == _h_T_1) begin // @[vga.scala 64:24]
        ram_377 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h179 == _T_37) begin // @[vga.scala 64:24]
        ram_377 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_377 <= _GEN_15605;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_378 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17a == _h_T_1) begin // @[vga.scala 64:24]
        ram_378 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17a == _T_37) begin // @[vga.scala 64:24]
        ram_378 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_378 <= _GEN_15606;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_379 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17b == _h_T_1) begin // @[vga.scala 64:24]
        ram_379 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17b == _T_37) begin // @[vga.scala 64:24]
        ram_379 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_379 <= _GEN_15607;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_380 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17c == _h_T_1) begin // @[vga.scala 64:24]
        ram_380 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17c == _T_37) begin // @[vga.scala 64:24]
        ram_380 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_380 <= _GEN_15608;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_381 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17d == _h_T_1) begin // @[vga.scala 64:24]
        ram_381 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17d == _T_37) begin // @[vga.scala 64:24]
        ram_381 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_381 <= _GEN_15609;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_382 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17e == _h_T_1) begin // @[vga.scala 64:24]
        ram_382 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17e == _T_37) begin // @[vga.scala 64:24]
        ram_382 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_382 <= _GEN_15610;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_383 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h17f == _h_T_1) begin // @[vga.scala 64:24]
        ram_383 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h17f == _T_37) begin // @[vga.scala 64:24]
        ram_383 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_383 <= _GEN_15611;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_384 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h180 == _h_T_1) begin // @[vga.scala 64:24]
        ram_384 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h180 == _T_37) begin // @[vga.scala 64:24]
        ram_384 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_384 <= _GEN_15612;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_385 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h181 == _h_T_1) begin // @[vga.scala 64:24]
        ram_385 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h181 == _T_37) begin // @[vga.scala 64:24]
        ram_385 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_385 <= _GEN_15613;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_386 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h182 == _h_T_1) begin // @[vga.scala 64:24]
        ram_386 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h182 == _T_37) begin // @[vga.scala 64:24]
        ram_386 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_386 <= _GEN_15614;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_387 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h183 == _h_T_1) begin // @[vga.scala 64:24]
        ram_387 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h183 == _T_37) begin // @[vga.scala 64:24]
        ram_387 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_387 <= _GEN_15615;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_388 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h184 == _h_T_1) begin // @[vga.scala 64:24]
        ram_388 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h184 == _T_37) begin // @[vga.scala 64:24]
        ram_388 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_388 <= _GEN_15616;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_389 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h185 == _h_T_1) begin // @[vga.scala 64:24]
        ram_389 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h185 == _T_37) begin // @[vga.scala 64:24]
        ram_389 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_389 <= _GEN_15617;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_390 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h186 == _h_T_1) begin // @[vga.scala 64:24]
        ram_390 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h186 == _T_37) begin // @[vga.scala 64:24]
        ram_390 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_390 <= _GEN_15618;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_391 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h187 == _h_T_1) begin // @[vga.scala 64:24]
        ram_391 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h187 == _T_37) begin // @[vga.scala 64:24]
        ram_391 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_391 <= _GEN_15619;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_392 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h188 == _h_T_1) begin // @[vga.scala 64:24]
        ram_392 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h188 == _T_37) begin // @[vga.scala 64:24]
        ram_392 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_392 <= _GEN_15620;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_393 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h189 == _h_T_1) begin // @[vga.scala 64:24]
        ram_393 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h189 == _T_37) begin // @[vga.scala 64:24]
        ram_393 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_393 <= _GEN_15621;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_394 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18a == _h_T_1) begin // @[vga.scala 64:24]
        ram_394 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18a == _T_37) begin // @[vga.scala 64:24]
        ram_394 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_394 <= _GEN_15622;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_395 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18b == _h_T_1) begin // @[vga.scala 64:24]
        ram_395 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18b == _T_37) begin // @[vga.scala 64:24]
        ram_395 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_395 <= _GEN_15623;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_396 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18c == _h_T_1) begin // @[vga.scala 64:24]
        ram_396 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18c == _T_37) begin // @[vga.scala 64:24]
        ram_396 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_396 <= _GEN_15624;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_397 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18d == _h_T_1) begin // @[vga.scala 64:24]
        ram_397 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18d == _T_37) begin // @[vga.scala 64:24]
        ram_397 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_397 <= _GEN_15625;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_398 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18e == _h_T_1) begin // @[vga.scala 64:24]
        ram_398 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18e == _T_37) begin // @[vga.scala 64:24]
        ram_398 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_398 <= _GEN_15626;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_399 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h18f == _h_T_1) begin // @[vga.scala 64:24]
        ram_399 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h18f == _T_37) begin // @[vga.scala 64:24]
        ram_399 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_399 <= _GEN_15627;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_400 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h190 == _h_T_1) begin // @[vga.scala 64:24]
        ram_400 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h190 == _T_37) begin // @[vga.scala 64:24]
        ram_400 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_400 <= _GEN_15628;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_401 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h191 == _h_T_1) begin // @[vga.scala 64:24]
        ram_401 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h191 == _T_37) begin // @[vga.scala 64:24]
        ram_401 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_401 <= _GEN_15629;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_402 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h192 == _h_T_1) begin // @[vga.scala 64:24]
        ram_402 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h192 == _T_37) begin // @[vga.scala 64:24]
        ram_402 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_402 <= _GEN_15630;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_403 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h193 == _h_T_1) begin // @[vga.scala 64:24]
        ram_403 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h193 == _T_37) begin // @[vga.scala 64:24]
        ram_403 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_403 <= _GEN_15631;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_404 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h194 == _h_T_1) begin // @[vga.scala 64:24]
        ram_404 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h194 == _T_37) begin // @[vga.scala 64:24]
        ram_404 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_404 <= _GEN_15632;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_405 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h195 == _h_T_1) begin // @[vga.scala 64:24]
        ram_405 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h195 == _T_37) begin // @[vga.scala 64:24]
        ram_405 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_405 <= _GEN_15633;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_406 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h196 == _h_T_1) begin // @[vga.scala 64:24]
        ram_406 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h196 == _T_37) begin // @[vga.scala 64:24]
        ram_406 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_406 <= _GEN_15634;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_407 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h197 == _h_T_1) begin // @[vga.scala 64:24]
        ram_407 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h197 == _T_37) begin // @[vga.scala 64:24]
        ram_407 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_407 <= _GEN_15635;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_408 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h198 == _h_T_1) begin // @[vga.scala 64:24]
        ram_408 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h198 == _T_37) begin // @[vga.scala 64:24]
        ram_408 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_408 <= _GEN_15636;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_409 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h199 == _h_T_1) begin // @[vga.scala 64:24]
        ram_409 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h199 == _T_37) begin // @[vga.scala 64:24]
        ram_409 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_409 <= _GEN_15637;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_410 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19a == _h_T_1) begin // @[vga.scala 64:24]
        ram_410 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19a == _T_37) begin // @[vga.scala 64:24]
        ram_410 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_410 <= _GEN_15638;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_411 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19b == _h_T_1) begin // @[vga.scala 64:24]
        ram_411 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19b == _T_37) begin // @[vga.scala 64:24]
        ram_411 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_411 <= _GEN_15639;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_412 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19c == _h_T_1) begin // @[vga.scala 64:24]
        ram_412 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19c == _T_37) begin // @[vga.scala 64:24]
        ram_412 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_412 <= _GEN_15640;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_413 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19d == _h_T_1) begin // @[vga.scala 64:24]
        ram_413 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19d == _T_37) begin // @[vga.scala 64:24]
        ram_413 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_413 <= _GEN_15641;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_414 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19e == _h_T_1) begin // @[vga.scala 64:24]
        ram_414 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19e == _T_37) begin // @[vga.scala 64:24]
        ram_414 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_414 <= _GEN_15642;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_415 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h19f == _h_T_1) begin // @[vga.scala 64:24]
        ram_415 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h19f == _T_37) begin // @[vga.scala 64:24]
        ram_415 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_415 <= _GEN_15643;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_416 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_416 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a0 == _T_37) begin // @[vga.scala 64:24]
        ram_416 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_416 <= _GEN_15644;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_417 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_417 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a1 == _T_37) begin // @[vga.scala 64:24]
        ram_417 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_417 <= _GEN_15645;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_418 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_418 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a2 == _T_37) begin // @[vga.scala 64:24]
        ram_418 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_418 <= _GEN_15646;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_419 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_419 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a3 == _T_37) begin // @[vga.scala 64:24]
        ram_419 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_419 <= _GEN_15647;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_420 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_420 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a4 == _T_37) begin // @[vga.scala 64:24]
        ram_420 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_420 <= _GEN_15648;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_421 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_421 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a5 == _T_37) begin // @[vga.scala 64:24]
        ram_421 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_421 <= _GEN_15649;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_422 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_422 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a6 == _T_37) begin // @[vga.scala 64:24]
        ram_422 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_422 <= _GEN_15650;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_423 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_423 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a7 == _T_37) begin // @[vga.scala 64:24]
        ram_423 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_423 <= _GEN_15651;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_424 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_424 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a8 == _T_37) begin // @[vga.scala 64:24]
        ram_424 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_424 <= _GEN_15652;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_425 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1a9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_425 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1a9 == _T_37) begin // @[vga.scala 64:24]
        ram_425 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_425 <= _GEN_15653;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_426 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1aa == _h_T_1) begin // @[vga.scala 64:24]
        ram_426 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1aa == _T_37) begin // @[vga.scala 64:24]
        ram_426 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_426 <= _GEN_15654;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_427 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ab == _h_T_1) begin // @[vga.scala 64:24]
        ram_427 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ab == _T_37) begin // @[vga.scala 64:24]
        ram_427 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_427 <= _GEN_15655;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_428 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ac == _h_T_1) begin // @[vga.scala 64:24]
        ram_428 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ac == _T_37) begin // @[vga.scala 64:24]
        ram_428 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_428 <= _GEN_15656;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_429 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ad == _h_T_1) begin // @[vga.scala 64:24]
        ram_429 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ad == _T_37) begin // @[vga.scala 64:24]
        ram_429 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_429 <= _GEN_15657;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_430 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ae == _h_T_1) begin // @[vga.scala 64:24]
        ram_430 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ae == _T_37) begin // @[vga.scala 64:24]
        ram_430 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_430 <= _GEN_15658;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_431 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1af == _h_T_1) begin // @[vga.scala 64:24]
        ram_431 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1af == _T_37) begin // @[vga.scala 64:24]
        ram_431 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_431 <= _GEN_15659;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_432 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_432 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b0 == _T_37) begin // @[vga.scala 64:24]
        ram_432 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_432 <= _GEN_15660;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_433 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_433 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b1 == _T_37) begin // @[vga.scala 64:24]
        ram_433 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_433 <= _GEN_15661;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_434 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_434 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b2 == _T_37) begin // @[vga.scala 64:24]
        ram_434 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_434 <= _GEN_15662;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_435 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_435 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b3 == _T_37) begin // @[vga.scala 64:24]
        ram_435 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_435 <= _GEN_15663;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_436 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_436 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b4 == _T_37) begin // @[vga.scala 64:24]
        ram_436 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_436 <= _GEN_15664;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_437 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_437 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b5 == _T_37) begin // @[vga.scala 64:24]
        ram_437 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_437 <= _GEN_15665;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_438 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_438 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b6 == _T_37) begin // @[vga.scala 64:24]
        ram_438 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_438 <= _GEN_15666;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_439 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_439 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b7 == _T_37) begin // @[vga.scala 64:24]
        ram_439 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_439 <= _GEN_15667;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_440 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_440 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b8 == _T_37) begin // @[vga.scala 64:24]
        ram_440 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_440 <= _GEN_15668;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_441 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1b9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_441 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1b9 == _T_37) begin // @[vga.scala 64:24]
        ram_441 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_441 <= _GEN_15669;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_442 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ba == _h_T_1) begin // @[vga.scala 64:24]
        ram_442 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ba == _T_37) begin // @[vga.scala 64:24]
        ram_442 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_442 <= _GEN_15670;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_443 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1bb == _h_T_1) begin // @[vga.scala 64:24]
        ram_443 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1bb == _T_37) begin // @[vga.scala 64:24]
        ram_443 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_443 <= _GEN_15671;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_444 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1bc == _h_T_1) begin // @[vga.scala 64:24]
        ram_444 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1bc == _T_37) begin // @[vga.scala 64:24]
        ram_444 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_444 <= _GEN_15672;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_445 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1bd == _h_T_1) begin // @[vga.scala 64:24]
        ram_445 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1bd == _T_37) begin // @[vga.scala 64:24]
        ram_445 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_445 <= _GEN_15673;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_446 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1be == _h_T_1) begin // @[vga.scala 64:24]
        ram_446 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1be == _T_37) begin // @[vga.scala 64:24]
        ram_446 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_446 <= _GEN_15674;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_447 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1bf == _h_T_1) begin // @[vga.scala 64:24]
        ram_447 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1bf == _T_37) begin // @[vga.scala 64:24]
        ram_447 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_447 <= _GEN_15675;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_448 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_448 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c0 == _T_37) begin // @[vga.scala 64:24]
        ram_448 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_448 <= _GEN_15676;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_449 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_449 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c1 == _T_37) begin // @[vga.scala 64:24]
        ram_449 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_449 <= _GEN_15677;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_450 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_450 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c2 == _T_37) begin // @[vga.scala 64:24]
        ram_450 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_450 <= _GEN_15678;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_451 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_451 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c3 == _T_37) begin // @[vga.scala 64:24]
        ram_451 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_451 <= _GEN_15679;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_452 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_452 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c4 == _T_37) begin // @[vga.scala 64:24]
        ram_452 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_452 <= _GEN_15680;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_453 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_453 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c5 == _T_37) begin // @[vga.scala 64:24]
        ram_453 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_453 <= _GEN_15681;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_454 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_454 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c6 == _T_37) begin // @[vga.scala 64:24]
        ram_454 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_454 <= _GEN_15682;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_455 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_455 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c7 == _T_37) begin // @[vga.scala 64:24]
        ram_455 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_455 <= _GEN_15683;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_456 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_456 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c8 == _T_37) begin // @[vga.scala 64:24]
        ram_456 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_456 <= _GEN_15684;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_457 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1c9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_457 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1c9 == _T_37) begin // @[vga.scala 64:24]
        ram_457 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_457 <= _GEN_15685;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_458 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ca == _h_T_1) begin // @[vga.scala 64:24]
        ram_458 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ca == _T_37) begin // @[vga.scala 64:24]
        ram_458 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_458 <= _GEN_15686;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_459 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1cb == _h_T_1) begin // @[vga.scala 64:24]
        ram_459 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1cb == _T_37) begin // @[vga.scala 64:24]
        ram_459 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_459 <= _GEN_15687;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_460 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1cc == _h_T_1) begin // @[vga.scala 64:24]
        ram_460 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1cc == _T_37) begin // @[vga.scala 64:24]
        ram_460 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_460 <= _GEN_15688;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_461 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1cd == _h_T_1) begin // @[vga.scala 64:24]
        ram_461 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1cd == _T_37) begin // @[vga.scala 64:24]
        ram_461 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_461 <= _GEN_15689;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_462 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ce == _h_T_1) begin // @[vga.scala 64:24]
        ram_462 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ce == _T_37) begin // @[vga.scala 64:24]
        ram_462 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_462 <= _GEN_15690;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_463 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1cf == _h_T_1) begin // @[vga.scala 64:24]
        ram_463 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1cf == _T_37) begin // @[vga.scala 64:24]
        ram_463 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_463 <= _GEN_15691;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_464 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_464 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d0 == _T_37) begin // @[vga.scala 64:24]
        ram_464 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_464 <= _GEN_15692;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_465 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_465 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d1 == _T_37) begin // @[vga.scala 64:24]
        ram_465 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_465 <= _GEN_15693;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_466 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_466 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d2 == _T_37) begin // @[vga.scala 64:24]
        ram_466 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_466 <= _GEN_15694;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_467 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_467 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d3 == _T_37) begin // @[vga.scala 64:24]
        ram_467 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_467 <= _GEN_15695;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_468 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_468 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d4 == _T_37) begin // @[vga.scala 64:24]
        ram_468 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_468 <= _GEN_15696;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_469 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_469 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d5 == _T_37) begin // @[vga.scala 64:24]
        ram_469 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_469 <= _GEN_15697;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_470 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_470 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d6 == _T_37) begin // @[vga.scala 64:24]
        ram_470 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_470 <= _GEN_15698;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_471 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_471 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d7 == _T_37) begin // @[vga.scala 64:24]
        ram_471 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_471 <= _GEN_15699;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_472 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_472 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d8 == _T_37) begin // @[vga.scala 64:24]
        ram_472 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_472 <= _GEN_15700;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_473 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1d9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_473 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1d9 == _T_37) begin // @[vga.scala 64:24]
        ram_473 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_473 <= _GEN_15701;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_474 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1da == _h_T_1) begin // @[vga.scala 64:24]
        ram_474 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1da == _T_37) begin // @[vga.scala 64:24]
        ram_474 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_474 <= _GEN_15702;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_475 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1db == _h_T_1) begin // @[vga.scala 64:24]
        ram_475 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1db == _T_37) begin // @[vga.scala 64:24]
        ram_475 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_475 <= _GEN_15703;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_476 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1dc == _h_T_1) begin // @[vga.scala 64:24]
        ram_476 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1dc == _T_37) begin // @[vga.scala 64:24]
        ram_476 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_476 <= _GEN_15704;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_477 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1dd == _h_T_1) begin // @[vga.scala 64:24]
        ram_477 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1dd == _T_37) begin // @[vga.scala 64:24]
        ram_477 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_477 <= _GEN_15705;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_478 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1de == _h_T_1) begin // @[vga.scala 64:24]
        ram_478 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1de == _T_37) begin // @[vga.scala 64:24]
        ram_478 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_478 <= _GEN_15706;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_479 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1df == _h_T_1) begin // @[vga.scala 64:24]
        ram_479 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1df == _T_37) begin // @[vga.scala 64:24]
        ram_479 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_479 <= _GEN_15707;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_480 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_480 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e0 == _T_37) begin // @[vga.scala 64:24]
        ram_480 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_480 <= _GEN_15708;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_481 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_481 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e1 == _T_37) begin // @[vga.scala 64:24]
        ram_481 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_481 <= _GEN_15709;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_482 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_482 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e2 == _T_37) begin // @[vga.scala 64:24]
        ram_482 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_482 <= _GEN_15710;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_483 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_483 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e3 == _T_37) begin // @[vga.scala 64:24]
        ram_483 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_483 <= _GEN_15711;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_484 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_484 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e4 == _T_37) begin // @[vga.scala 64:24]
        ram_484 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_484 <= _GEN_15712;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_485 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_485 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e5 == _T_37) begin // @[vga.scala 64:24]
        ram_485 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_485 <= _GEN_15713;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_486 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_486 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e6 == _T_37) begin // @[vga.scala 64:24]
        ram_486 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_486 <= _GEN_15714;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_487 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_487 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e7 == _T_37) begin // @[vga.scala 64:24]
        ram_487 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_487 <= _GEN_15715;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_488 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_488 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e8 == _T_37) begin // @[vga.scala 64:24]
        ram_488 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_488 <= _GEN_15716;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_489 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1e9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_489 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1e9 == _T_37) begin // @[vga.scala 64:24]
        ram_489 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_489 <= _GEN_15717;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_490 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ea == _h_T_1) begin // @[vga.scala 64:24]
        ram_490 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ea == _T_37) begin // @[vga.scala 64:24]
        ram_490 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_490 <= _GEN_15718;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_491 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1eb == _h_T_1) begin // @[vga.scala 64:24]
        ram_491 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1eb == _T_37) begin // @[vga.scala 64:24]
        ram_491 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_491 <= _GEN_15719;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_492 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ec == _h_T_1) begin // @[vga.scala 64:24]
        ram_492 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ec == _T_37) begin // @[vga.scala 64:24]
        ram_492 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_492 <= _GEN_15720;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_493 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ed == _h_T_1) begin // @[vga.scala 64:24]
        ram_493 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ed == _T_37) begin // @[vga.scala 64:24]
        ram_493 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_493 <= _GEN_15721;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_494 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ee == _h_T_1) begin // @[vga.scala 64:24]
        ram_494 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ee == _T_37) begin // @[vga.scala 64:24]
        ram_494 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_494 <= _GEN_15722;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_495 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ef == _h_T_1) begin // @[vga.scala 64:24]
        ram_495 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ef == _T_37) begin // @[vga.scala 64:24]
        ram_495 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_495 <= _GEN_15723;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_496 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f0 == _h_T_1) begin // @[vga.scala 64:24]
        ram_496 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f0 == _T_37) begin // @[vga.scala 64:24]
        ram_496 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_496 <= _GEN_15724;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_497 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f1 == _h_T_1) begin // @[vga.scala 64:24]
        ram_497 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f1 == _T_37) begin // @[vga.scala 64:24]
        ram_497 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_497 <= _GEN_15725;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_498 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f2 == _h_T_1) begin // @[vga.scala 64:24]
        ram_498 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f2 == _T_37) begin // @[vga.scala 64:24]
        ram_498 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_498 <= _GEN_15726;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_499 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f3 == _h_T_1) begin // @[vga.scala 64:24]
        ram_499 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f3 == _T_37) begin // @[vga.scala 64:24]
        ram_499 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_499 <= _GEN_15727;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_500 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f4 == _h_T_1) begin // @[vga.scala 64:24]
        ram_500 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f4 == _T_37) begin // @[vga.scala 64:24]
        ram_500 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_500 <= _GEN_15728;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_501 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f5 == _h_T_1) begin // @[vga.scala 64:24]
        ram_501 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f5 == _T_37) begin // @[vga.scala 64:24]
        ram_501 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_501 <= _GEN_15729;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_502 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f6 == _h_T_1) begin // @[vga.scala 64:24]
        ram_502 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f6 == _T_37) begin // @[vga.scala 64:24]
        ram_502 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_502 <= _GEN_15730;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_503 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f7 == _h_T_1) begin // @[vga.scala 64:24]
        ram_503 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f7 == _T_37) begin // @[vga.scala 64:24]
        ram_503 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_503 <= _GEN_15731;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_504 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f8 == _h_T_1) begin // @[vga.scala 64:24]
        ram_504 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f8 == _T_37) begin // @[vga.scala 64:24]
        ram_504 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_504 <= _GEN_15732;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_505 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1f9 == _h_T_1) begin // @[vga.scala 64:24]
        ram_505 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1f9 == _T_37) begin // @[vga.scala 64:24]
        ram_505 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_505 <= _GEN_15733;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_506 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1fa == _h_T_1) begin // @[vga.scala 64:24]
        ram_506 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1fa == _T_37) begin // @[vga.scala 64:24]
        ram_506 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_506 <= _GEN_15734;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_507 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1fb == _h_T_1) begin // @[vga.scala 64:24]
        ram_507 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1fb == _T_37) begin // @[vga.scala 64:24]
        ram_507 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_507 <= _GEN_15735;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_508 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1fc == _h_T_1) begin // @[vga.scala 64:24]
        ram_508 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1fc == _T_37) begin // @[vga.scala 64:24]
        ram_508 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_508 <= _GEN_15736;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_509 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1fd == _h_T_1) begin // @[vga.scala 64:24]
        ram_509 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1fd == _T_37) begin // @[vga.scala 64:24]
        ram_509 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_509 <= _GEN_15737;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_510 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1fe == _h_T_1) begin // @[vga.scala 64:24]
        ram_510 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1fe == _T_37) begin // @[vga.scala 64:24]
        ram_510 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_510 <= _GEN_15738;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_511 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h1ff == _h_T_1) begin // @[vga.scala 64:24]
        ram_511 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h1ff == _T_37) begin // @[vga.scala 64:24]
        ram_511 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_511 <= _GEN_15739;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_512 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h200 == _h_T_1) begin // @[vga.scala 64:24]
        ram_512 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h200 == _T_37) begin // @[vga.scala 64:24]
        ram_512 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_512 <= _GEN_15740;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_513 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h201 == _h_T_1) begin // @[vga.scala 64:24]
        ram_513 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h201 == _T_37) begin // @[vga.scala 64:24]
        ram_513 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_513 <= _GEN_15741;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_514 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h202 == _h_T_1) begin // @[vga.scala 64:24]
        ram_514 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h202 == _T_37) begin // @[vga.scala 64:24]
        ram_514 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_514 <= _GEN_15742;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_515 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h203 == _h_T_1) begin // @[vga.scala 64:24]
        ram_515 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h203 == _T_37) begin // @[vga.scala 64:24]
        ram_515 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_515 <= _GEN_15743;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_516 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h204 == _h_T_1) begin // @[vga.scala 64:24]
        ram_516 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h204 == _T_37) begin // @[vga.scala 64:24]
        ram_516 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_516 <= _GEN_15744;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_517 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h205 == _h_T_1) begin // @[vga.scala 64:24]
        ram_517 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h205 == _T_37) begin // @[vga.scala 64:24]
        ram_517 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_517 <= _GEN_15745;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_518 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h206 == _h_T_1) begin // @[vga.scala 64:24]
        ram_518 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h206 == _T_37) begin // @[vga.scala 64:24]
        ram_518 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_518 <= _GEN_15746;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_519 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h207 == _h_T_1) begin // @[vga.scala 64:24]
        ram_519 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h207 == _T_37) begin // @[vga.scala 64:24]
        ram_519 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_519 <= _GEN_15747;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_520 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h208 == _h_T_1) begin // @[vga.scala 64:24]
        ram_520 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h208 == _T_37) begin // @[vga.scala 64:24]
        ram_520 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_520 <= _GEN_15748;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_521 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h209 == _h_T_1) begin // @[vga.scala 64:24]
        ram_521 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h209 == _T_37) begin // @[vga.scala 64:24]
        ram_521 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_521 <= _GEN_15749;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_522 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h20a == _h_T_1) begin // @[vga.scala 64:24]
        ram_522 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h20a == _T_37) begin // @[vga.scala 64:24]
        ram_522 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_522 <= _GEN_15750;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_523 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h20b == _h_T_1) begin // @[vga.scala 64:24]
        ram_523 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h20b == _T_37) begin // @[vga.scala 64:24]
        ram_523 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_523 <= _GEN_15751;
      end
    end
    if (reset) begin // @[vga.scala 46:20]
      ram_524 <= 288'h0; // @[vga.scala 46:20]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      if (10'h20c == _h_T_1) begin // @[vga.scala 64:24]
        ram_524 <= _ram_T_441[287:0]; // @[vga.scala 64:24]
      end else if (10'h20c == _T_37) begin // @[vga.scala 64:24]
        ram_524 <= _ram_T_415[287:0]; // @[vga.scala 64:24]
      end else begin
        ram_524 <= _GEN_15752;
      end
    end
    if (reset) begin // @[vga.scala 47:18]
      h <= 10'h0; // @[vga.scala 47:18]
    end else if (h == 10'h200 & v == 9'h120) begin // @[vga.scala 54:35]
      h <= 10'h1; // @[vga.scala 55:10]
    end else if (_T_1) begin // @[vga.scala 56:26]
      h <= _h_T_1; // @[vga.scala 57:10]
    end
    if (reset) begin // @[vga.scala 48:18]
      v <= 9'h0; // @[vga.scala 48:18]
    end else if (io_now != 2'h0) begin // @[vga.scala 62:23]
      v <= _v_T_1; // @[vga.scala 66:10]
    end else if (_T_1) begin // @[vga.scala 59:20]
      v <= 9'h0; // @[vga.scala 60:10]
    end
    if (_T_40[0]) begin // @[vga.scala 69:42]
      rdwrPort <= 24'hffffff; // @[vga.scala 70:17]
    end else begin
      rdwrPort <= 24'h0; // @[vga.scala 72:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
  integer initvar;
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vga_mem_ram_MPORT_en_pipe_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  vga_mem_ram_MPORT_addr_pipe_0 = _RAND_1[11:0];
  _RAND_2 = {1{`RANDOM}};
  vga_mem_ram_MPORT_1_en_pipe_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  vga_mem_ram_MPORT_1_addr_pipe_0 = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  vga_mem_ram_MPORT_2_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vga_mem_ram_MPORT_2_addr_pipe_0 = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  vga_mem_ram_MPORT_3_en_pipe_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  vga_mem_ram_MPORT_3_addr_pipe_0 = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  vga_mem_ram_MPORT_4_en_pipe_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  vga_mem_ram_MPORT_4_addr_pipe_0 = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  vga_mem_ram_MPORT_5_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vga_mem_ram_MPORT_5_addr_pipe_0 = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  vga_mem_ram_MPORT_6_en_pipe_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  vga_mem_ram_MPORT_6_addr_pipe_0 = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  vga_mem_ram_MPORT_7_en_pipe_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  vga_mem_ram_MPORT_7_addr_pipe_0 = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  vga_mem_ram_MPORT_8_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  vga_mem_ram_MPORT_8_addr_pipe_0 = _RAND_17[11:0];
  _RAND_18 = {1{`RANDOM}};
  vga_mem_ram_MPORT_9_en_pipe_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  vga_mem_ram_MPORT_9_addr_pipe_0 = _RAND_19[11:0];
  _RAND_20 = {1{`RANDOM}};
  vga_mem_ram_MPORT_10_en_pipe_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  vga_mem_ram_MPORT_10_addr_pipe_0 = _RAND_21[11:0];
  _RAND_22 = {1{`RANDOM}};
  vga_mem_ram_MPORT_11_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  vga_mem_ram_MPORT_11_addr_pipe_0 = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  vga_mem_ram_MPORT_12_en_pipe_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  vga_mem_ram_MPORT_12_addr_pipe_0 = _RAND_25[11:0];
  _RAND_26 = {1{`RANDOM}};
  vga_mem_ram_MPORT_13_en_pipe_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vga_mem_ram_MPORT_13_addr_pipe_0 = _RAND_27[11:0];
  _RAND_28 = {1{`RANDOM}};
  vga_mem_ram_MPORT_14_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  vga_mem_ram_MPORT_14_addr_pipe_0 = _RAND_29[11:0];
  _RAND_30 = {1{`RANDOM}};
  vga_mem_ram_MPORT_15_en_pipe_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  vga_mem_ram_MPORT_15_addr_pipe_0 = _RAND_31[11:0];
  _RAND_32 = {1{`RANDOM}};
  vga_mem_ram_MPORT_16_en_pipe_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  vga_mem_ram_MPORT_16_addr_pipe_0 = _RAND_33[11:0];
  _RAND_34 = {1{`RANDOM}};
  vga_mem_ram_MPORT_17_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  vga_mem_ram_MPORT_17_addr_pipe_0 = _RAND_35[11:0];
  _RAND_36 = {1{`RANDOM}};
  vga_mem_ram_MPORT_18_en_pipe_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  vga_mem_ram_MPORT_18_addr_pipe_0 = _RAND_37[11:0];
  _RAND_38 = {1{`RANDOM}};
  vga_mem_ram_MPORT_19_en_pipe_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  vga_mem_ram_MPORT_19_addr_pipe_0 = _RAND_39[11:0];
  _RAND_40 = {1{`RANDOM}};
  vga_mem_ram_MPORT_20_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  vga_mem_ram_MPORT_20_addr_pipe_0 = _RAND_41[11:0];
  _RAND_42 = {1{`RANDOM}};
  vga_mem_ram_MPORT_21_en_pipe_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  vga_mem_ram_MPORT_21_addr_pipe_0 = _RAND_43[11:0];
  _RAND_44 = {1{`RANDOM}};
  vga_mem_ram_MPORT_22_en_pipe_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  vga_mem_ram_MPORT_22_addr_pipe_0 = _RAND_45[11:0];
  _RAND_46 = {1{`RANDOM}};
  vga_mem_ram_MPORT_23_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  vga_mem_ram_MPORT_23_addr_pipe_0 = _RAND_47[11:0];
  _RAND_48 = {1{`RANDOM}};
  vga_mem_ram_MPORT_24_en_pipe_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  vga_mem_ram_MPORT_24_addr_pipe_0 = _RAND_49[11:0];
  _RAND_50 = {1{`RANDOM}};
  vga_mem_ram_MPORT_25_en_pipe_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  vga_mem_ram_MPORT_25_addr_pipe_0 = _RAND_51[11:0];
  _RAND_52 = {1{`RANDOM}};
  vga_mem_ram_MPORT_26_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vga_mem_ram_MPORT_26_addr_pipe_0 = _RAND_53[11:0];
  _RAND_54 = {1{`RANDOM}};
  vga_mem_ram_MPORT_27_en_pipe_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  vga_mem_ram_MPORT_27_addr_pipe_0 = _RAND_55[11:0];
  _RAND_56 = {1{`RANDOM}};
  vga_mem_ram_MPORT_28_en_pipe_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  vga_mem_ram_MPORT_28_addr_pipe_0 = _RAND_57[11:0];
  _RAND_58 = {1{`RANDOM}};
  vga_mem_ram_MPORT_29_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  vga_mem_ram_MPORT_29_addr_pipe_0 = _RAND_59[11:0];
  _RAND_60 = {1{`RANDOM}};
  vga_mem_ram_MPORT_30_en_pipe_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  vga_mem_ram_MPORT_30_addr_pipe_0 = _RAND_61[11:0];
  _RAND_62 = {1{`RANDOM}};
  vga_mem_ram_MPORT_31_en_pipe_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  vga_mem_ram_MPORT_31_addr_pipe_0 = _RAND_63[11:0];
  _RAND_64 = {1{`RANDOM}};
  vga_mem_ram_MPORT_32_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  vga_mem_ram_MPORT_32_addr_pipe_0 = _RAND_65[11:0];
  _RAND_66 = {1{`RANDOM}};
  vga_mem_ram_MPORT_33_en_pipe_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  vga_mem_ram_MPORT_33_addr_pipe_0 = _RAND_67[11:0];
  _RAND_68 = {1{`RANDOM}};
  vga_mem_ram_MPORT_34_en_pipe_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  vga_mem_ram_MPORT_34_addr_pipe_0 = _RAND_69[11:0];
  _RAND_70 = {1{`RANDOM}};
  vga_mem_ram_MPORT_35_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  vga_mem_ram_MPORT_35_addr_pipe_0 = _RAND_71[11:0];
  _RAND_72 = {1{`RANDOM}};
  vga_mem_ram_MPORT_36_en_pipe_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  vga_mem_ram_MPORT_36_addr_pipe_0 = _RAND_73[11:0];
  _RAND_74 = {1{`RANDOM}};
  vga_mem_ram_MPORT_37_en_pipe_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  vga_mem_ram_MPORT_37_addr_pipe_0 = _RAND_75[11:0];
  _RAND_76 = {1{`RANDOM}};
  vga_mem_ram_MPORT_38_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  vga_mem_ram_MPORT_38_addr_pipe_0 = _RAND_77[11:0];
  _RAND_78 = {1{`RANDOM}};
  vga_mem_ram_MPORT_39_en_pipe_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  vga_mem_ram_MPORT_39_addr_pipe_0 = _RAND_79[11:0];
  _RAND_80 = {1{`RANDOM}};
  vga_mem_ram_MPORT_40_en_pipe_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  vga_mem_ram_MPORT_40_addr_pipe_0 = _RAND_81[11:0];
  _RAND_82 = {1{`RANDOM}};
  vga_mem_ram_MPORT_41_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  vga_mem_ram_MPORT_41_addr_pipe_0 = _RAND_83[11:0];
  _RAND_84 = {1{`RANDOM}};
  vga_mem_ram_MPORT_42_en_pipe_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  vga_mem_ram_MPORT_42_addr_pipe_0 = _RAND_85[11:0];
  _RAND_86 = {1{`RANDOM}};
  vga_mem_ram_MPORT_43_en_pipe_0 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  vga_mem_ram_MPORT_43_addr_pipe_0 = _RAND_87[11:0];
  _RAND_88 = {1{`RANDOM}};
  vga_mem_ram_MPORT_44_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  vga_mem_ram_MPORT_44_addr_pipe_0 = _RAND_89[11:0];
  _RAND_90 = {1{`RANDOM}};
  vga_mem_ram_MPORT_45_en_pipe_0 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  vga_mem_ram_MPORT_45_addr_pipe_0 = _RAND_91[11:0];
  _RAND_92 = {1{`RANDOM}};
  vga_mem_ram_MPORT_46_en_pipe_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  vga_mem_ram_MPORT_46_addr_pipe_0 = _RAND_93[11:0];
  _RAND_94 = {1{`RANDOM}};
  vga_mem_ram_MPORT_47_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  vga_mem_ram_MPORT_47_addr_pipe_0 = _RAND_95[11:0];
  _RAND_96 = {1{`RANDOM}};
  vga_mem_ram_MPORT_48_en_pipe_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  vga_mem_ram_MPORT_48_addr_pipe_0 = _RAND_97[11:0];
  _RAND_98 = {1{`RANDOM}};
  vga_mem_ram_MPORT_49_en_pipe_0 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  vga_mem_ram_MPORT_49_addr_pipe_0 = _RAND_99[11:0];
  _RAND_100 = {1{`RANDOM}};
  vga_mem_ram_MPORT_50_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  vga_mem_ram_MPORT_50_addr_pipe_0 = _RAND_101[11:0];
  _RAND_102 = {1{`RANDOM}};
  vga_mem_ram_MPORT_51_en_pipe_0 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  vga_mem_ram_MPORT_51_addr_pipe_0 = _RAND_103[11:0];
  _RAND_104 = {1{`RANDOM}};
  vga_mem_ram_MPORT_52_en_pipe_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  vga_mem_ram_MPORT_52_addr_pipe_0 = _RAND_105[11:0];
  _RAND_106 = {1{`RANDOM}};
  vga_mem_ram_MPORT_53_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  vga_mem_ram_MPORT_53_addr_pipe_0 = _RAND_107[11:0];
  _RAND_108 = {1{`RANDOM}};
  vga_mem_ram_MPORT_54_en_pipe_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  vga_mem_ram_MPORT_54_addr_pipe_0 = _RAND_109[11:0];
  _RAND_110 = {1{`RANDOM}};
  vga_mem_ram_MPORT_55_en_pipe_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  vga_mem_ram_MPORT_55_addr_pipe_0 = _RAND_111[11:0];
  _RAND_112 = {1{`RANDOM}};
  vga_mem_ram_MPORT_56_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  vga_mem_ram_MPORT_56_addr_pipe_0 = _RAND_113[11:0];
  _RAND_114 = {1{`RANDOM}};
  vga_mem_ram_MPORT_57_en_pipe_0 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  vga_mem_ram_MPORT_57_addr_pipe_0 = _RAND_115[11:0];
  _RAND_116 = {1{`RANDOM}};
  vga_mem_ram_MPORT_58_en_pipe_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  vga_mem_ram_MPORT_58_addr_pipe_0 = _RAND_117[11:0];
  _RAND_118 = {1{`RANDOM}};
  vga_mem_ram_MPORT_59_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  vga_mem_ram_MPORT_59_addr_pipe_0 = _RAND_119[11:0];
  _RAND_120 = {1{`RANDOM}};
  vga_mem_ram_MPORT_60_en_pipe_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  vga_mem_ram_MPORT_60_addr_pipe_0 = _RAND_121[11:0];
  _RAND_122 = {1{`RANDOM}};
  vga_mem_ram_MPORT_61_en_pipe_0 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  vga_mem_ram_MPORT_61_addr_pipe_0 = _RAND_123[11:0];
  _RAND_124 = {1{`RANDOM}};
  vga_mem_ram_MPORT_62_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  vga_mem_ram_MPORT_62_addr_pipe_0 = _RAND_125[11:0];
  _RAND_126 = {1{`RANDOM}};
  vga_mem_ram_MPORT_63_en_pipe_0 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  vga_mem_ram_MPORT_63_addr_pipe_0 = _RAND_127[11:0];
  _RAND_128 = {1{`RANDOM}};
  vga_mem_ram_MPORT_64_en_pipe_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  vga_mem_ram_MPORT_64_addr_pipe_0 = _RAND_129[11:0];
  _RAND_130 = {1{`RANDOM}};
  vga_mem_ram_MPORT_65_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  vga_mem_ram_MPORT_65_addr_pipe_0 = _RAND_131[11:0];
  _RAND_132 = {1{`RANDOM}};
  vga_mem_ram_MPORT_66_en_pipe_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  vga_mem_ram_MPORT_66_addr_pipe_0 = _RAND_133[11:0];
  _RAND_134 = {1{`RANDOM}};
  vga_mem_ram_MPORT_67_en_pipe_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  vga_mem_ram_MPORT_67_addr_pipe_0 = _RAND_135[11:0];
  _RAND_136 = {1{`RANDOM}};
  vga_mem_ram_MPORT_68_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  vga_mem_ram_MPORT_68_addr_pipe_0 = _RAND_137[11:0];
  _RAND_138 = {1{`RANDOM}};
  vga_mem_ram_MPORT_69_en_pipe_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  vga_mem_ram_MPORT_69_addr_pipe_0 = _RAND_139[11:0];
  _RAND_140 = {1{`RANDOM}};
  vga_mem_ram_MPORT_70_en_pipe_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  vga_mem_ram_MPORT_70_addr_pipe_0 = _RAND_141[11:0];
  _RAND_142 = {1{`RANDOM}};
  vga_mem_ram_MPORT_71_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  vga_mem_ram_MPORT_71_addr_pipe_0 = _RAND_143[11:0];
  _RAND_144 = {1{`RANDOM}};
  vga_mem_ram_MPORT_72_en_pipe_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  vga_mem_ram_MPORT_72_addr_pipe_0 = _RAND_145[11:0];
  _RAND_146 = {1{`RANDOM}};
  vga_mem_ram_MPORT_73_en_pipe_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  vga_mem_ram_MPORT_73_addr_pipe_0 = _RAND_147[11:0];
  _RAND_148 = {1{`RANDOM}};
  vga_mem_ram_MPORT_74_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  vga_mem_ram_MPORT_74_addr_pipe_0 = _RAND_149[11:0];
  _RAND_150 = {1{`RANDOM}};
  vga_mem_ram_MPORT_75_en_pipe_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  vga_mem_ram_MPORT_75_addr_pipe_0 = _RAND_151[11:0];
  _RAND_152 = {1{`RANDOM}};
  vga_mem_ram_MPORT_76_en_pipe_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  vga_mem_ram_MPORT_76_addr_pipe_0 = _RAND_153[11:0];
  _RAND_154 = {1{`RANDOM}};
  vga_mem_ram_MPORT_77_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  vga_mem_ram_MPORT_77_addr_pipe_0 = _RAND_155[11:0];
  _RAND_156 = {1{`RANDOM}};
  vga_mem_ram_MPORT_78_en_pipe_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  vga_mem_ram_MPORT_78_addr_pipe_0 = _RAND_157[11:0];
  _RAND_158 = {1{`RANDOM}};
  vga_mem_ram_MPORT_79_en_pipe_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  vga_mem_ram_MPORT_79_addr_pipe_0 = _RAND_159[11:0];
  _RAND_160 = {1{`RANDOM}};
  vga_mem_ram_MPORT_80_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  vga_mem_ram_MPORT_80_addr_pipe_0 = _RAND_161[11:0];
  _RAND_162 = {1{`RANDOM}};
  vga_mem_ram_MPORT_81_en_pipe_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  vga_mem_ram_MPORT_81_addr_pipe_0 = _RAND_163[11:0];
  _RAND_164 = {1{`RANDOM}};
  vga_mem_ram_MPORT_82_en_pipe_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  vga_mem_ram_MPORT_82_addr_pipe_0 = _RAND_165[11:0];
  _RAND_166 = {1{`RANDOM}};
  vga_mem_ram_MPORT_83_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  vga_mem_ram_MPORT_83_addr_pipe_0 = _RAND_167[11:0];
  _RAND_168 = {1{`RANDOM}};
  vga_mem_ram_MPORT_84_en_pipe_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  vga_mem_ram_MPORT_84_addr_pipe_0 = _RAND_169[11:0];
  _RAND_170 = {1{`RANDOM}};
  vga_mem_ram_MPORT_85_en_pipe_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  vga_mem_ram_MPORT_85_addr_pipe_0 = _RAND_171[11:0];
  _RAND_172 = {1{`RANDOM}};
  vga_mem_ram_MPORT_86_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  vga_mem_ram_MPORT_86_addr_pipe_0 = _RAND_173[11:0];
  _RAND_174 = {1{`RANDOM}};
  vga_mem_ram_MPORT_87_en_pipe_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  vga_mem_ram_MPORT_87_addr_pipe_0 = _RAND_175[11:0];
  _RAND_176 = {1{`RANDOM}};
  vga_mem_ram_MPORT_88_en_pipe_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  vga_mem_ram_MPORT_88_addr_pipe_0 = _RAND_177[11:0];
  _RAND_178 = {1{`RANDOM}};
  vga_mem_ram_MPORT_89_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  vga_mem_ram_MPORT_89_addr_pipe_0 = _RAND_179[11:0];
  _RAND_180 = {1{`RANDOM}};
  vga_mem_ram_MPORT_90_en_pipe_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  vga_mem_ram_MPORT_90_addr_pipe_0 = _RAND_181[11:0];
  _RAND_182 = {1{`RANDOM}};
  vga_mem_ram_MPORT_91_en_pipe_0 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  vga_mem_ram_MPORT_91_addr_pipe_0 = _RAND_183[11:0];
  _RAND_184 = {1{`RANDOM}};
  vga_mem_ram_MPORT_92_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  vga_mem_ram_MPORT_92_addr_pipe_0 = _RAND_185[11:0];
  _RAND_186 = {1{`RANDOM}};
  vga_mem_ram_MPORT_93_en_pipe_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  vga_mem_ram_MPORT_93_addr_pipe_0 = _RAND_187[11:0];
  _RAND_188 = {1{`RANDOM}};
  vga_mem_ram_MPORT_94_en_pipe_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  vga_mem_ram_MPORT_94_addr_pipe_0 = _RAND_189[11:0];
  _RAND_190 = {1{`RANDOM}};
  vga_mem_ram_MPORT_95_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  vga_mem_ram_MPORT_95_addr_pipe_0 = _RAND_191[11:0];
  _RAND_192 = {1{`RANDOM}};
  vga_mem_ram_MPORT_96_en_pipe_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  vga_mem_ram_MPORT_96_addr_pipe_0 = _RAND_193[11:0];
  _RAND_194 = {1{`RANDOM}};
  vga_mem_ram_MPORT_97_en_pipe_0 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  vga_mem_ram_MPORT_97_addr_pipe_0 = _RAND_195[11:0];
  _RAND_196 = {1{`RANDOM}};
  vga_mem_ram_MPORT_98_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  vga_mem_ram_MPORT_98_addr_pipe_0 = _RAND_197[11:0];
  _RAND_198 = {1{`RANDOM}};
  vga_mem_ram_MPORT_99_en_pipe_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  vga_mem_ram_MPORT_99_addr_pipe_0 = _RAND_199[11:0];
  _RAND_200 = {1{`RANDOM}};
  vga_mem_ram_MPORT_100_en_pipe_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  vga_mem_ram_MPORT_100_addr_pipe_0 = _RAND_201[11:0];
  _RAND_202 = {1{`RANDOM}};
  vga_mem_ram_MPORT_101_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  vga_mem_ram_MPORT_101_addr_pipe_0 = _RAND_203[11:0];
  _RAND_204 = {1{`RANDOM}};
  vga_mem_ram_MPORT_102_en_pipe_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  vga_mem_ram_MPORT_102_addr_pipe_0 = _RAND_205[11:0];
  _RAND_206 = {1{`RANDOM}};
  vga_mem_ram_MPORT_103_en_pipe_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  vga_mem_ram_MPORT_103_addr_pipe_0 = _RAND_207[11:0];
  _RAND_208 = {1{`RANDOM}};
  vga_mem_ram_MPORT_104_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  vga_mem_ram_MPORT_104_addr_pipe_0 = _RAND_209[11:0];
  _RAND_210 = {1{`RANDOM}};
  vga_mem_ram_MPORT_105_en_pipe_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  vga_mem_ram_MPORT_105_addr_pipe_0 = _RAND_211[11:0];
  _RAND_212 = {1{`RANDOM}};
  vga_mem_ram_MPORT_106_en_pipe_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  vga_mem_ram_MPORT_106_addr_pipe_0 = _RAND_213[11:0];
  _RAND_214 = {1{`RANDOM}};
  vga_mem_ram_MPORT_107_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  vga_mem_ram_MPORT_107_addr_pipe_0 = _RAND_215[11:0];
  _RAND_216 = {1{`RANDOM}};
  vga_mem_ram_MPORT_108_en_pipe_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  vga_mem_ram_MPORT_108_addr_pipe_0 = _RAND_217[11:0];
  _RAND_218 = {1{`RANDOM}};
  vga_mem_ram_MPORT_109_en_pipe_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  vga_mem_ram_MPORT_109_addr_pipe_0 = _RAND_219[11:0];
  _RAND_220 = {1{`RANDOM}};
  vga_mem_ram_MPORT_110_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  vga_mem_ram_MPORT_110_addr_pipe_0 = _RAND_221[11:0];
  _RAND_222 = {1{`RANDOM}};
  vga_mem_ram_MPORT_111_en_pipe_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  vga_mem_ram_MPORT_111_addr_pipe_0 = _RAND_223[11:0];
  _RAND_224 = {1{`RANDOM}};
  vga_mem_ram_MPORT_112_en_pipe_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  vga_mem_ram_MPORT_112_addr_pipe_0 = _RAND_225[11:0];
  _RAND_226 = {1{`RANDOM}};
  vga_mem_ram_MPORT_113_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  vga_mem_ram_MPORT_113_addr_pipe_0 = _RAND_227[11:0];
  _RAND_228 = {1{`RANDOM}};
  vga_mem_ram_MPORT_114_en_pipe_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  vga_mem_ram_MPORT_114_addr_pipe_0 = _RAND_229[11:0];
  _RAND_230 = {1{`RANDOM}};
  vga_mem_ram_MPORT_115_en_pipe_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  vga_mem_ram_MPORT_115_addr_pipe_0 = _RAND_231[11:0];
  _RAND_232 = {1{`RANDOM}};
  vga_mem_ram_MPORT_116_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  vga_mem_ram_MPORT_116_addr_pipe_0 = _RAND_233[11:0];
  _RAND_234 = {1{`RANDOM}};
  vga_mem_ram_MPORT_117_en_pipe_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  vga_mem_ram_MPORT_117_addr_pipe_0 = _RAND_235[11:0];
  _RAND_236 = {1{`RANDOM}};
  vga_mem_ram_MPORT_118_en_pipe_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  vga_mem_ram_MPORT_118_addr_pipe_0 = _RAND_237[11:0];
  _RAND_238 = {1{`RANDOM}};
  vga_mem_ram_MPORT_119_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  vga_mem_ram_MPORT_119_addr_pipe_0 = _RAND_239[11:0];
  _RAND_240 = {1{`RANDOM}};
  vga_mem_ram_MPORT_120_en_pipe_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  vga_mem_ram_MPORT_120_addr_pipe_0 = _RAND_241[11:0];
  _RAND_242 = {1{`RANDOM}};
  vga_mem_ram_MPORT_121_en_pipe_0 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  vga_mem_ram_MPORT_121_addr_pipe_0 = _RAND_243[11:0];
  _RAND_244 = {1{`RANDOM}};
  vga_mem_ram_MPORT_122_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  vga_mem_ram_MPORT_122_addr_pipe_0 = _RAND_245[11:0];
  _RAND_246 = {1{`RANDOM}};
  vga_mem_ram_MPORT_123_en_pipe_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  vga_mem_ram_MPORT_123_addr_pipe_0 = _RAND_247[11:0];
  _RAND_248 = {1{`RANDOM}};
  vga_mem_ram_MPORT_124_en_pipe_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  vga_mem_ram_MPORT_124_addr_pipe_0 = _RAND_249[11:0];
  _RAND_250 = {1{`RANDOM}};
  vga_mem_ram_MPORT_125_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  vga_mem_ram_MPORT_125_addr_pipe_0 = _RAND_251[11:0];
  _RAND_252 = {1{`RANDOM}};
  vga_mem_ram_MPORT_126_en_pipe_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  vga_mem_ram_MPORT_126_addr_pipe_0 = _RAND_253[11:0];
  _RAND_254 = {1{`RANDOM}};
  vga_mem_ram_MPORT_127_en_pipe_0 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  vga_mem_ram_MPORT_127_addr_pipe_0 = _RAND_255[11:0];
  _RAND_256 = {1{`RANDOM}};
  vga_mem_ram_MPORT_128_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  vga_mem_ram_MPORT_128_addr_pipe_0 = _RAND_257[11:0];
  _RAND_258 = {1{`RANDOM}};
  vga_mem_ram_MPORT_129_en_pipe_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  vga_mem_ram_MPORT_129_addr_pipe_0 = _RAND_259[11:0];
  _RAND_260 = {1{`RANDOM}};
  vga_mem_ram_MPORT_130_en_pipe_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  vga_mem_ram_MPORT_130_addr_pipe_0 = _RAND_261[11:0];
  _RAND_262 = {1{`RANDOM}};
  vga_mem_ram_MPORT_131_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  vga_mem_ram_MPORT_131_addr_pipe_0 = _RAND_263[11:0];
  _RAND_264 = {1{`RANDOM}};
  vga_mem_ram_MPORT_132_en_pipe_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  vga_mem_ram_MPORT_132_addr_pipe_0 = _RAND_265[11:0];
  _RAND_266 = {1{`RANDOM}};
  vga_mem_ram_MPORT_133_en_pipe_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  vga_mem_ram_MPORT_133_addr_pipe_0 = _RAND_267[11:0];
  _RAND_268 = {1{`RANDOM}};
  vga_mem_ram_MPORT_134_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  vga_mem_ram_MPORT_134_addr_pipe_0 = _RAND_269[11:0];
  _RAND_270 = {1{`RANDOM}};
  vga_mem_ram_MPORT_135_en_pipe_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  vga_mem_ram_MPORT_135_addr_pipe_0 = _RAND_271[11:0];
  _RAND_272 = {1{`RANDOM}};
  vga_mem_ram_MPORT_136_en_pipe_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  vga_mem_ram_MPORT_136_addr_pipe_0 = _RAND_273[11:0];
  _RAND_274 = {1{`RANDOM}};
  vga_mem_ram_MPORT_137_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  vga_mem_ram_MPORT_137_addr_pipe_0 = _RAND_275[11:0];
  _RAND_276 = {1{`RANDOM}};
  vga_mem_ram_MPORT_138_en_pipe_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  vga_mem_ram_MPORT_138_addr_pipe_0 = _RAND_277[11:0];
  _RAND_278 = {1{`RANDOM}};
  vga_mem_ram_MPORT_139_en_pipe_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  vga_mem_ram_MPORT_139_addr_pipe_0 = _RAND_279[11:0];
  _RAND_280 = {1{`RANDOM}};
  vga_mem_ram_MPORT_140_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  vga_mem_ram_MPORT_140_addr_pipe_0 = _RAND_281[11:0];
  _RAND_282 = {1{`RANDOM}};
  vga_mem_ram_MPORT_141_en_pipe_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  vga_mem_ram_MPORT_141_addr_pipe_0 = _RAND_283[11:0];
  _RAND_284 = {1{`RANDOM}};
  vga_mem_ram_MPORT_142_en_pipe_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  vga_mem_ram_MPORT_142_addr_pipe_0 = _RAND_285[11:0];
  _RAND_286 = {1{`RANDOM}};
  vga_mem_ram_MPORT_143_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  vga_mem_ram_MPORT_143_addr_pipe_0 = _RAND_287[11:0];
  _RAND_288 = {1{`RANDOM}};
  vga_mem_ram_MPORT_144_en_pipe_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  vga_mem_ram_MPORT_144_addr_pipe_0 = _RAND_289[11:0];
  _RAND_290 = {1{`RANDOM}};
  vga_mem_ram_MPORT_145_en_pipe_0 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  vga_mem_ram_MPORT_145_addr_pipe_0 = _RAND_291[11:0];
  _RAND_292 = {1{`RANDOM}};
  vga_mem_ram_MPORT_146_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  vga_mem_ram_MPORT_146_addr_pipe_0 = _RAND_293[11:0];
  _RAND_294 = {1{`RANDOM}};
  vga_mem_ram_MPORT_147_en_pipe_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  vga_mem_ram_MPORT_147_addr_pipe_0 = _RAND_295[11:0];
  _RAND_296 = {1{`RANDOM}};
  vga_mem_ram_MPORT_148_en_pipe_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  vga_mem_ram_MPORT_148_addr_pipe_0 = _RAND_297[11:0];
  _RAND_298 = {1{`RANDOM}};
  vga_mem_ram_MPORT_149_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  vga_mem_ram_MPORT_149_addr_pipe_0 = _RAND_299[11:0];
  _RAND_300 = {1{`RANDOM}};
  vga_mem_ram_MPORT_150_en_pipe_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  vga_mem_ram_MPORT_150_addr_pipe_0 = _RAND_301[11:0];
  _RAND_302 = {1{`RANDOM}};
  vga_mem_ram_MPORT_151_en_pipe_0 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  vga_mem_ram_MPORT_151_addr_pipe_0 = _RAND_303[11:0];
  _RAND_304 = {1{`RANDOM}};
  vga_mem_ram_MPORT_152_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  vga_mem_ram_MPORT_152_addr_pipe_0 = _RAND_305[11:0];
  _RAND_306 = {9{`RANDOM}};
  ram_0 = _RAND_306[287:0];
  _RAND_307 = {9{`RANDOM}};
  ram_1 = _RAND_307[287:0];
  _RAND_308 = {9{`RANDOM}};
  ram_2 = _RAND_308[287:0];
  _RAND_309 = {9{`RANDOM}};
  ram_3 = _RAND_309[287:0];
  _RAND_310 = {9{`RANDOM}};
  ram_4 = _RAND_310[287:0];
  _RAND_311 = {9{`RANDOM}};
  ram_5 = _RAND_311[287:0];
  _RAND_312 = {9{`RANDOM}};
  ram_6 = _RAND_312[287:0];
  _RAND_313 = {9{`RANDOM}};
  ram_7 = _RAND_313[287:0];
  _RAND_314 = {9{`RANDOM}};
  ram_8 = _RAND_314[287:0];
  _RAND_315 = {9{`RANDOM}};
  ram_9 = _RAND_315[287:0];
  _RAND_316 = {9{`RANDOM}};
  ram_10 = _RAND_316[287:0];
  _RAND_317 = {9{`RANDOM}};
  ram_11 = _RAND_317[287:0];
  _RAND_318 = {9{`RANDOM}};
  ram_12 = _RAND_318[287:0];
  _RAND_319 = {9{`RANDOM}};
  ram_13 = _RAND_319[287:0];
  _RAND_320 = {9{`RANDOM}};
  ram_14 = _RAND_320[287:0];
  _RAND_321 = {9{`RANDOM}};
  ram_15 = _RAND_321[287:0];
  _RAND_322 = {9{`RANDOM}};
  ram_16 = _RAND_322[287:0];
  _RAND_323 = {9{`RANDOM}};
  ram_17 = _RAND_323[287:0];
  _RAND_324 = {9{`RANDOM}};
  ram_18 = _RAND_324[287:0];
  _RAND_325 = {9{`RANDOM}};
  ram_19 = _RAND_325[287:0];
  _RAND_326 = {9{`RANDOM}};
  ram_20 = _RAND_326[287:0];
  _RAND_327 = {9{`RANDOM}};
  ram_21 = _RAND_327[287:0];
  _RAND_328 = {9{`RANDOM}};
  ram_22 = _RAND_328[287:0];
  _RAND_329 = {9{`RANDOM}};
  ram_23 = _RAND_329[287:0];
  _RAND_330 = {9{`RANDOM}};
  ram_24 = _RAND_330[287:0];
  _RAND_331 = {9{`RANDOM}};
  ram_25 = _RAND_331[287:0];
  _RAND_332 = {9{`RANDOM}};
  ram_26 = _RAND_332[287:0];
  _RAND_333 = {9{`RANDOM}};
  ram_27 = _RAND_333[287:0];
  _RAND_334 = {9{`RANDOM}};
  ram_28 = _RAND_334[287:0];
  _RAND_335 = {9{`RANDOM}};
  ram_29 = _RAND_335[287:0];
  _RAND_336 = {9{`RANDOM}};
  ram_30 = _RAND_336[287:0];
  _RAND_337 = {9{`RANDOM}};
  ram_31 = _RAND_337[287:0];
  _RAND_338 = {9{`RANDOM}};
  ram_32 = _RAND_338[287:0];
  _RAND_339 = {9{`RANDOM}};
  ram_33 = _RAND_339[287:0];
  _RAND_340 = {9{`RANDOM}};
  ram_34 = _RAND_340[287:0];
  _RAND_341 = {9{`RANDOM}};
  ram_35 = _RAND_341[287:0];
  _RAND_342 = {9{`RANDOM}};
  ram_36 = _RAND_342[287:0];
  _RAND_343 = {9{`RANDOM}};
  ram_37 = _RAND_343[287:0];
  _RAND_344 = {9{`RANDOM}};
  ram_38 = _RAND_344[287:0];
  _RAND_345 = {9{`RANDOM}};
  ram_39 = _RAND_345[287:0];
  _RAND_346 = {9{`RANDOM}};
  ram_40 = _RAND_346[287:0];
  _RAND_347 = {9{`RANDOM}};
  ram_41 = _RAND_347[287:0];
  _RAND_348 = {9{`RANDOM}};
  ram_42 = _RAND_348[287:0];
  _RAND_349 = {9{`RANDOM}};
  ram_43 = _RAND_349[287:0];
  _RAND_350 = {9{`RANDOM}};
  ram_44 = _RAND_350[287:0];
  _RAND_351 = {9{`RANDOM}};
  ram_45 = _RAND_351[287:0];
  _RAND_352 = {9{`RANDOM}};
  ram_46 = _RAND_352[287:0];
  _RAND_353 = {9{`RANDOM}};
  ram_47 = _RAND_353[287:0];
  _RAND_354 = {9{`RANDOM}};
  ram_48 = _RAND_354[287:0];
  _RAND_355 = {9{`RANDOM}};
  ram_49 = _RAND_355[287:0];
  _RAND_356 = {9{`RANDOM}};
  ram_50 = _RAND_356[287:0];
  _RAND_357 = {9{`RANDOM}};
  ram_51 = _RAND_357[287:0];
  _RAND_358 = {9{`RANDOM}};
  ram_52 = _RAND_358[287:0];
  _RAND_359 = {9{`RANDOM}};
  ram_53 = _RAND_359[287:0];
  _RAND_360 = {9{`RANDOM}};
  ram_54 = _RAND_360[287:0];
  _RAND_361 = {9{`RANDOM}};
  ram_55 = _RAND_361[287:0];
  _RAND_362 = {9{`RANDOM}};
  ram_56 = _RAND_362[287:0];
  _RAND_363 = {9{`RANDOM}};
  ram_57 = _RAND_363[287:0];
  _RAND_364 = {9{`RANDOM}};
  ram_58 = _RAND_364[287:0];
  _RAND_365 = {9{`RANDOM}};
  ram_59 = _RAND_365[287:0];
  _RAND_366 = {9{`RANDOM}};
  ram_60 = _RAND_366[287:0];
  _RAND_367 = {9{`RANDOM}};
  ram_61 = _RAND_367[287:0];
  _RAND_368 = {9{`RANDOM}};
  ram_62 = _RAND_368[287:0];
  _RAND_369 = {9{`RANDOM}};
  ram_63 = _RAND_369[287:0];
  _RAND_370 = {9{`RANDOM}};
  ram_64 = _RAND_370[287:0];
  _RAND_371 = {9{`RANDOM}};
  ram_65 = _RAND_371[287:0];
  _RAND_372 = {9{`RANDOM}};
  ram_66 = _RAND_372[287:0];
  _RAND_373 = {9{`RANDOM}};
  ram_67 = _RAND_373[287:0];
  _RAND_374 = {9{`RANDOM}};
  ram_68 = _RAND_374[287:0];
  _RAND_375 = {9{`RANDOM}};
  ram_69 = _RAND_375[287:0];
  _RAND_376 = {9{`RANDOM}};
  ram_70 = _RAND_376[287:0];
  _RAND_377 = {9{`RANDOM}};
  ram_71 = _RAND_377[287:0];
  _RAND_378 = {9{`RANDOM}};
  ram_72 = _RAND_378[287:0];
  _RAND_379 = {9{`RANDOM}};
  ram_73 = _RAND_379[287:0];
  _RAND_380 = {9{`RANDOM}};
  ram_74 = _RAND_380[287:0];
  _RAND_381 = {9{`RANDOM}};
  ram_75 = _RAND_381[287:0];
  _RAND_382 = {9{`RANDOM}};
  ram_76 = _RAND_382[287:0];
  _RAND_383 = {9{`RANDOM}};
  ram_77 = _RAND_383[287:0];
  _RAND_384 = {9{`RANDOM}};
  ram_78 = _RAND_384[287:0];
  _RAND_385 = {9{`RANDOM}};
  ram_79 = _RAND_385[287:0];
  _RAND_386 = {9{`RANDOM}};
  ram_80 = _RAND_386[287:0];
  _RAND_387 = {9{`RANDOM}};
  ram_81 = _RAND_387[287:0];
  _RAND_388 = {9{`RANDOM}};
  ram_82 = _RAND_388[287:0];
  _RAND_389 = {9{`RANDOM}};
  ram_83 = _RAND_389[287:0];
  _RAND_390 = {9{`RANDOM}};
  ram_84 = _RAND_390[287:0];
  _RAND_391 = {9{`RANDOM}};
  ram_85 = _RAND_391[287:0];
  _RAND_392 = {9{`RANDOM}};
  ram_86 = _RAND_392[287:0];
  _RAND_393 = {9{`RANDOM}};
  ram_87 = _RAND_393[287:0];
  _RAND_394 = {9{`RANDOM}};
  ram_88 = _RAND_394[287:0];
  _RAND_395 = {9{`RANDOM}};
  ram_89 = _RAND_395[287:0];
  _RAND_396 = {9{`RANDOM}};
  ram_90 = _RAND_396[287:0];
  _RAND_397 = {9{`RANDOM}};
  ram_91 = _RAND_397[287:0];
  _RAND_398 = {9{`RANDOM}};
  ram_92 = _RAND_398[287:0];
  _RAND_399 = {9{`RANDOM}};
  ram_93 = _RAND_399[287:0];
  _RAND_400 = {9{`RANDOM}};
  ram_94 = _RAND_400[287:0];
  _RAND_401 = {9{`RANDOM}};
  ram_95 = _RAND_401[287:0];
  _RAND_402 = {9{`RANDOM}};
  ram_96 = _RAND_402[287:0];
  _RAND_403 = {9{`RANDOM}};
  ram_97 = _RAND_403[287:0];
  _RAND_404 = {9{`RANDOM}};
  ram_98 = _RAND_404[287:0];
  _RAND_405 = {9{`RANDOM}};
  ram_99 = _RAND_405[287:0];
  _RAND_406 = {9{`RANDOM}};
  ram_100 = _RAND_406[287:0];
  _RAND_407 = {9{`RANDOM}};
  ram_101 = _RAND_407[287:0];
  _RAND_408 = {9{`RANDOM}};
  ram_102 = _RAND_408[287:0];
  _RAND_409 = {9{`RANDOM}};
  ram_103 = _RAND_409[287:0];
  _RAND_410 = {9{`RANDOM}};
  ram_104 = _RAND_410[287:0];
  _RAND_411 = {9{`RANDOM}};
  ram_105 = _RAND_411[287:0];
  _RAND_412 = {9{`RANDOM}};
  ram_106 = _RAND_412[287:0];
  _RAND_413 = {9{`RANDOM}};
  ram_107 = _RAND_413[287:0];
  _RAND_414 = {9{`RANDOM}};
  ram_108 = _RAND_414[287:0];
  _RAND_415 = {9{`RANDOM}};
  ram_109 = _RAND_415[287:0];
  _RAND_416 = {9{`RANDOM}};
  ram_110 = _RAND_416[287:0];
  _RAND_417 = {9{`RANDOM}};
  ram_111 = _RAND_417[287:0];
  _RAND_418 = {9{`RANDOM}};
  ram_112 = _RAND_418[287:0];
  _RAND_419 = {9{`RANDOM}};
  ram_113 = _RAND_419[287:0];
  _RAND_420 = {9{`RANDOM}};
  ram_114 = _RAND_420[287:0];
  _RAND_421 = {9{`RANDOM}};
  ram_115 = _RAND_421[287:0];
  _RAND_422 = {9{`RANDOM}};
  ram_116 = _RAND_422[287:0];
  _RAND_423 = {9{`RANDOM}};
  ram_117 = _RAND_423[287:0];
  _RAND_424 = {9{`RANDOM}};
  ram_118 = _RAND_424[287:0];
  _RAND_425 = {9{`RANDOM}};
  ram_119 = _RAND_425[287:0];
  _RAND_426 = {9{`RANDOM}};
  ram_120 = _RAND_426[287:0];
  _RAND_427 = {9{`RANDOM}};
  ram_121 = _RAND_427[287:0];
  _RAND_428 = {9{`RANDOM}};
  ram_122 = _RAND_428[287:0];
  _RAND_429 = {9{`RANDOM}};
  ram_123 = _RAND_429[287:0];
  _RAND_430 = {9{`RANDOM}};
  ram_124 = _RAND_430[287:0];
  _RAND_431 = {9{`RANDOM}};
  ram_125 = _RAND_431[287:0];
  _RAND_432 = {9{`RANDOM}};
  ram_126 = _RAND_432[287:0];
  _RAND_433 = {9{`RANDOM}};
  ram_127 = _RAND_433[287:0];
  _RAND_434 = {9{`RANDOM}};
  ram_128 = _RAND_434[287:0];
  _RAND_435 = {9{`RANDOM}};
  ram_129 = _RAND_435[287:0];
  _RAND_436 = {9{`RANDOM}};
  ram_130 = _RAND_436[287:0];
  _RAND_437 = {9{`RANDOM}};
  ram_131 = _RAND_437[287:0];
  _RAND_438 = {9{`RANDOM}};
  ram_132 = _RAND_438[287:0];
  _RAND_439 = {9{`RANDOM}};
  ram_133 = _RAND_439[287:0];
  _RAND_440 = {9{`RANDOM}};
  ram_134 = _RAND_440[287:0];
  _RAND_441 = {9{`RANDOM}};
  ram_135 = _RAND_441[287:0];
  _RAND_442 = {9{`RANDOM}};
  ram_136 = _RAND_442[287:0];
  _RAND_443 = {9{`RANDOM}};
  ram_137 = _RAND_443[287:0];
  _RAND_444 = {9{`RANDOM}};
  ram_138 = _RAND_444[287:0];
  _RAND_445 = {9{`RANDOM}};
  ram_139 = _RAND_445[287:0];
  _RAND_446 = {9{`RANDOM}};
  ram_140 = _RAND_446[287:0];
  _RAND_447 = {9{`RANDOM}};
  ram_141 = _RAND_447[287:0];
  _RAND_448 = {9{`RANDOM}};
  ram_142 = _RAND_448[287:0];
  _RAND_449 = {9{`RANDOM}};
  ram_143 = _RAND_449[287:0];
  _RAND_450 = {9{`RANDOM}};
  ram_144 = _RAND_450[287:0];
  _RAND_451 = {9{`RANDOM}};
  ram_145 = _RAND_451[287:0];
  _RAND_452 = {9{`RANDOM}};
  ram_146 = _RAND_452[287:0];
  _RAND_453 = {9{`RANDOM}};
  ram_147 = _RAND_453[287:0];
  _RAND_454 = {9{`RANDOM}};
  ram_148 = _RAND_454[287:0];
  _RAND_455 = {9{`RANDOM}};
  ram_149 = _RAND_455[287:0];
  _RAND_456 = {9{`RANDOM}};
  ram_150 = _RAND_456[287:0];
  _RAND_457 = {9{`RANDOM}};
  ram_151 = _RAND_457[287:0];
  _RAND_458 = {9{`RANDOM}};
  ram_152 = _RAND_458[287:0];
  _RAND_459 = {9{`RANDOM}};
  ram_153 = _RAND_459[287:0];
  _RAND_460 = {9{`RANDOM}};
  ram_154 = _RAND_460[287:0];
  _RAND_461 = {9{`RANDOM}};
  ram_155 = _RAND_461[287:0];
  _RAND_462 = {9{`RANDOM}};
  ram_156 = _RAND_462[287:0];
  _RAND_463 = {9{`RANDOM}};
  ram_157 = _RAND_463[287:0];
  _RAND_464 = {9{`RANDOM}};
  ram_158 = _RAND_464[287:0];
  _RAND_465 = {9{`RANDOM}};
  ram_159 = _RAND_465[287:0];
  _RAND_466 = {9{`RANDOM}};
  ram_160 = _RAND_466[287:0];
  _RAND_467 = {9{`RANDOM}};
  ram_161 = _RAND_467[287:0];
  _RAND_468 = {9{`RANDOM}};
  ram_162 = _RAND_468[287:0];
  _RAND_469 = {9{`RANDOM}};
  ram_163 = _RAND_469[287:0];
  _RAND_470 = {9{`RANDOM}};
  ram_164 = _RAND_470[287:0];
  _RAND_471 = {9{`RANDOM}};
  ram_165 = _RAND_471[287:0];
  _RAND_472 = {9{`RANDOM}};
  ram_166 = _RAND_472[287:0];
  _RAND_473 = {9{`RANDOM}};
  ram_167 = _RAND_473[287:0];
  _RAND_474 = {9{`RANDOM}};
  ram_168 = _RAND_474[287:0];
  _RAND_475 = {9{`RANDOM}};
  ram_169 = _RAND_475[287:0];
  _RAND_476 = {9{`RANDOM}};
  ram_170 = _RAND_476[287:0];
  _RAND_477 = {9{`RANDOM}};
  ram_171 = _RAND_477[287:0];
  _RAND_478 = {9{`RANDOM}};
  ram_172 = _RAND_478[287:0];
  _RAND_479 = {9{`RANDOM}};
  ram_173 = _RAND_479[287:0];
  _RAND_480 = {9{`RANDOM}};
  ram_174 = _RAND_480[287:0];
  _RAND_481 = {9{`RANDOM}};
  ram_175 = _RAND_481[287:0];
  _RAND_482 = {9{`RANDOM}};
  ram_176 = _RAND_482[287:0];
  _RAND_483 = {9{`RANDOM}};
  ram_177 = _RAND_483[287:0];
  _RAND_484 = {9{`RANDOM}};
  ram_178 = _RAND_484[287:0];
  _RAND_485 = {9{`RANDOM}};
  ram_179 = _RAND_485[287:0];
  _RAND_486 = {9{`RANDOM}};
  ram_180 = _RAND_486[287:0];
  _RAND_487 = {9{`RANDOM}};
  ram_181 = _RAND_487[287:0];
  _RAND_488 = {9{`RANDOM}};
  ram_182 = _RAND_488[287:0];
  _RAND_489 = {9{`RANDOM}};
  ram_183 = _RAND_489[287:0];
  _RAND_490 = {9{`RANDOM}};
  ram_184 = _RAND_490[287:0];
  _RAND_491 = {9{`RANDOM}};
  ram_185 = _RAND_491[287:0];
  _RAND_492 = {9{`RANDOM}};
  ram_186 = _RAND_492[287:0];
  _RAND_493 = {9{`RANDOM}};
  ram_187 = _RAND_493[287:0];
  _RAND_494 = {9{`RANDOM}};
  ram_188 = _RAND_494[287:0];
  _RAND_495 = {9{`RANDOM}};
  ram_189 = _RAND_495[287:0];
  _RAND_496 = {9{`RANDOM}};
  ram_190 = _RAND_496[287:0];
  _RAND_497 = {9{`RANDOM}};
  ram_191 = _RAND_497[287:0];
  _RAND_498 = {9{`RANDOM}};
  ram_192 = _RAND_498[287:0];
  _RAND_499 = {9{`RANDOM}};
  ram_193 = _RAND_499[287:0];
  _RAND_500 = {9{`RANDOM}};
  ram_194 = _RAND_500[287:0];
  _RAND_501 = {9{`RANDOM}};
  ram_195 = _RAND_501[287:0];
  _RAND_502 = {9{`RANDOM}};
  ram_196 = _RAND_502[287:0];
  _RAND_503 = {9{`RANDOM}};
  ram_197 = _RAND_503[287:0];
  _RAND_504 = {9{`RANDOM}};
  ram_198 = _RAND_504[287:0];
  _RAND_505 = {9{`RANDOM}};
  ram_199 = _RAND_505[287:0];
  _RAND_506 = {9{`RANDOM}};
  ram_200 = _RAND_506[287:0];
  _RAND_507 = {9{`RANDOM}};
  ram_201 = _RAND_507[287:0];
  _RAND_508 = {9{`RANDOM}};
  ram_202 = _RAND_508[287:0];
  _RAND_509 = {9{`RANDOM}};
  ram_203 = _RAND_509[287:0];
  _RAND_510 = {9{`RANDOM}};
  ram_204 = _RAND_510[287:0];
  _RAND_511 = {9{`RANDOM}};
  ram_205 = _RAND_511[287:0];
  _RAND_512 = {9{`RANDOM}};
  ram_206 = _RAND_512[287:0];
  _RAND_513 = {9{`RANDOM}};
  ram_207 = _RAND_513[287:0];
  _RAND_514 = {9{`RANDOM}};
  ram_208 = _RAND_514[287:0];
  _RAND_515 = {9{`RANDOM}};
  ram_209 = _RAND_515[287:0];
  _RAND_516 = {9{`RANDOM}};
  ram_210 = _RAND_516[287:0];
  _RAND_517 = {9{`RANDOM}};
  ram_211 = _RAND_517[287:0];
  _RAND_518 = {9{`RANDOM}};
  ram_212 = _RAND_518[287:0];
  _RAND_519 = {9{`RANDOM}};
  ram_213 = _RAND_519[287:0];
  _RAND_520 = {9{`RANDOM}};
  ram_214 = _RAND_520[287:0];
  _RAND_521 = {9{`RANDOM}};
  ram_215 = _RAND_521[287:0];
  _RAND_522 = {9{`RANDOM}};
  ram_216 = _RAND_522[287:0];
  _RAND_523 = {9{`RANDOM}};
  ram_217 = _RAND_523[287:0];
  _RAND_524 = {9{`RANDOM}};
  ram_218 = _RAND_524[287:0];
  _RAND_525 = {9{`RANDOM}};
  ram_219 = _RAND_525[287:0];
  _RAND_526 = {9{`RANDOM}};
  ram_220 = _RAND_526[287:0];
  _RAND_527 = {9{`RANDOM}};
  ram_221 = _RAND_527[287:0];
  _RAND_528 = {9{`RANDOM}};
  ram_222 = _RAND_528[287:0];
  _RAND_529 = {9{`RANDOM}};
  ram_223 = _RAND_529[287:0];
  _RAND_530 = {9{`RANDOM}};
  ram_224 = _RAND_530[287:0];
  _RAND_531 = {9{`RANDOM}};
  ram_225 = _RAND_531[287:0];
  _RAND_532 = {9{`RANDOM}};
  ram_226 = _RAND_532[287:0];
  _RAND_533 = {9{`RANDOM}};
  ram_227 = _RAND_533[287:0];
  _RAND_534 = {9{`RANDOM}};
  ram_228 = _RAND_534[287:0];
  _RAND_535 = {9{`RANDOM}};
  ram_229 = _RAND_535[287:0];
  _RAND_536 = {9{`RANDOM}};
  ram_230 = _RAND_536[287:0];
  _RAND_537 = {9{`RANDOM}};
  ram_231 = _RAND_537[287:0];
  _RAND_538 = {9{`RANDOM}};
  ram_232 = _RAND_538[287:0];
  _RAND_539 = {9{`RANDOM}};
  ram_233 = _RAND_539[287:0];
  _RAND_540 = {9{`RANDOM}};
  ram_234 = _RAND_540[287:0];
  _RAND_541 = {9{`RANDOM}};
  ram_235 = _RAND_541[287:0];
  _RAND_542 = {9{`RANDOM}};
  ram_236 = _RAND_542[287:0];
  _RAND_543 = {9{`RANDOM}};
  ram_237 = _RAND_543[287:0];
  _RAND_544 = {9{`RANDOM}};
  ram_238 = _RAND_544[287:0];
  _RAND_545 = {9{`RANDOM}};
  ram_239 = _RAND_545[287:0];
  _RAND_546 = {9{`RANDOM}};
  ram_240 = _RAND_546[287:0];
  _RAND_547 = {9{`RANDOM}};
  ram_241 = _RAND_547[287:0];
  _RAND_548 = {9{`RANDOM}};
  ram_242 = _RAND_548[287:0];
  _RAND_549 = {9{`RANDOM}};
  ram_243 = _RAND_549[287:0];
  _RAND_550 = {9{`RANDOM}};
  ram_244 = _RAND_550[287:0];
  _RAND_551 = {9{`RANDOM}};
  ram_245 = _RAND_551[287:0];
  _RAND_552 = {9{`RANDOM}};
  ram_246 = _RAND_552[287:0];
  _RAND_553 = {9{`RANDOM}};
  ram_247 = _RAND_553[287:0];
  _RAND_554 = {9{`RANDOM}};
  ram_248 = _RAND_554[287:0];
  _RAND_555 = {9{`RANDOM}};
  ram_249 = _RAND_555[287:0];
  _RAND_556 = {9{`RANDOM}};
  ram_250 = _RAND_556[287:0];
  _RAND_557 = {9{`RANDOM}};
  ram_251 = _RAND_557[287:0];
  _RAND_558 = {9{`RANDOM}};
  ram_252 = _RAND_558[287:0];
  _RAND_559 = {9{`RANDOM}};
  ram_253 = _RAND_559[287:0];
  _RAND_560 = {9{`RANDOM}};
  ram_254 = _RAND_560[287:0];
  _RAND_561 = {9{`RANDOM}};
  ram_255 = _RAND_561[287:0];
  _RAND_562 = {9{`RANDOM}};
  ram_256 = _RAND_562[287:0];
  _RAND_563 = {9{`RANDOM}};
  ram_257 = _RAND_563[287:0];
  _RAND_564 = {9{`RANDOM}};
  ram_258 = _RAND_564[287:0];
  _RAND_565 = {9{`RANDOM}};
  ram_259 = _RAND_565[287:0];
  _RAND_566 = {9{`RANDOM}};
  ram_260 = _RAND_566[287:0];
  _RAND_567 = {9{`RANDOM}};
  ram_261 = _RAND_567[287:0];
  _RAND_568 = {9{`RANDOM}};
  ram_262 = _RAND_568[287:0];
  _RAND_569 = {9{`RANDOM}};
  ram_263 = _RAND_569[287:0];
  _RAND_570 = {9{`RANDOM}};
  ram_264 = _RAND_570[287:0];
  _RAND_571 = {9{`RANDOM}};
  ram_265 = _RAND_571[287:0];
  _RAND_572 = {9{`RANDOM}};
  ram_266 = _RAND_572[287:0];
  _RAND_573 = {9{`RANDOM}};
  ram_267 = _RAND_573[287:0];
  _RAND_574 = {9{`RANDOM}};
  ram_268 = _RAND_574[287:0];
  _RAND_575 = {9{`RANDOM}};
  ram_269 = _RAND_575[287:0];
  _RAND_576 = {9{`RANDOM}};
  ram_270 = _RAND_576[287:0];
  _RAND_577 = {9{`RANDOM}};
  ram_271 = _RAND_577[287:0];
  _RAND_578 = {9{`RANDOM}};
  ram_272 = _RAND_578[287:0];
  _RAND_579 = {9{`RANDOM}};
  ram_273 = _RAND_579[287:0];
  _RAND_580 = {9{`RANDOM}};
  ram_274 = _RAND_580[287:0];
  _RAND_581 = {9{`RANDOM}};
  ram_275 = _RAND_581[287:0];
  _RAND_582 = {9{`RANDOM}};
  ram_276 = _RAND_582[287:0];
  _RAND_583 = {9{`RANDOM}};
  ram_277 = _RAND_583[287:0];
  _RAND_584 = {9{`RANDOM}};
  ram_278 = _RAND_584[287:0];
  _RAND_585 = {9{`RANDOM}};
  ram_279 = _RAND_585[287:0];
  _RAND_586 = {9{`RANDOM}};
  ram_280 = _RAND_586[287:0];
  _RAND_587 = {9{`RANDOM}};
  ram_281 = _RAND_587[287:0];
  _RAND_588 = {9{`RANDOM}};
  ram_282 = _RAND_588[287:0];
  _RAND_589 = {9{`RANDOM}};
  ram_283 = _RAND_589[287:0];
  _RAND_590 = {9{`RANDOM}};
  ram_284 = _RAND_590[287:0];
  _RAND_591 = {9{`RANDOM}};
  ram_285 = _RAND_591[287:0];
  _RAND_592 = {9{`RANDOM}};
  ram_286 = _RAND_592[287:0];
  _RAND_593 = {9{`RANDOM}};
  ram_287 = _RAND_593[287:0];
  _RAND_594 = {9{`RANDOM}};
  ram_288 = _RAND_594[287:0];
  _RAND_595 = {9{`RANDOM}};
  ram_289 = _RAND_595[287:0];
  _RAND_596 = {9{`RANDOM}};
  ram_290 = _RAND_596[287:0];
  _RAND_597 = {9{`RANDOM}};
  ram_291 = _RAND_597[287:0];
  _RAND_598 = {9{`RANDOM}};
  ram_292 = _RAND_598[287:0];
  _RAND_599 = {9{`RANDOM}};
  ram_293 = _RAND_599[287:0];
  _RAND_600 = {9{`RANDOM}};
  ram_294 = _RAND_600[287:0];
  _RAND_601 = {9{`RANDOM}};
  ram_295 = _RAND_601[287:0];
  _RAND_602 = {9{`RANDOM}};
  ram_296 = _RAND_602[287:0];
  _RAND_603 = {9{`RANDOM}};
  ram_297 = _RAND_603[287:0];
  _RAND_604 = {9{`RANDOM}};
  ram_298 = _RAND_604[287:0];
  _RAND_605 = {9{`RANDOM}};
  ram_299 = _RAND_605[287:0];
  _RAND_606 = {9{`RANDOM}};
  ram_300 = _RAND_606[287:0];
  _RAND_607 = {9{`RANDOM}};
  ram_301 = _RAND_607[287:0];
  _RAND_608 = {9{`RANDOM}};
  ram_302 = _RAND_608[287:0];
  _RAND_609 = {9{`RANDOM}};
  ram_303 = _RAND_609[287:0];
  _RAND_610 = {9{`RANDOM}};
  ram_304 = _RAND_610[287:0];
  _RAND_611 = {9{`RANDOM}};
  ram_305 = _RAND_611[287:0];
  _RAND_612 = {9{`RANDOM}};
  ram_306 = _RAND_612[287:0];
  _RAND_613 = {9{`RANDOM}};
  ram_307 = _RAND_613[287:0];
  _RAND_614 = {9{`RANDOM}};
  ram_308 = _RAND_614[287:0];
  _RAND_615 = {9{`RANDOM}};
  ram_309 = _RAND_615[287:0];
  _RAND_616 = {9{`RANDOM}};
  ram_310 = _RAND_616[287:0];
  _RAND_617 = {9{`RANDOM}};
  ram_311 = _RAND_617[287:0];
  _RAND_618 = {9{`RANDOM}};
  ram_312 = _RAND_618[287:0];
  _RAND_619 = {9{`RANDOM}};
  ram_313 = _RAND_619[287:0];
  _RAND_620 = {9{`RANDOM}};
  ram_314 = _RAND_620[287:0];
  _RAND_621 = {9{`RANDOM}};
  ram_315 = _RAND_621[287:0];
  _RAND_622 = {9{`RANDOM}};
  ram_316 = _RAND_622[287:0];
  _RAND_623 = {9{`RANDOM}};
  ram_317 = _RAND_623[287:0];
  _RAND_624 = {9{`RANDOM}};
  ram_318 = _RAND_624[287:0];
  _RAND_625 = {9{`RANDOM}};
  ram_319 = _RAND_625[287:0];
  _RAND_626 = {9{`RANDOM}};
  ram_320 = _RAND_626[287:0];
  _RAND_627 = {9{`RANDOM}};
  ram_321 = _RAND_627[287:0];
  _RAND_628 = {9{`RANDOM}};
  ram_322 = _RAND_628[287:0];
  _RAND_629 = {9{`RANDOM}};
  ram_323 = _RAND_629[287:0];
  _RAND_630 = {9{`RANDOM}};
  ram_324 = _RAND_630[287:0];
  _RAND_631 = {9{`RANDOM}};
  ram_325 = _RAND_631[287:0];
  _RAND_632 = {9{`RANDOM}};
  ram_326 = _RAND_632[287:0];
  _RAND_633 = {9{`RANDOM}};
  ram_327 = _RAND_633[287:0];
  _RAND_634 = {9{`RANDOM}};
  ram_328 = _RAND_634[287:0];
  _RAND_635 = {9{`RANDOM}};
  ram_329 = _RAND_635[287:0];
  _RAND_636 = {9{`RANDOM}};
  ram_330 = _RAND_636[287:0];
  _RAND_637 = {9{`RANDOM}};
  ram_331 = _RAND_637[287:0];
  _RAND_638 = {9{`RANDOM}};
  ram_332 = _RAND_638[287:0];
  _RAND_639 = {9{`RANDOM}};
  ram_333 = _RAND_639[287:0];
  _RAND_640 = {9{`RANDOM}};
  ram_334 = _RAND_640[287:0];
  _RAND_641 = {9{`RANDOM}};
  ram_335 = _RAND_641[287:0];
  _RAND_642 = {9{`RANDOM}};
  ram_336 = _RAND_642[287:0];
  _RAND_643 = {9{`RANDOM}};
  ram_337 = _RAND_643[287:0];
  _RAND_644 = {9{`RANDOM}};
  ram_338 = _RAND_644[287:0];
  _RAND_645 = {9{`RANDOM}};
  ram_339 = _RAND_645[287:0];
  _RAND_646 = {9{`RANDOM}};
  ram_340 = _RAND_646[287:0];
  _RAND_647 = {9{`RANDOM}};
  ram_341 = _RAND_647[287:0];
  _RAND_648 = {9{`RANDOM}};
  ram_342 = _RAND_648[287:0];
  _RAND_649 = {9{`RANDOM}};
  ram_343 = _RAND_649[287:0];
  _RAND_650 = {9{`RANDOM}};
  ram_344 = _RAND_650[287:0];
  _RAND_651 = {9{`RANDOM}};
  ram_345 = _RAND_651[287:0];
  _RAND_652 = {9{`RANDOM}};
  ram_346 = _RAND_652[287:0];
  _RAND_653 = {9{`RANDOM}};
  ram_347 = _RAND_653[287:0];
  _RAND_654 = {9{`RANDOM}};
  ram_348 = _RAND_654[287:0];
  _RAND_655 = {9{`RANDOM}};
  ram_349 = _RAND_655[287:0];
  _RAND_656 = {9{`RANDOM}};
  ram_350 = _RAND_656[287:0];
  _RAND_657 = {9{`RANDOM}};
  ram_351 = _RAND_657[287:0];
  _RAND_658 = {9{`RANDOM}};
  ram_352 = _RAND_658[287:0];
  _RAND_659 = {9{`RANDOM}};
  ram_353 = _RAND_659[287:0];
  _RAND_660 = {9{`RANDOM}};
  ram_354 = _RAND_660[287:0];
  _RAND_661 = {9{`RANDOM}};
  ram_355 = _RAND_661[287:0];
  _RAND_662 = {9{`RANDOM}};
  ram_356 = _RAND_662[287:0];
  _RAND_663 = {9{`RANDOM}};
  ram_357 = _RAND_663[287:0];
  _RAND_664 = {9{`RANDOM}};
  ram_358 = _RAND_664[287:0];
  _RAND_665 = {9{`RANDOM}};
  ram_359 = _RAND_665[287:0];
  _RAND_666 = {9{`RANDOM}};
  ram_360 = _RAND_666[287:0];
  _RAND_667 = {9{`RANDOM}};
  ram_361 = _RAND_667[287:0];
  _RAND_668 = {9{`RANDOM}};
  ram_362 = _RAND_668[287:0];
  _RAND_669 = {9{`RANDOM}};
  ram_363 = _RAND_669[287:0];
  _RAND_670 = {9{`RANDOM}};
  ram_364 = _RAND_670[287:0];
  _RAND_671 = {9{`RANDOM}};
  ram_365 = _RAND_671[287:0];
  _RAND_672 = {9{`RANDOM}};
  ram_366 = _RAND_672[287:0];
  _RAND_673 = {9{`RANDOM}};
  ram_367 = _RAND_673[287:0];
  _RAND_674 = {9{`RANDOM}};
  ram_368 = _RAND_674[287:0];
  _RAND_675 = {9{`RANDOM}};
  ram_369 = _RAND_675[287:0];
  _RAND_676 = {9{`RANDOM}};
  ram_370 = _RAND_676[287:0];
  _RAND_677 = {9{`RANDOM}};
  ram_371 = _RAND_677[287:0];
  _RAND_678 = {9{`RANDOM}};
  ram_372 = _RAND_678[287:0];
  _RAND_679 = {9{`RANDOM}};
  ram_373 = _RAND_679[287:0];
  _RAND_680 = {9{`RANDOM}};
  ram_374 = _RAND_680[287:0];
  _RAND_681 = {9{`RANDOM}};
  ram_375 = _RAND_681[287:0];
  _RAND_682 = {9{`RANDOM}};
  ram_376 = _RAND_682[287:0];
  _RAND_683 = {9{`RANDOM}};
  ram_377 = _RAND_683[287:0];
  _RAND_684 = {9{`RANDOM}};
  ram_378 = _RAND_684[287:0];
  _RAND_685 = {9{`RANDOM}};
  ram_379 = _RAND_685[287:0];
  _RAND_686 = {9{`RANDOM}};
  ram_380 = _RAND_686[287:0];
  _RAND_687 = {9{`RANDOM}};
  ram_381 = _RAND_687[287:0];
  _RAND_688 = {9{`RANDOM}};
  ram_382 = _RAND_688[287:0];
  _RAND_689 = {9{`RANDOM}};
  ram_383 = _RAND_689[287:0];
  _RAND_690 = {9{`RANDOM}};
  ram_384 = _RAND_690[287:0];
  _RAND_691 = {9{`RANDOM}};
  ram_385 = _RAND_691[287:0];
  _RAND_692 = {9{`RANDOM}};
  ram_386 = _RAND_692[287:0];
  _RAND_693 = {9{`RANDOM}};
  ram_387 = _RAND_693[287:0];
  _RAND_694 = {9{`RANDOM}};
  ram_388 = _RAND_694[287:0];
  _RAND_695 = {9{`RANDOM}};
  ram_389 = _RAND_695[287:0];
  _RAND_696 = {9{`RANDOM}};
  ram_390 = _RAND_696[287:0];
  _RAND_697 = {9{`RANDOM}};
  ram_391 = _RAND_697[287:0];
  _RAND_698 = {9{`RANDOM}};
  ram_392 = _RAND_698[287:0];
  _RAND_699 = {9{`RANDOM}};
  ram_393 = _RAND_699[287:0];
  _RAND_700 = {9{`RANDOM}};
  ram_394 = _RAND_700[287:0];
  _RAND_701 = {9{`RANDOM}};
  ram_395 = _RAND_701[287:0];
  _RAND_702 = {9{`RANDOM}};
  ram_396 = _RAND_702[287:0];
  _RAND_703 = {9{`RANDOM}};
  ram_397 = _RAND_703[287:0];
  _RAND_704 = {9{`RANDOM}};
  ram_398 = _RAND_704[287:0];
  _RAND_705 = {9{`RANDOM}};
  ram_399 = _RAND_705[287:0];
  _RAND_706 = {9{`RANDOM}};
  ram_400 = _RAND_706[287:0];
  _RAND_707 = {9{`RANDOM}};
  ram_401 = _RAND_707[287:0];
  _RAND_708 = {9{`RANDOM}};
  ram_402 = _RAND_708[287:0];
  _RAND_709 = {9{`RANDOM}};
  ram_403 = _RAND_709[287:0];
  _RAND_710 = {9{`RANDOM}};
  ram_404 = _RAND_710[287:0];
  _RAND_711 = {9{`RANDOM}};
  ram_405 = _RAND_711[287:0];
  _RAND_712 = {9{`RANDOM}};
  ram_406 = _RAND_712[287:0];
  _RAND_713 = {9{`RANDOM}};
  ram_407 = _RAND_713[287:0];
  _RAND_714 = {9{`RANDOM}};
  ram_408 = _RAND_714[287:0];
  _RAND_715 = {9{`RANDOM}};
  ram_409 = _RAND_715[287:0];
  _RAND_716 = {9{`RANDOM}};
  ram_410 = _RAND_716[287:0];
  _RAND_717 = {9{`RANDOM}};
  ram_411 = _RAND_717[287:0];
  _RAND_718 = {9{`RANDOM}};
  ram_412 = _RAND_718[287:0];
  _RAND_719 = {9{`RANDOM}};
  ram_413 = _RAND_719[287:0];
  _RAND_720 = {9{`RANDOM}};
  ram_414 = _RAND_720[287:0];
  _RAND_721 = {9{`RANDOM}};
  ram_415 = _RAND_721[287:0];
  _RAND_722 = {9{`RANDOM}};
  ram_416 = _RAND_722[287:0];
  _RAND_723 = {9{`RANDOM}};
  ram_417 = _RAND_723[287:0];
  _RAND_724 = {9{`RANDOM}};
  ram_418 = _RAND_724[287:0];
  _RAND_725 = {9{`RANDOM}};
  ram_419 = _RAND_725[287:0];
  _RAND_726 = {9{`RANDOM}};
  ram_420 = _RAND_726[287:0];
  _RAND_727 = {9{`RANDOM}};
  ram_421 = _RAND_727[287:0];
  _RAND_728 = {9{`RANDOM}};
  ram_422 = _RAND_728[287:0];
  _RAND_729 = {9{`RANDOM}};
  ram_423 = _RAND_729[287:0];
  _RAND_730 = {9{`RANDOM}};
  ram_424 = _RAND_730[287:0];
  _RAND_731 = {9{`RANDOM}};
  ram_425 = _RAND_731[287:0];
  _RAND_732 = {9{`RANDOM}};
  ram_426 = _RAND_732[287:0];
  _RAND_733 = {9{`RANDOM}};
  ram_427 = _RAND_733[287:0];
  _RAND_734 = {9{`RANDOM}};
  ram_428 = _RAND_734[287:0];
  _RAND_735 = {9{`RANDOM}};
  ram_429 = _RAND_735[287:0];
  _RAND_736 = {9{`RANDOM}};
  ram_430 = _RAND_736[287:0];
  _RAND_737 = {9{`RANDOM}};
  ram_431 = _RAND_737[287:0];
  _RAND_738 = {9{`RANDOM}};
  ram_432 = _RAND_738[287:0];
  _RAND_739 = {9{`RANDOM}};
  ram_433 = _RAND_739[287:0];
  _RAND_740 = {9{`RANDOM}};
  ram_434 = _RAND_740[287:0];
  _RAND_741 = {9{`RANDOM}};
  ram_435 = _RAND_741[287:0];
  _RAND_742 = {9{`RANDOM}};
  ram_436 = _RAND_742[287:0];
  _RAND_743 = {9{`RANDOM}};
  ram_437 = _RAND_743[287:0];
  _RAND_744 = {9{`RANDOM}};
  ram_438 = _RAND_744[287:0];
  _RAND_745 = {9{`RANDOM}};
  ram_439 = _RAND_745[287:0];
  _RAND_746 = {9{`RANDOM}};
  ram_440 = _RAND_746[287:0];
  _RAND_747 = {9{`RANDOM}};
  ram_441 = _RAND_747[287:0];
  _RAND_748 = {9{`RANDOM}};
  ram_442 = _RAND_748[287:0];
  _RAND_749 = {9{`RANDOM}};
  ram_443 = _RAND_749[287:0];
  _RAND_750 = {9{`RANDOM}};
  ram_444 = _RAND_750[287:0];
  _RAND_751 = {9{`RANDOM}};
  ram_445 = _RAND_751[287:0];
  _RAND_752 = {9{`RANDOM}};
  ram_446 = _RAND_752[287:0];
  _RAND_753 = {9{`RANDOM}};
  ram_447 = _RAND_753[287:0];
  _RAND_754 = {9{`RANDOM}};
  ram_448 = _RAND_754[287:0];
  _RAND_755 = {9{`RANDOM}};
  ram_449 = _RAND_755[287:0];
  _RAND_756 = {9{`RANDOM}};
  ram_450 = _RAND_756[287:0];
  _RAND_757 = {9{`RANDOM}};
  ram_451 = _RAND_757[287:0];
  _RAND_758 = {9{`RANDOM}};
  ram_452 = _RAND_758[287:0];
  _RAND_759 = {9{`RANDOM}};
  ram_453 = _RAND_759[287:0];
  _RAND_760 = {9{`RANDOM}};
  ram_454 = _RAND_760[287:0];
  _RAND_761 = {9{`RANDOM}};
  ram_455 = _RAND_761[287:0];
  _RAND_762 = {9{`RANDOM}};
  ram_456 = _RAND_762[287:0];
  _RAND_763 = {9{`RANDOM}};
  ram_457 = _RAND_763[287:0];
  _RAND_764 = {9{`RANDOM}};
  ram_458 = _RAND_764[287:0];
  _RAND_765 = {9{`RANDOM}};
  ram_459 = _RAND_765[287:0];
  _RAND_766 = {9{`RANDOM}};
  ram_460 = _RAND_766[287:0];
  _RAND_767 = {9{`RANDOM}};
  ram_461 = _RAND_767[287:0];
  _RAND_768 = {9{`RANDOM}};
  ram_462 = _RAND_768[287:0];
  _RAND_769 = {9{`RANDOM}};
  ram_463 = _RAND_769[287:0];
  _RAND_770 = {9{`RANDOM}};
  ram_464 = _RAND_770[287:0];
  _RAND_771 = {9{`RANDOM}};
  ram_465 = _RAND_771[287:0];
  _RAND_772 = {9{`RANDOM}};
  ram_466 = _RAND_772[287:0];
  _RAND_773 = {9{`RANDOM}};
  ram_467 = _RAND_773[287:0];
  _RAND_774 = {9{`RANDOM}};
  ram_468 = _RAND_774[287:0];
  _RAND_775 = {9{`RANDOM}};
  ram_469 = _RAND_775[287:0];
  _RAND_776 = {9{`RANDOM}};
  ram_470 = _RAND_776[287:0];
  _RAND_777 = {9{`RANDOM}};
  ram_471 = _RAND_777[287:0];
  _RAND_778 = {9{`RANDOM}};
  ram_472 = _RAND_778[287:0];
  _RAND_779 = {9{`RANDOM}};
  ram_473 = _RAND_779[287:0];
  _RAND_780 = {9{`RANDOM}};
  ram_474 = _RAND_780[287:0];
  _RAND_781 = {9{`RANDOM}};
  ram_475 = _RAND_781[287:0];
  _RAND_782 = {9{`RANDOM}};
  ram_476 = _RAND_782[287:0];
  _RAND_783 = {9{`RANDOM}};
  ram_477 = _RAND_783[287:0];
  _RAND_784 = {9{`RANDOM}};
  ram_478 = _RAND_784[287:0];
  _RAND_785 = {9{`RANDOM}};
  ram_479 = _RAND_785[287:0];
  _RAND_786 = {9{`RANDOM}};
  ram_480 = _RAND_786[287:0];
  _RAND_787 = {9{`RANDOM}};
  ram_481 = _RAND_787[287:0];
  _RAND_788 = {9{`RANDOM}};
  ram_482 = _RAND_788[287:0];
  _RAND_789 = {9{`RANDOM}};
  ram_483 = _RAND_789[287:0];
  _RAND_790 = {9{`RANDOM}};
  ram_484 = _RAND_790[287:0];
  _RAND_791 = {9{`RANDOM}};
  ram_485 = _RAND_791[287:0];
  _RAND_792 = {9{`RANDOM}};
  ram_486 = _RAND_792[287:0];
  _RAND_793 = {9{`RANDOM}};
  ram_487 = _RAND_793[287:0];
  _RAND_794 = {9{`RANDOM}};
  ram_488 = _RAND_794[287:0];
  _RAND_795 = {9{`RANDOM}};
  ram_489 = _RAND_795[287:0];
  _RAND_796 = {9{`RANDOM}};
  ram_490 = _RAND_796[287:0];
  _RAND_797 = {9{`RANDOM}};
  ram_491 = _RAND_797[287:0];
  _RAND_798 = {9{`RANDOM}};
  ram_492 = _RAND_798[287:0];
  _RAND_799 = {9{`RANDOM}};
  ram_493 = _RAND_799[287:0];
  _RAND_800 = {9{`RANDOM}};
  ram_494 = _RAND_800[287:0];
  _RAND_801 = {9{`RANDOM}};
  ram_495 = _RAND_801[287:0];
  _RAND_802 = {9{`RANDOM}};
  ram_496 = _RAND_802[287:0];
  _RAND_803 = {9{`RANDOM}};
  ram_497 = _RAND_803[287:0];
  _RAND_804 = {9{`RANDOM}};
  ram_498 = _RAND_804[287:0];
  _RAND_805 = {9{`RANDOM}};
  ram_499 = _RAND_805[287:0];
  _RAND_806 = {9{`RANDOM}};
  ram_500 = _RAND_806[287:0];
  _RAND_807 = {9{`RANDOM}};
  ram_501 = _RAND_807[287:0];
  _RAND_808 = {9{`RANDOM}};
  ram_502 = _RAND_808[287:0];
  _RAND_809 = {9{`RANDOM}};
  ram_503 = _RAND_809[287:0];
  _RAND_810 = {9{`RANDOM}};
  ram_504 = _RAND_810[287:0];
  _RAND_811 = {9{`RANDOM}};
  ram_505 = _RAND_811[287:0];
  _RAND_812 = {9{`RANDOM}};
  ram_506 = _RAND_812[287:0];
  _RAND_813 = {9{`RANDOM}};
  ram_507 = _RAND_813[287:0];
  _RAND_814 = {9{`RANDOM}};
  ram_508 = _RAND_814[287:0];
  _RAND_815 = {9{`RANDOM}};
  ram_509 = _RAND_815[287:0];
  _RAND_816 = {9{`RANDOM}};
  ram_510 = _RAND_816[287:0];
  _RAND_817 = {9{`RANDOM}};
  ram_511 = _RAND_817[287:0];
  _RAND_818 = {9{`RANDOM}};
  ram_512 = _RAND_818[287:0];
  _RAND_819 = {9{`RANDOM}};
  ram_513 = _RAND_819[287:0];
  _RAND_820 = {9{`RANDOM}};
  ram_514 = _RAND_820[287:0];
  _RAND_821 = {9{`RANDOM}};
  ram_515 = _RAND_821[287:0];
  _RAND_822 = {9{`RANDOM}};
  ram_516 = _RAND_822[287:0];
  _RAND_823 = {9{`RANDOM}};
  ram_517 = _RAND_823[287:0];
  _RAND_824 = {9{`RANDOM}};
  ram_518 = _RAND_824[287:0];
  _RAND_825 = {9{`RANDOM}};
  ram_519 = _RAND_825[287:0];
  _RAND_826 = {9{`RANDOM}};
  ram_520 = _RAND_826[287:0];
  _RAND_827 = {9{`RANDOM}};
  ram_521 = _RAND_827[287:0];
  _RAND_828 = {9{`RANDOM}};
  ram_522 = _RAND_828[287:0];
  _RAND_829 = {9{`RANDOM}};
  ram_523 = _RAND_829[287:0];
  _RAND_830 = {9{`RANDOM}};
  ram_524 = _RAND_830[287:0];
  _RAND_831 = {1{`RANDOM}};
  h = _RAND_831[9:0];
  _RAND_832 = {1{`RANDOM}};
  v = _RAND_832[8:0];
  _RAND_833 = {1{`RANDOM}};
  rdwrPort = _RAND_833[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
  $readmemh("resource/vga_font.txt", vga_mem);
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module vga(
  input        clock,
  input        reset,
  input  [1:0] io_now,
  input  [7:0] io_ascii,
  output       io_VGA_HSYNC,
  output       io_VGA_VSYNC,
  output       io_VGA_BLANK_N,
  output [7:0] io_VGA_R,
  output [7:0] io_VGA_G,
  output [7:0] io_VGA_B
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  v1_clock; // @[vga.scala 20:18]
  wire  v1_reset; // @[vga.scala 20:18]
  wire [23:0] v1_io_vga_data; // @[vga.scala 20:18]
  wire [9:0] v1_io_h_addr; // @[vga.scala 20:18]
  wire [9:0] v1_io_v_addr; // @[vga.scala 20:18]
  wire  v1_io_hsync; // @[vga.scala 20:18]
  wire  v1_io_vsync; // @[vga.scala 20:18]
  wire  v1_io_valid; // @[vga.scala 20:18]
  wire [7:0] v1_io_vga_r; // @[vga.scala 20:18]
  wire [7:0] v1_io_vga_g; // @[vga.scala 20:18]
  wire [7:0] v1_io_vga_b; // @[vga.scala 20:18]
  wire  vm_clock; // @[vga.scala 31:18]
  wire  vm_reset; // @[vga.scala 31:18]
  wire [1:0] vm_io_now; // @[vga.scala 31:18]
  wire [7:0] vm_io_ascii; // @[vga.scala 31:18]
  wire [9:0] vm_io_h_addr; // @[vga.scala 31:18]
  wire [8:0] vm_io_v_addr; // @[vga.scala 31:18]
  wire [23:0] vm_io_vga_data; // @[vga.scala 31:18]
  reg [9:0] h_addr; // @[vga.scala 16:19]
  reg [9:0] v_addr; // @[vga.scala 17:19]
  reg [23:0] vga_data; // @[vga.scala 18:21]
  vga_ctrl v1 ( // @[vga.scala 20:18]
    .clock(v1_clock),
    .reset(v1_reset),
    .io_vga_data(v1_io_vga_data),
    .io_h_addr(v1_io_h_addr),
    .io_v_addr(v1_io_v_addr),
    .io_hsync(v1_io_hsync),
    .io_vsync(v1_io_vsync),
    .io_valid(v1_io_valid),
    .io_vga_r(v1_io_vga_r),
    .io_vga_g(v1_io_vga_g),
    .io_vga_b(v1_io_vga_b)
  );
  vmem vm ( // @[vga.scala 31:18]
    .clock(vm_clock),
    .reset(vm_reset),
    .io_now(vm_io_now),
    .io_ascii(vm_io_ascii),
    .io_h_addr(vm_io_h_addr),
    .io_v_addr(vm_io_v_addr),
    .io_vga_data(vm_io_vga_data)
  );
  assign io_VGA_HSYNC = v1_io_hsync; // @[vga.scala 24:17]
  assign io_VGA_VSYNC = v1_io_vsync; // @[vga.scala 25:17]
  assign io_VGA_BLANK_N = v1_io_valid; // @[vga.scala 26:19]
  assign io_VGA_R = v1_io_vga_r; // @[vga.scala 27:13]
  assign io_VGA_G = v1_io_vga_g; // @[vga.scala 28:13]
  assign io_VGA_B = v1_io_vga_b; // @[vga.scala 29:13]
  assign v1_clock = clock;
  assign v1_reset = reset;
  assign v1_io_vga_data = vga_data; // @[vga.scala 21:19]
  assign vm_clock = clock;
  assign vm_reset = reset;
  assign vm_io_now = io_now; // @[vga.scala 32:14]
  assign vm_io_ascii = io_ascii; // @[vga.scala 33:16]
  assign vm_io_h_addr = h_addr; // @[vga.scala 34:17]
  assign vm_io_v_addr = v_addr[8:0]; // @[vga.scala 35:25]
  always @(posedge clock) begin
    h_addr <= v1_io_h_addr; // @[vga.scala 22:11]
    v_addr <= v1_io_v_addr; // @[vga.scala 23:11]
    vga_data <= vm_io_vga_data; // @[vga.scala 36:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  h_addr = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  v_addr = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  vga_data = _RAND_2[23:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input        clock,
  input        reset,
  input        io_ps2_clk,
  input        io_ps2_data,
  output       io_VGA_HSYNC,
  output       io_VGA_VSYNC,
  output       io_VGA_BLANK_N,
  output [7:0] io_VGA_R,
  output [7:0] io_VGA_G,
  output [7:0] io_VGA_B,
  output [7:0] io_bcd8seg_0,
  output [7:0] io_bcd8seg_1,
  output [7:0] io_bcd8seg_2,
  output [7:0] io_bcd8seg_3,
  output [7:0] io_bcd8seg_4,
  output [7:0] io_bcd8seg_5,
  output [7:0] io_bcd8seg_6,
  output [7:0] io_bcd8seg_7
);
  wire  PS2_clock; // @[top.scala 21:19]
  wire  PS2_reset; // @[top.scala 21:19]
  wire  PS2_io_ps2_clk; // @[top.scala 21:19]
  wire  PS2_io_ps2_data; // @[top.scala 21:19]
  wire [7:0] PS2_io_ascii; // @[top.scala 21:19]
  wire [1:0] PS2_io_now; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_0; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_1; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_2; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_3; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_4; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_5; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_6; // @[top.scala 21:19]
  wire [7:0] PS2_io_bcd8seg_7; // @[top.scala 21:19]
  wire  VGA_clock; // @[top.scala 27:19]
  wire  VGA_reset; // @[top.scala 27:19]
  wire [1:0] VGA_io_now; // @[top.scala 27:19]
  wire [7:0] VGA_io_ascii; // @[top.scala 27:19]
  wire  VGA_io_VGA_HSYNC; // @[top.scala 27:19]
  wire  VGA_io_VGA_VSYNC; // @[top.scala 27:19]
  wire  VGA_io_VGA_BLANK_N; // @[top.scala 27:19]
  wire [7:0] VGA_io_VGA_R; // @[top.scala 27:19]
  wire [7:0] VGA_io_VGA_G; // @[top.scala 27:19]
  wire [7:0] VGA_io_VGA_B; // @[top.scala 27:19]
  ps2 PS2 ( // @[top.scala 21:19]
    .clock(PS2_clock),
    .reset(PS2_reset),
    .io_ps2_clk(PS2_io_ps2_clk),
    .io_ps2_data(PS2_io_ps2_data),
    .io_ascii(PS2_io_ascii),
    .io_now(PS2_io_now),
    .io_bcd8seg_0(PS2_io_bcd8seg_0),
    .io_bcd8seg_1(PS2_io_bcd8seg_1),
    .io_bcd8seg_2(PS2_io_bcd8seg_2),
    .io_bcd8seg_3(PS2_io_bcd8seg_3),
    .io_bcd8seg_4(PS2_io_bcd8seg_4),
    .io_bcd8seg_5(PS2_io_bcd8seg_5),
    .io_bcd8seg_6(PS2_io_bcd8seg_6),
    .io_bcd8seg_7(PS2_io_bcd8seg_7)
  );
  vga VGA ( // @[top.scala 27:19]
    .clock(VGA_clock),
    .reset(VGA_reset),
    .io_now(VGA_io_now),
    .io_ascii(VGA_io_ascii),
    .io_VGA_HSYNC(VGA_io_VGA_HSYNC),
    .io_VGA_VSYNC(VGA_io_VGA_VSYNC),
    .io_VGA_BLANK_N(VGA_io_VGA_BLANK_N),
    .io_VGA_R(VGA_io_VGA_R),
    .io_VGA_G(VGA_io_VGA_G),
    .io_VGA_B(VGA_io_VGA_B)
  );
  assign io_VGA_HSYNC = VGA_io_VGA_HSYNC; // @[top.scala 30:17]
  assign io_VGA_VSYNC = VGA_io_VGA_VSYNC; // @[top.scala 31:17]
  assign io_VGA_BLANK_N = VGA_io_VGA_BLANK_N; // @[top.scala 32:19]
  assign io_VGA_R = VGA_io_VGA_R; // @[top.scala 33:13]
  assign io_VGA_G = VGA_io_VGA_G; // @[top.scala 34:13]
  assign io_VGA_B = VGA_io_VGA_B; // @[top.scala 35:13]
  assign io_bcd8seg_0 = PS2_io_bcd8seg_0; // @[top.scala 25:15]
  assign io_bcd8seg_1 = PS2_io_bcd8seg_1; // @[top.scala 25:15]
  assign io_bcd8seg_2 = PS2_io_bcd8seg_2; // @[top.scala 25:15]
  assign io_bcd8seg_3 = PS2_io_bcd8seg_3; // @[top.scala 25:15]
  assign io_bcd8seg_4 = PS2_io_bcd8seg_4; // @[top.scala 25:15]
  assign io_bcd8seg_5 = PS2_io_bcd8seg_5; // @[top.scala 25:15]
  assign io_bcd8seg_6 = PS2_io_bcd8seg_6; // @[top.scala 25:15]
  assign io_bcd8seg_7 = PS2_io_bcd8seg_7; // @[top.scala 25:15]
  assign PS2_clock = clock;
  assign PS2_reset = reset;
  assign PS2_io_ps2_clk = io_ps2_clk; // @[top.scala 23:19]
  assign PS2_io_ps2_data = io_ps2_data; // @[top.scala 24:20]
  assign VGA_clock = clock;
  assign VGA_reset = reset;
  assign VGA_io_now = PS2_io_now; // @[top.scala 29:15]
  assign VGA_io_ascii = PS2_io_ascii; // @[top.scala 28:17]
endmodule
