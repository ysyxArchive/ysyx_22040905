module ICache(
  input          clock,
  input          reset,
  output         io_in_ar_ready,
  input          io_in_ar_valid,
  input  [31:0]  io_in_ar_bits_addr,
  output         io_in_r_valid,
  output [63:0]  io_in_r_bits_data,
  input          io_mem_ar_ready,
  output         io_mem_ar_valid,
  output [31:0]  io_mem_ar_bits_addr,
  output [7:0]   io_mem_ar_bits_len,
  output         io_mem_r_ready,
  input          io_mem_r_valid,
  input  [63:0]  io_mem_r_bits_data,
  input          io_mem_r_bits_last,
  input  [127:0] io_ram_bits_Q0,
  input  [127:0] io_ram_bits_Q1,
  output         io_ram_bits_CEN,
  output         io_ram_bits_WEN,
  output [127:0] io_ram_bits_BWEN,
  output [6:0]   io_ram_bits_A,
  output [127:0] io_ram_bits_D,
  output         io_ram_bits_WAY,
  input          io_flush,
  output [63:0]  io_hitrate
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
`endif // RANDOMIZE_REG_INIT
  wire  lfsr8_clock; // @[icache.scala 54:21]
  wire  lfsr8_reset; // @[icache.scala 54:21]
  wire  lfsr8_io_en; // @[icache.scala 54:21]
  wire [7:0] lfsr8_io_out; // @[icache.scala 54:21]
  reg [41:0] cache_tag_0; // @[icache.scala 30:26]
  reg [41:0] cache_tag_1; // @[icache.scala 30:26]
  reg [41:0] cache_tag_2; // @[icache.scala 30:26]
  reg [41:0] cache_tag_3; // @[icache.scala 30:26]
  reg [41:0] cache_tag_4; // @[icache.scala 30:26]
  reg [41:0] cache_tag_5; // @[icache.scala 30:26]
  reg [41:0] cache_tag_6; // @[icache.scala 30:26]
  reg [41:0] cache_tag_7; // @[icache.scala 30:26]
  reg [41:0] cache_tag_8; // @[icache.scala 30:26]
  reg [41:0] cache_tag_9; // @[icache.scala 30:26]
  reg [41:0] cache_tag_10; // @[icache.scala 30:26]
  reg [41:0] cache_tag_11; // @[icache.scala 30:26]
  reg [41:0] cache_tag_12; // @[icache.scala 30:26]
  reg [41:0] cache_tag_13; // @[icache.scala 30:26]
  reg [41:0] cache_tag_14; // @[icache.scala 30:26]
  reg [41:0] cache_tag_15; // @[icache.scala 30:26]
  reg [41:0] cache_tag_16; // @[icache.scala 30:26]
  reg [41:0] cache_tag_17; // @[icache.scala 30:26]
  reg [41:0] cache_tag_18; // @[icache.scala 30:26]
  reg [41:0] cache_tag_19; // @[icache.scala 30:26]
  reg [41:0] cache_tag_20; // @[icache.scala 30:26]
  reg [41:0] cache_tag_21; // @[icache.scala 30:26]
  reg [41:0] cache_tag_22; // @[icache.scala 30:26]
  reg [41:0] cache_tag_23; // @[icache.scala 30:26]
  reg [41:0] cache_tag_24; // @[icache.scala 30:26]
  reg [41:0] cache_tag_25; // @[icache.scala 30:26]
  reg [41:0] cache_tag_26; // @[icache.scala 30:26]
  reg [41:0] cache_tag_27; // @[icache.scala 30:26]
  reg [41:0] cache_tag_28; // @[icache.scala 30:26]
  reg [41:0] cache_tag_29; // @[icache.scala 30:26]
  reg [41:0] cache_tag_30; // @[icache.scala 30:26]
  reg [41:0] cache_tag_31; // @[icache.scala 30:26]
  reg [41:0] cache_tag_32; // @[icache.scala 30:26]
  reg [41:0] cache_tag_33; // @[icache.scala 30:26]
  reg [41:0] cache_tag_34; // @[icache.scala 30:26]
  reg [41:0] cache_tag_35; // @[icache.scala 30:26]
  reg [41:0] cache_tag_36; // @[icache.scala 30:26]
  reg [41:0] cache_tag_37; // @[icache.scala 30:26]
  reg [41:0] cache_tag_38; // @[icache.scala 30:26]
  reg [41:0] cache_tag_39; // @[icache.scala 30:26]
  reg [41:0] cache_tag_40; // @[icache.scala 30:26]
  reg [41:0] cache_tag_41; // @[icache.scala 30:26]
  reg [41:0] cache_tag_42; // @[icache.scala 30:26]
  reg [41:0] cache_tag_43; // @[icache.scala 30:26]
  reg [41:0] cache_tag_44; // @[icache.scala 30:26]
  reg [41:0] cache_tag_45; // @[icache.scala 30:26]
  reg [41:0] cache_tag_46; // @[icache.scala 30:26]
  reg [41:0] cache_tag_47; // @[icache.scala 30:26]
  reg [41:0] cache_tag_48; // @[icache.scala 30:26]
  reg [41:0] cache_tag_49; // @[icache.scala 30:26]
  reg [41:0] cache_tag_50; // @[icache.scala 30:26]
  reg [41:0] cache_tag_51; // @[icache.scala 30:26]
  reg [41:0] cache_tag_52; // @[icache.scala 30:26]
  reg [41:0] cache_tag_53; // @[icache.scala 30:26]
  reg [41:0] cache_tag_54; // @[icache.scala 30:26]
  reg [41:0] cache_tag_55; // @[icache.scala 30:26]
  reg [41:0] cache_tag_56; // @[icache.scala 30:26]
  reg [41:0] cache_tag_57; // @[icache.scala 30:26]
  reg [41:0] cache_tag_58; // @[icache.scala 30:26]
  reg [41:0] cache_tag_59; // @[icache.scala 30:26]
  reg [41:0] cache_tag_60; // @[icache.scala 30:26]
  reg [41:0] cache_tag_61; // @[icache.scala 30:26]
  reg [41:0] cache_tag_62; // @[icache.scala 30:26]
  reg [41:0] cache_tag_63; // @[icache.scala 30:26]
  reg [41:0] cache_tag_64; // @[icache.scala 30:26]
  reg [41:0] cache_tag_65; // @[icache.scala 30:26]
  reg [41:0] cache_tag_66; // @[icache.scala 30:26]
  reg [41:0] cache_tag_67; // @[icache.scala 30:26]
  reg [41:0] cache_tag_68; // @[icache.scala 30:26]
  reg [41:0] cache_tag_69; // @[icache.scala 30:26]
  reg [41:0] cache_tag_70; // @[icache.scala 30:26]
  reg [41:0] cache_tag_71; // @[icache.scala 30:26]
  reg [41:0] cache_tag_72; // @[icache.scala 30:26]
  reg [41:0] cache_tag_73; // @[icache.scala 30:26]
  reg [41:0] cache_tag_74; // @[icache.scala 30:26]
  reg [41:0] cache_tag_75; // @[icache.scala 30:26]
  reg [41:0] cache_tag_76; // @[icache.scala 30:26]
  reg [41:0] cache_tag_77; // @[icache.scala 30:26]
  reg [41:0] cache_tag_78; // @[icache.scala 30:26]
  reg [41:0] cache_tag_79; // @[icache.scala 30:26]
  reg [41:0] cache_tag_80; // @[icache.scala 30:26]
  reg [41:0] cache_tag_81; // @[icache.scala 30:26]
  reg [41:0] cache_tag_82; // @[icache.scala 30:26]
  reg [41:0] cache_tag_83; // @[icache.scala 30:26]
  reg [41:0] cache_tag_84; // @[icache.scala 30:26]
  reg [41:0] cache_tag_85; // @[icache.scala 30:26]
  reg [41:0] cache_tag_86; // @[icache.scala 30:26]
  reg [41:0] cache_tag_87; // @[icache.scala 30:26]
  reg [41:0] cache_tag_88; // @[icache.scala 30:26]
  reg [41:0] cache_tag_89; // @[icache.scala 30:26]
  reg [41:0] cache_tag_90; // @[icache.scala 30:26]
  reg [41:0] cache_tag_91; // @[icache.scala 30:26]
  reg [41:0] cache_tag_92; // @[icache.scala 30:26]
  reg [41:0] cache_tag_93; // @[icache.scala 30:26]
  reg [41:0] cache_tag_94; // @[icache.scala 30:26]
  reg [41:0] cache_tag_95; // @[icache.scala 30:26]
  reg [41:0] cache_tag_96; // @[icache.scala 30:26]
  reg [41:0] cache_tag_97; // @[icache.scala 30:26]
  reg [41:0] cache_tag_98; // @[icache.scala 30:26]
  reg [41:0] cache_tag_99; // @[icache.scala 30:26]
  reg [41:0] cache_tag_100; // @[icache.scala 30:26]
  reg [41:0] cache_tag_101; // @[icache.scala 30:26]
  reg [41:0] cache_tag_102; // @[icache.scala 30:26]
  reg [41:0] cache_tag_103; // @[icache.scala 30:26]
  reg [41:0] cache_tag_104; // @[icache.scala 30:26]
  reg [41:0] cache_tag_105; // @[icache.scala 30:26]
  reg [41:0] cache_tag_106; // @[icache.scala 30:26]
  reg [41:0] cache_tag_107; // @[icache.scala 30:26]
  reg [41:0] cache_tag_108; // @[icache.scala 30:26]
  reg [41:0] cache_tag_109; // @[icache.scala 30:26]
  reg [41:0] cache_tag_110; // @[icache.scala 30:26]
  reg [41:0] cache_tag_111; // @[icache.scala 30:26]
  reg [41:0] cache_tag_112; // @[icache.scala 30:26]
  reg [41:0] cache_tag_113; // @[icache.scala 30:26]
  reg [41:0] cache_tag_114; // @[icache.scala 30:26]
  reg [41:0] cache_tag_115; // @[icache.scala 30:26]
  reg [41:0] cache_tag_116; // @[icache.scala 30:26]
  reg [41:0] cache_tag_117; // @[icache.scala 30:26]
  reg [41:0] cache_tag_118; // @[icache.scala 30:26]
  reg [41:0] cache_tag_119; // @[icache.scala 30:26]
  reg [41:0] cache_tag_120; // @[icache.scala 30:26]
  reg [41:0] cache_tag_121; // @[icache.scala 30:26]
  reg [41:0] cache_tag_122; // @[icache.scala 30:26]
  reg [41:0] cache_tag_123; // @[icache.scala 30:26]
  reg [41:0] cache_tag_124; // @[icache.scala 30:26]
  reg [41:0] cache_tag_125; // @[icache.scala 30:26]
  reg [41:0] cache_tag_126; // @[icache.scala 30:26]
  reg [41:0] cache_tag_127; // @[icache.scala 30:26]
  reg  valid_0_0; // @[icache.scala 31:22]
  reg  valid_0_1; // @[icache.scala 31:22]
  reg  valid_1_0; // @[icache.scala 31:22]
  reg  valid_1_1; // @[icache.scala 31:22]
  reg  valid_2_0; // @[icache.scala 31:22]
  reg  valid_2_1; // @[icache.scala 31:22]
  reg  valid_3_0; // @[icache.scala 31:22]
  reg  valid_3_1; // @[icache.scala 31:22]
  reg  valid_4_0; // @[icache.scala 31:22]
  reg  valid_4_1; // @[icache.scala 31:22]
  reg  valid_5_0; // @[icache.scala 31:22]
  reg  valid_5_1; // @[icache.scala 31:22]
  reg  valid_6_0; // @[icache.scala 31:22]
  reg  valid_6_1; // @[icache.scala 31:22]
  reg  valid_7_0; // @[icache.scala 31:22]
  reg  valid_7_1; // @[icache.scala 31:22]
  reg  valid_8_0; // @[icache.scala 31:22]
  reg  valid_8_1; // @[icache.scala 31:22]
  reg  valid_9_0; // @[icache.scala 31:22]
  reg  valid_9_1; // @[icache.scala 31:22]
  reg  valid_10_0; // @[icache.scala 31:22]
  reg  valid_10_1; // @[icache.scala 31:22]
  reg  valid_11_0; // @[icache.scala 31:22]
  reg  valid_11_1; // @[icache.scala 31:22]
  reg  valid_12_0; // @[icache.scala 31:22]
  reg  valid_12_1; // @[icache.scala 31:22]
  reg  valid_13_0; // @[icache.scala 31:22]
  reg  valid_13_1; // @[icache.scala 31:22]
  reg  valid_14_0; // @[icache.scala 31:22]
  reg  valid_14_1; // @[icache.scala 31:22]
  reg  valid_15_0; // @[icache.scala 31:22]
  reg  valid_15_1; // @[icache.scala 31:22]
  reg  valid_16_0; // @[icache.scala 31:22]
  reg  valid_16_1; // @[icache.scala 31:22]
  reg  valid_17_0; // @[icache.scala 31:22]
  reg  valid_17_1; // @[icache.scala 31:22]
  reg  valid_18_0; // @[icache.scala 31:22]
  reg  valid_18_1; // @[icache.scala 31:22]
  reg  valid_19_0; // @[icache.scala 31:22]
  reg  valid_19_1; // @[icache.scala 31:22]
  reg  valid_20_0; // @[icache.scala 31:22]
  reg  valid_20_1; // @[icache.scala 31:22]
  reg  valid_21_0; // @[icache.scala 31:22]
  reg  valid_21_1; // @[icache.scala 31:22]
  reg  valid_22_0; // @[icache.scala 31:22]
  reg  valid_22_1; // @[icache.scala 31:22]
  reg  valid_23_0; // @[icache.scala 31:22]
  reg  valid_23_1; // @[icache.scala 31:22]
  reg  valid_24_0; // @[icache.scala 31:22]
  reg  valid_24_1; // @[icache.scala 31:22]
  reg  valid_25_0; // @[icache.scala 31:22]
  reg  valid_25_1; // @[icache.scala 31:22]
  reg  valid_26_0; // @[icache.scala 31:22]
  reg  valid_26_1; // @[icache.scala 31:22]
  reg  valid_27_0; // @[icache.scala 31:22]
  reg  valid_27_1; // @[icache.scala 31:22]
  reg  valid_28_0; // @[icache.scala 31:22]
  reg  valid_28_1; // @[icache.scala 31:22]
  reg  valid_29_0; // @[icache.scala 31:22]
  reg  valid_29_1; // @[icache.scala 31:22]
  reg  valid_30_0; // @[icache.scala 31:22]
  reg  valid_30_1; // @[icache.scala 31:22]
  reg  valid_31_0; // @[icache.scala 31:22]
  reg  valid_31_1; // @[icache.scala 31:22]
  reg  valid_32_0; // @[icache.scala 31:22]
  reg  valid_32_1; // @[icache.scala 31:22]
  reg  valid_33_0; // @[icache.scala 31:22]
  reg  valid_33_1; // @[icache.scala 31:22]
  reg  valid_34_0; // @[icache.scala 31:22]
  reg  valid_34_1; // @[icache.scala 31:22]
  reg  valid_35_0; // @[icache.scala 31:22]
  reg  valid_35_1; // @[icache.scala 31:22]
  reg  valid_36_0; // @[icache.scala 31:22]
  reg  valid_36_1; // @[icache.scala 31:22]
  reg  valid_37_0; // @[icache.scala 31:22]
  reg  valid_37_1; // @[icache.scala 31:22]
  reg  valid_38_0; // @[icache.scala 31:22]
  reg  valid_38_1; // @[icache.scala 31:22]
  reg  valid_39_0; // @[icache.scala 31:22]
  reg  valid_39_1; // @[icache.scala 31:22]
  reg  valid_40_0; // @[icache.scala 31:22]
  reg  valid_40_1; // @[icache.scala 31:22]
  reg  valid_41_0; // @[icache.scala 31:22]
  reg  valid_41_1; // @[icache.scala 31:22]
  reg  valid_42_0; // @[icache.scala 31:22]
  reg  valid_42_1; // @[icache.scala 31:22]
  reg  valid_43_0; // @[icache.scala 31:22]
  reg  valid_43_1; // @[icache.scala 31:22]
  reg  valid_44_0; // @[icache.scala 31:22]
  reg  valid_44_1; // @[icache.scala 31:22]
  reg  valid_45_0; // @[icache.scala 31:22]
  reg  valid_45_1; // @[icache.scala 31:22]
  reg  valid_46_0; // @[icache.scala 31:22]
  reg  valid_46_1; // @[icache.scala 31:22]
  reg  valid_47_0; // @[icache.scala 31:22]
  reg  valid_47_1; // @[icache.scala 31:22]
  reg  valid_48_0; // @[icache.scala 31:22]
  reg  valid_48_1; // @[icache.scala 31:22]
  reg  valid_49_0; // @[icache.scala 31:22]
  reg  valid_49_1; // @[icache.scala 31:22]
  reg  valid_50_0; // @[icache.scala 31:22]
  reg  valid_50_1; // @[icache.scala 31:22]
  reg  valid_51_0; // @[icache.scala 31:22]
  reg  valid_51_1; // @[icache.scala 31:22]
  reg  valid_52_0; // @[icache.scala 31:22]
  reg  valid_52_1; // @[icache.scala 31:22]
  reg  valid_53_0; // @[icache.scala 31:22]
  reg  valid_53_1; // @[icache.scala 31:22]
  reg  valid_54_0; // @[icache.scala 31:22]
  reg  valid_54_1; // @[icache.scala 31:22]
  reg  valid_55_0; // @[icache.scala 31:22]
  reg  valid_55_1; // @[icache.scala 31:22]
  reg  valid_56_0; // @[icache.scala 31:22]
  reg  valid_56_1; // @[icache.scala 31:22]
  reg  valid_57_0; // @[icache.scala 31:22]
  reg  valid_57_1; // @[icache.scala 31:22]
  reg  valid_58_0; // @[icache.scala 31:22]
  reg  valid_58_1; // @[icache.scala 31:22]
  reg  valid_59_0; // @[icache.scala 31:22]
  reg  valid_59_1; // @[icache.scala 31:22]
  reg  valid_60_0; // @[icache.scala 31:22]
  reg  valid_60_1; // @[icache.scala 31:22]
  reg  valid_61_0; // @[icache.scala 31:22]
  reg  valid_61_1; // @[icache.scala 31:22]
  reg  valid_62_0; // @[icache.scala 31:22]
  reg  valid_62_1; // @[icache.scala 31:22]
  reg  valid_63_0; // @[icache.scala 31:22]
  reg  valid_63_1; // @[icache.scala 31:22]
  reg  valid_64_0; // @[icache.scala 31:22]
  reg  valid_64_1; // @[icache.scala 31:22]
  reg  valid_65_0; // @[icache.scala 31:22]
  reg  valid_65_1; // @[icache.scala 31:22]
  reg  valid_66_0; // @[icache.scala 31:22]
  reg  valid_66_1; // @[icache.scala 31:22]
  reg  valid_67_0; // @[icache.scala 31:22]
  reg  valid_67_1; // @[icache.scala 31:22]
  reg  valid_68_0; // @[icache.scala 31:22]
  reg  valid_68_1; // @[icache.scala 31:22]
  reg  valid_69_0; // @[icache.scala 31:22]
  reg  valid_69_1; // @[icache.scala 31:22]
  reg  valid_70_0; // @[icache.scala 31:22]
  reg  valid_70_1; // @[icache.scala 31:22]
  reg  valid_71_0; // @[icache.scala 31:22]
  reg  valid_71_1; // @[icache.scala 31:22]
  reg  valid_72_0; // @[icache.scala 31:22]
  reg  valid_72_1; // @[icache.scala 31:22]
  reg  valid_73_0; // @[icache.scala 31:22]
  reg  valid_73_1; // @[icache.scala 31:22]
  reg  valid_74_0; // @[icache.scala 31:22]
  reg  valid_74_1; // @[icache.scala 31:22]
  reg  valid_75_0; // @[icache.scala 31:22]
  reg  valid_75_1; // @[icache.scala 31:22]
  reg  valid_76_0; // @[icache.scala 31:22]
  reg  valid_76_1; // @[icache.scala 31:22]
  reg  valid_77_0; // @[icache.scala 31:22]
  reg  valid_77_1; // @[icache.scala 31:22]
  reg  valid_78_0; // @[icache.scala 31:22]
  reg  valid_78_1; // @[icache.scala 31:22]
  reg  valid_79_0; // @[icache.scala 31:22]
  reg  valid_79_1; // @[icache.scala 31:22]
  reg  valid_80_0; // @[icache.scala 31:22]
  reg  valid_80_1; // @[icache.scala 31:22]
  reg  valid_81_0; // @[icache.scala 31:22]
  reg  valid_81_1; // @[icache.scala 31:22]
  reg  valid_82_0; // @[icache.scala 31:22]
  reg  valid_82_1; // @[icache.scala 31:22]
  reg  valid_83_0; // @[icache.scala 31:22]
  reg  valid_83_1; // @[icache.scala 31:22]
  reg  valid_84_0; // @[icache.scala 31:22]
  reg  valid_84_1; // @[icache.scala 31:22]
  reg  valid_85_0; // @[icache.scala 31:22]
  reg  valid_85_1; // @[icache.scala 31:22]
  reg  valid_86_0; // @[icache.scala 31:22]
  reg  valid_86_1; // @[icache.scala 31:22]
  reg  valid_87_0; // @[icache.scala 31:22]
  reg  valid_87_1; // @[icache.scala 31:22]
  reg  valid_88_0; // @[icache.scala 31:22]
  reg  valid_88_1; // @[icache.scala 31:22]
  reg  valid_89_0; // @[icache.scala 31:22]
  reg  valid_89_1; // @[icache.scala 31:22]
  reg  valid_90_0; // @[icache.scala 31:22]
  reg  valid_90_1; // @[icache.scala 31:22]
  reg  valid_91_0; // @[icache.scala 31:22]
  reg  valid_91_1; // @[icache.scala 31:22]
  reg  valid_92_0; // @[icache.scala 31:22]
  reg  valid_92_1; // @[icache.scala 31:22]
  reg  valid_93_0; // @[icache.scala 31:22]
  reg  valid_93_1; // @[icache.scala 31:22]
  reg  valid_94_0; // @[icache.scala 31:22]
  reg  valid_94_1; // @[icache.scala 31:22]
  reg  valid_95_0; // @[icache.scala 31:22]
  reg  valid_95_1; // @[icache.scala 31:22]
  reg  valid_96_0; // @[icache.scala 31:22]
  reg  valid_96_1; // @[icache.scala 31:22]
  reg  valid_97_0; // @[icache.scala 31:22]
  reg  valid_97_1; // @[icache.scala 31:22]
  reg  valid_98_0; // @[icache.scala 31:22]
  reg  valid_98_1; // @[icache.scala 31:22]
  reg  valid_99_0; // @[icache.scala 31:22]
  reg  valid_99_1; // @[icache.scala 31:22]
  reg  valid_100_0; // @[icache.scala 31:22]
  reg  valid_100_1; // @[icache.scala 31:22]
  reg  valid_101_0; // @[icache.scala 31:22]
  reg  valid_101_1; // @[icache.scala 31:22]
  reg  valid_102_0; // @[icache.scala 31:22]
  reg  valid_102_1; // @[icache.scala 31:22]
  reg  valid_103_0; // @[icache.scala 31:22]
  reg  valid_103_1; // @[icache.scala 31:22]
  reg  valid_104_0; // @[icache.scala 31:22]
  reg  valid_104_1; // @[icache.scala 31:22]
  reg  valid_105_0; // @[icache.scala 31:22]
  reg  valid_105_1; // @[icache.scala 31:22]
  reg  valid_106_0; // @[icache.scala 31:22]
  reg  valid_106_1; // @[icache.scala 31:22]
  reg  valid_107_0; // @[icache.scala 31:22]
  reg  valid_107_1; // @[icache.scala 31:22]
  reg  valid_108_0; // @[icache.scala 31:22]
  reg  valid_108_1; // @[icache.scala 31:22]
  reg  valid_109_0; // @[icache.scala 31:22]
  reg  valid_109_1; // @[icache.scala 31:22]
  reg  valid_110_0; // @[icache.scala 31:22]
  reg  valid_110_1; // @[icache.scala 31:22]
  reg  valid_111_0; // @[icache.scala 31:22]
  reg  valid_111_1; // @[icache.scala 31:22]
  reg  valid_112_0; // @[icache.scala 31:22]
  reg  valid_112_1; // @[icache.scala 31:22]
  reg  valid_113_0; // @[icache.scala 31:22]
  reg  valid_113_1; // @[icache.scala 31:22]
  reg  valid_114_0; // @[icache.scala 31:22]
  reg  valid_114_1; // @[icache.scala 31:22]
  reg  valid_115_0; // @[icache.scala 31:22]
  reg  valid_115_1; // @[icache.scala 31:22]
  reg  valid_116_0; // @[icache.scala 31:22]
  reg  valid_116_1; // @[icache.scala 31:22]
  reg  valid_117_0; // @[icache.scala 31:22]
  reg  valid_117_1; // @[icache.scala 31:22]
  reg  valid_118_0; // @[icache.scala 31:22]
  reg  valid_118_1; // @[icache.scala 31:22]
  reg  valid_119_0; // @[icache.scala 31:22]
  reg  valid_119_1; // @[icache.scala 31:22]
  reg  valid_120_0; // @[icache.scala 31:22]
  reg  valid_120_1; // @[icache.scala 31:22]
  reg  valid_121_0; // @[icache.scala 31:22]
  reg  valid_121_1; // @[icache.scala 31:22]
  reg  valid_122_0; // @[icache.scala 31:22]
  reg  valid_122_1; // @[icache.scala 31:22]
  reg  valid_123_0; // @[icache.scala 31:22]
  reg  valid_123_1; // @[icache.scala 31:22]
  reg  valid_124_0; // @[icache.scala 31:22]
  reg  valid_124_1; // @[icache.scala 31:22]
  reg  valid_125_0; // @[icache.scala 31:22]
  reg  valid_125_1; // @[icache.scala 31:22]
  reg  valid_126_0; // @[icache.scala 31:22]
  reg  valid_126_1; // @[icache.scala 31:22]
  reg  valid_127_0; // @[icache.scala 31:22]
  reg  valid_127_1; // @[icache.scala 31:22]
  reg [1:0] state; // @[icache.scala 36:22]
  wire  req = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 52:35]
  reg [31:0] addr; // @[icache.scala 39:21]
  reg  uncache; // @[icache.scala 40:24]
  wire [20:0] tag = addr[31:11]; // @[icache.scala 41:17]
  wire [6:0] offset = {addr[3:0], 3'h0}; // @[icache.scala 42:42]
  wire [6:0] idx = addr[10:4]; // @[icache.scala 43:17]
  wire [41:0] _GEN_1 = 7'h1 == idx ? cache_tag_1 : cache_tag_0; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_2 = 7'h2 == idx ? cache_tag_2 : _GEN_1; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_3 = 7'h3 == idx ? cache_tag_3 : _GEN_2; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_4 = 7'h4 == idx ? cache_tag_4 : _GEN_3; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_5 = 7'h5 == idx ? cache_tag_5 : _GEN_4; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_6 = 7'h6 == idx ? cache_tag_6 : _GEN_5; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_7 = 7'h7 == idx ? cache_tag_7 : _GEN_6; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_8 = 7'h8 == idx ? cache_tag_8 : _GEN_7; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_9 = 7'h9 == idx ? cache_tag_9 : _GEN_8; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_10 = 7'ha == idx ? cache_tag_10 : _GEN_9; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_11 = 7'hb == idx ? cache_tag_11 : _GEN_10; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_12 = 7'hc == idx ? cache_tag_12 : _GEN_11; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_13 = 7'hd == idx ? cache_tag_13 : _GEN_12; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_14 = 7'he == idx ? cache_tag_14 : _GEN_13; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_15 = 7'hf == idx ? cache_tag_15 : _GEN_14; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_16 = 7'h10 == idx ? cache_tag_16 : _GEN_15; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_17 = 7'h11 == idx ? cache_tag_17 : _GEN_16; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_18 = 7'h12 == idx ? cache_tag_18 : _GEN_17; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_19 = 7'h13 == idx ? cache_tag_19 : _GEN_18; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_20 = 7'h14 == idx ? cache_tag_20 : _GEN_19; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_21 = 7'h15 == idx ? cache_tag_21 : _GEN_20; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_22 = 7'h16 == idx ? cache_tag_22 : _GEN_21; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_23 = 7'h17 == idx ? cache_tag_23 : _GEN_22; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_24 = 7'h18 == idx ? cache_tag_24 : _GEN_23; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_25 = 7'h19 == idx ? cache_tag_25 : _GEN_24; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_26 = 7'h1a == idx ? cache_tag_26 : _GEN_25; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_27 = 7'h1b == idx ? cache_tag_27 : _GEN_26; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_28 = 7'h1c == idx ? cache_tag_28 : _GEN_27; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_29 = 7'h1d == idx ? cache_tag_29 : _GEN_28; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_30 = 7'h1e == idx ? cache_tag_30 : _GEN_29; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_31 = 7'h1f == idx ? cache_tag_31 : _GEN_30; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_32 = 7'h20 == idx ? cache_tag_32 : _GEN_31; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_33 = 7'h21 == idx ? cache_tag_33 : _GEN_32; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_34 = 7'h22 == idx ? cache_tag_34 : _GEN_33; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_35 = 7'h23 == idx ? cache_tag_35 : _GEN_34; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_36 = 7'h24 == idx ? cache_tag_36 : _GEN_35; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_37 = 7'h25 == idx ? cache_tag_37 : _GEN_36; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_38 = 7'h26 == idx ? cache_tag_38 : _GEN_37; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_39 = 7'h27 == idx ? cache_tag_39 : _GEN_38; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_40 = 7'h28 == idx ? cache_tag_40 : _GEN_39; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_41 = 7'h29 == idx ? cache_tag_41 : _GEN_40; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_42 = 7'h2a == idx ? cache_tag_42 : _GEN_41; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_43 = 7'h2b == idx ? cache_tag_43 : _GEN_42; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_44 = 7'h2c == idx ? cache_tag_44 : _GEN_43; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_45 = 7'h2d == idx ? cache_tag_45 : _GEN_44; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_46 = 7'h2e == idx ? cache_tag_46 : _GEN_45; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_47 = 7'h2f == idx ? cache_tag_47 : _GEN_46; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_48 = 7'h30 == idx ? cache_tag_48 : _GEN_47; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_49 = 7'h31 == idx ? cache_tag_49 : _GEN_48; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_50 = 7'h32 == idx ? cache_tag_50 : _GEN_49; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_51 = 7'h33 == idx ? cache_tag_51 : _GEN_50; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_52 = 7'h34 == idx ? cache_tag_52 : _GEN_51; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_53 = 7'h35 == idx ? cache_tag_53 : _GEN_52; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_54 = 7'h36 == idx ? cache_tag_54 : _GEN_53; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_55 = 7'h37 == idx ? cache_tag_55 : _GEN_54; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_56 = 7'h38 == idx ? cache_tag_56 : _GEN_55; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_57 = 7'h39 == idx ? cache_tag_57 : _GEN_56; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_58 = 7'h3a == idx ? cache_tag_58 : _GEN_57; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_59 = 7'h3b == idx ? cache_tag_59 : _GEN_58; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_60 = 7'h3c == idx ? cache_tag_60 : _GEN_59; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_61 = 7'h3d == idx ? cache_tag_61 : _GEN_60; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_62 = 7'h3e == idx ? cache_tag_62 : _GEN_61; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_63 = 7'h3f == idx ? cache_tag_63 : _GEN_62; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_64 = 7'h40 == idx ? cache_tag_64 : _GEN_63; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_65 = 7'h41 == idx ? cache_tag_65 : _GEN_64; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_66 = 7'h42 == idx ? cache_tag_66 : _GEN_65; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_67 = 7'h43 == idx ? cache_tag_67 : _GEN_66; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_68 = 7'h44 == idx ? cache_tag_68 : _GEN_67; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_69 = 7'h45 == idx ? cache_tag_69 : _GEN_68; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_70 = 7'h46 == idx ? cache_tag_70 : _GEN_69; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_71 = 7'h47 == idx ? cache_tag_71 : _GEN_70; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_72 = 7'h48 == idx ? cache_tag_72 : _GEN_71; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_73 = 7'h49 == idx ? cache_tag_73 : _GEN_72; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_74 = 7'h4a == idx ? cache_tag_74 : _GEN_73; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_75 = 7'h4b == idx ? cache_tag_75 : _GEN_74; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_76 = 7'h4c == idx ? cache_tag_76 : _GEN_75; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_77 = 7'h4d == idx ? cache_tag_77 : _GEN_76; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_78 = 7'h4e == idx ? cache_tag_78 : _GEN_77; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_79 = 7'h4f == idx ? cache_tag_79 : _GEN_78; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_80 = 7'h50 == idx ? cache_tag_80 : _GEN_79; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_81 = 7'h51 == idx ? cache_tag_81 : _GEN_80; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_82 = 7'h52 == idx ? cache_tag_82 : _GEN_81; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_83 = 7'h53 == idx ? cache_tag_83 : _GEN_82; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_84 = 7'h54 == idx ? cache_tag_84 : _GEN_83; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_85 = 7'h55 == idx ? cache_tag_85 : _GEN_84; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_86 = 7'h56 == idx ? cache_tag_86 : _GEN_85; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_87 = 7'h57 == idx ? cache_tag_87 : _GEN_86; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_88 = 7'h58 == idx ? cache_tag_88 : _GEN_87; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_89 = 7'h59 == idx ? cache_tag_89 : _GEN_88; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_90 = 7'h5a == idx ? cache_tag_90 : _GEN_89; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_91 = 7'h5b == idx ? cache_tag_91 : _GEN_90; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_92 = 7'h5c == idx ? cache_tag_92 : _GEN_91; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_93 = 7'h5d == idx ? cache_tag_93 : _GEN_92; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_94 = 7'h5e == idx ? cache_tag_94 : _GEN_93; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_95 = 7'h5f == idx ? cache_tag_95 : _GEN_94; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_96 = 7'h60 == idx ? cache_tag_96 : _GEN_95; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_97 = 7'h61 == idx ? cache_tag_97 : _GEN_96; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_98 = 7'h62 == idx ? cache_tag_98 : _GEN_97; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_99 = 7'h63 == idx ? cache_tag_99 : _GEN_98; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_100 = 7'h64 == idx ? cache_tag_100 : _GEN_99; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_101 = 7'h65 == idx ? cache_tag_101 : _GEN_100; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_102 = 7'h66 == idx ? cache_tag_102 : _GEN_101; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_103 = 7'h67 == idx ? cache_tag_103 : _GEN_102; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_104 = 7'h68 == idx ? cache_tag_104 : _GEN_103; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_105 = 7'h69 == idx ? cache_tag_105 : _GEN_104; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_106 = 7'h6a == idx ? cache_tag_106 : _GEN_105; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_107 = 7'h6b == idx ? cache_tag_107 : _GEN_106; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_108 = 7'h6c == idx ? cache_tag_108 : _GEN_107; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_109 = 7'h6d == idx ? cache_tag_109 : _GEN_108; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_110 = 7'h6e == idx ? cache_tag_110 : _GEN_109; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_111 = 7'h6f == idx ? cache_tag_111 : _GEN_110; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_112 = 7'h70 == idx ? cache_tag_112 : _GEN_111; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_113 = 7'h71 == idx ? cache_tag_113 : _GEN_112; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_114 = 7'h72 == idx ? cache_tag_114 : _GEN_113; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_115 = 7'h73 == idx ? cache_tag_115 : _GEN_114; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_116 = 7'h74 == idx ? cache_tag_116 : _GEN_115; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_117 = 7'h75 == idx ? cache_tag_117 : _GEN_116; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_118 = 7'h76 == idx ? cache_tag_118 : _GEN_117; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_119 = 7'h77 == idx ? cache_tag_119 : _GEN_118; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_120 = 7'h78 == idx ? cache_tag_120 : _GEN_119; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_121 = 7'h79 == idx ? cache_tag_121 : _GEN_120; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_122 = 7'h7a == idx ? cache_tag_122 : _GEN_121; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_123 = 7'h7b == idx ? cache_tag_123 : _GEN_122; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_124 = 7'h7c == idx ? cache_tag_124 : _GEN_123; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_125 = 7'h7d == idx ? cache_tag_125 : _GEN_124; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_126 = 7'h7e == idx ? cache_tag_126 : _GEN_125; // @[icache.scala 50:{33,33}]
  wire [41:0] _GEN_127 = 7'h7f == idx ? cache_tag_127 : _GEN_126; // @[icache.scala 50:{33,33}]
  wire  _GEN_129 = 7'h1 == idx ? valid_1_0 : valid_0_0; // @[icache.scala 50:{70,70}]
  wire  _GEN_130 = 7'h2 == idx ? valid_2_0 : _GEN_129; // @[icache.scala 50:{70,70}]
  wire  _GEN_131 = 7'h3 == idx ? valid_3_0 : _GEN_130; // @[icache.scala 50:{70,70}]
  wire  _GEN_132 = 7'h4 == idx ? valid_4_0 : _GEN_131; // @[icache.scala 50:{70,70}]
  wire  _GEN_133 = 7'h5 == idx ? valid_5_0 : _GEN_132; // @[icache.scala 50:{70,70}]
  wire  _GEN_134 = 7'h6 == idx ? valid_6_0 : _GEN_133; // @[icache.scala 50:{70,70}]
  wire  _GEN_135 = 7'h7 == idx ? valid_7_0 : _GEN_134; // @[icache.scala 50:{70,70}]
  wire  _GEN_136 = 7'h8 == idx ? valid_8_0 : _GEN_135; // @[icache.scala 50:{70,70}]
  wire  _GEN_137 = 7'h9 == idx ? valid_9_0 : _GEN_136; // @[icache.scala 50:{70,70}]
  wire  _GEN_138 = 7'ha == idx ? valid_10_0 : _GEN_137; // @[icache.scala 50:{70,70}]
  wire  _GEN_139 = 7'hb == idx ? valid_11_0 : _GEN_138; // @[icache.scala 50:{70,70}]
  wire  _GEN_140 = 7'hc == idx ? valid_12_0 : _GEN_139; // @[icache.scala 50:{70,70}]
  wire  _GEN_141 = 7'hd == idx ? valid_13_0 : _GEN_140; // @[icache.scala 50:{70,70}]
  wire  _GEN_142 = 7'he == idx ? valid_14_0 : _GEN_141; // @[icache.scala 50:{70,70}]
  wire  _GEN_143 = 7'hf == idx ? valid_15_0 : _GEN_142; // @[icache.scala 50:{70,70}]
  wire  _GEN_144 = 7'h10 == idx ? valid_16_0 : _GEN_143; // @[icache.scala 50:{70,70}]
  wire  _GEN_145 = 7'h11 == idx ? valid_17_0 : _GEN_144; // @[icache.scala 50:{70,70}]
  wire  _GEN_146 = 7'h12 == idx ? valid_18_0 : _GEN_145; // @[icache.scala 50:{70,70}]
  wire  _GEN_147 = 7'h13 == idx ? valid_19_0 : _GEN_146; // @[icache.scala 50:{70,70}]
  wire  _GEN_148 = 7'h14 == idx ? valid_20_0 : _GEN_147; // @[icache.scala 50:{70,70}]
  wire  _GEN_149 = 7'h15 == idx ? valid_21_0 : _GEN_148; // @[icache.scala 50:{70,70}]
  wire  _GEN_150 = 7'h16 == idx ? valid_22_0 : _GEN_149; // @[icache.scala 50:{70,70}]
  wire  _GEN_151 = 7'h17 == idx ? valid_23_0 : _GEN_150; // @[icache.scala 50:{70,70}]
  wire  _GEN_152 = 7'h18 == idx ? valid_24_0 : _GEN_151; // @[icache.scala 50:{70,70}]
  wire  _GEN_153 = 7'h19 == idx ? valid_25_0 : _GEN_152; // @[icache.scala 50:{70,70}]
  wire  _GEN_154 = 7'h1a == idx ? valid_26_0 : _GEN_153; // @[icache.scala 50:{70,70}]
  wire  _GEN_155 = 7'h1b == idx ? valid_27_0 : _GEN_154; // @[icache.scala 50:{70,70}]
  wire  _GEN_156 = 7'h1c == idx ? valid_28_0 : _GEN_155; // @[icache.scala 50:{70,70}]
  wire  _GEN_157 = 7'h1d == idx ? valid_29_0 : _GEN_156; // @[icache.scala 50:{70,70}]
  wire  _GEN_158 = 7'h1e == idx ? valid_30_0 : _GEN_157; // @[icache.scala 50:{70,70}]
  wire  _GEN_159 = 7'h1f == idx ? valid_31_0 : _GEN_158; // @[icache.scala 50:{70,70}]
  wire  _GEN_160 = 7'h20 == idx ? valid_32_0 : _GEN_159; // @[icache.scala 50:{70,70}]
  wire  _GEN_161 = 7'h21 == idx ? valid_33_0 : _GEN_160; // @[icache.scala 50:{70,70}]
  wire  _GEN_162 = 7'h22 == idx ? valid_34_0 : _GEN_161; // @[icache.scala 50:{70,70}]
  wire  _GEN_163 = 7'h23 == idx ? valid_35_0 : _GEN_162; // @[icache.scala 50:{70,70}]
  wire  _GEN_164 = 7'h24 == idx ? valid_36_0 : _GEN_163; // @[icache.scala 50:{70,70}]
  wire  _GEN_165 = 7'h25 == idx ? valid_37_0 : _GEN_164; // @[icache.scala 50:{70,70}]
  wire  _GEN_166 = 7'h26 == idx ? valid_38_0 : _GEN_165; // @[icache.scala 50:{70,70}]
  wire  _GEN_167 = 7'h27 == idx ? valid_39_0 : _GEN_166; // @[icache.scala 50:{70,70}]
  wire  _GEN_168 = 7'h28 == idx ? valid_40_0 : _GEN_167; // @[icache.scala 50:{70,70}]
  wire  _GEN_169 = 7'h29 == idx ? valid_41_0 : _GEN_168; // @[icache.scala 50:{70,70}]
  wire  _GEN_170 = 7'h2a == idx ? valid_42_0 : _GEN_169; // @[icache.scala 50:{70,70}]
  wire  _GEN_171 = 7'h2b == idx ? valid_43_0 : _GEN_170; // @[icache.scala 50:{70,70}]
  wire  _GEN_172 = 7'h2c == idx ? valid_44_0 : _GEN_171; // @[icache.scala 50:{70,70}]
  wire  _GEN_173 = 7'h2d == idx ? valid_45_0 : _GEN_172; // @[icache.scala 50:{70,70}]
  wire  _GEN_174 = 7'h2e == idx ? valid_46_0 : _GEN_173; // @[icache.scala 50:{70,70}]
  wire  _GEN_175 = 7'h2f == idx ? valid_47_0 : _GEN_174; // @[icache.scala 50:{70,70}]
  wire  _GEN_176 = 7'h30 == idx ? valid_48_0 : _GEN_175; // @[icache.scala 50:{70,70}]
  wire  _GEN_177 = 7'h31 == idx ? valid_49_0 : _GEN_176; // @[icache.scala 50:{70,70}]
  wire  _GEN_178 = 7'h32 == idx ? valid_50_0 : _GEN_177; // @[icache.scala 50:{70,70}]
  wire  _GEN_179 = 7'h33 == idx ? valid_51_0 : _GEN_178; // @[icache.scala 50:{70,70}]
  wire  _GEN_180 = 7'h34 == idx ? valid_52_0 : _GEN_179; // @[icache.scala 50:{70,70}]
  wire  _GEN_181 = 7'h35 == idx ? valid_53_0 : _GEN_180; // @[icache.scala 50:{70,70}]
  wire  _GEN_182 = 7'h36 == idx ? valid_54_0 : _GEN_181; // @[icache.scala 50:{70,70}]
  wire  _GEN_183 = 7'h37 == idx ? valid_55_0 : _GEN_182; // @[icache.scala 50:{70,70}]
  wire  _GEN_184 = 7'h38 == idx ? valid_56_0 : _GEN_183; // @[icache.scala 50:{70,70}]
  wire  _GEN_185 = 7'h39 == idx ? valid_57_0 : _GEN_184; // @[icache.scala 50:{70,70}]
  wire  _GEN_186 = 7'h3a == idx ? valid_58_0 : _GEN_185; // @[icache.scala 50:{70,70}]
  wire  _GEN_187 = 7'h3b == idx ? valid_59_0 : _GEN_186; // @[icache.scala 50:{70,70}]
  wire  _GEN_188 = 7'h3c == idx ? valid_60_0 : _GEN_187; // @[icache.scala 50:{70,70}]
  wire  _GEN_189 = 7'h3d == idx ? valid_61_0 : _GEN_188; // @[icache.scala 50:{70,70}]
  wire  _GEN_190 = 7'h3e == idx ? valid_62_0 : _GEN_189; // @[icache.scala 50:{70,70}]
  wire  _GEN_191 = 7'h3f == idx ? valid_63_0 : _GEN_190; // @[icache.scala 50:{70,70}]
  wire  _GEN_192 = 7'h40 == idx ? valid_64_0 : _GEN_191; // @[icache.scala 50:{70,70}]
  wire  _GEN_193 = 7'h41 == idx ? valid_65_0 : _GEN_192; // @[icache.scala 50:{70,70}]
  wire  _GEN_194 = 7'h42 == idx ? valid_66_0 : _GEN_193; // @[icache.scala 50:{70,70}]
  wire  _GEN_195 = 7'h43 == idx ? valid_67_0 : _GEN_194; // @[icache.scala 50:{70,70}]
  wire  _GEN_196 = 7'h44 == idx ? valid_68_0 : _GEN_195; // @[icache.scala 50:{70,70}]
  wire  _GEN_197 = 7'h45 == idx ? valid_69_0 : _GEN_196; // @[icache.scala 50:{70,70}]
  wire  _GEN_198 = 7'h46 == idx ? valid_70_0 : _GEN_197; // @[icache.scala 50:{70,70}]
  wire  _GEN_199 = 7'h47 == idx ? valid_71_0 : _GEN_198; // @[icache.scala 50:{70,70}]
  wire  _GEN_200 = 7'h48 == idx ? valid_72_0 : _GEN_199; // @[icache.scala 50:{70,70}]
  wire  _GEN_201 = 7'h49 == idx ? valid_73_0 : _GEN_200; // @[icache.scala 50:{70,70}]
  wire  _GEN_202 = 7'h4a == idx ? valid_74_0 : _GEN_201; // @[icache.scala 50:{70,70}]
  wire  _GEN_203 = 7'h4b == idx ? valid_75_0 : _GEN_202; // @[icache.scala 50:{70,70}]
  wire  _GEN_204 = 7'h4c == idx ? valid_76_0 : _GEN_203; // @[icache.scala 50:{70,70}]
  wire  _GEN_205 = 7'h4d == idx ? valid_77_0 : _GEN_204; // @[icache.scala 50:{70,70}]
  wire  _GEN_206 = 7'h4e == idx ? valid_78_0 : _GEN_205; // @[icache.scala 50:{70,70}]
  wire  _GEN_207 = 7'h4f == idx ? valid_79_0 : _GEN_206; // @[icache.scala 50:{70,70}]
  wire  _GEN_208 = 7'h50 == idx ? valid_80_0 : _GEN_207; // @[icache.scala 50:{70,70}]
  wire  _GEN_209 = 7'h51 == idx ? valid_81_0 : _GEN_208; // @[icache.scala 50:{70,70}]
  wire  _GEN_210 = 7'h52 == idx ? valid_82_0 : _GEN_209; // @[icache.scala 50:{70,70}]
  wire  _GEN_211 = 7'h53 == idx ? valid_83_0 : _GEN_210; // @[icache.scala 50:{70,70}]
  wire  _GEN_212 = 7'h54 == idx ? valid_84_0 : _GEN_211; // @[icache.scala 50:{70,70}]
  wire  _GEN_213 = 7'h55 == idx ? valid_85_0 : _GEN_212; // @[icache.scala 50:{70,70}]
  wire  _GEN_214 = 7'h56 == idx ? valid_86_0 : _GEN_213; // @[icache.scala 50:{70,70}]
  wire  _GEN_215 = 7'h57 == idx ? valid_87_0 : _GEN_214; // @[icache.scala 50:{70,70}]
  wire  _GEN_216 = 7'h58 == idx ? valid_88_0 : _GEN_215; // @[icache.scala 50:{70,70}]
  wire  _GEN_217 = 7'h59 == idx ? valid_89_0 : _GEN_216; // @[icache.scala 50:{70,70}]
  wire  _GEN_218 = 7'h5a == idx ? valid_90_0 : _GEN_217; // @[icache.scala 50:{70,70}]
  wire  _GEN_219 = 7'h5b == idx ? valid_91_0 : _GEN_218; // @[icache.scala 50:{70,70}]
  wire  _GEN_220 = 7'h5c == idx ? valid_92_0 : _GEN_219; // @[icache.scala 50:{70,70}]
  wire  _GEN_221 = 7'h5d == idx ? valid_93_0 : _GEN_220; // @[icache.scala 50:{70,70}]
  wire  _GEN_222 = 7'h5e == idx ? valid_94_0 : _GEN_221; // @[icache.scala 50:{70,70}]
  wire  _GEN_223 = 7'h5f == idx ? valid_95_0 : _GEN_222; // @[icache.scala 50:{70,70}]
  wire  _GEN_224 = 7'h60 == idx ? valid_96_0 : _GEN_223; // @[icache.scala 50:{70,70}]
  wire  _GEN_225 = 7'h61 == idx ? valid_97_0 : _GEN_224; // @[icache.scala 50:{70,70}]
  wire  _GEN_226 = 7'h62 == idx ? valid_98_0 : _GEN_225; // @[icache.scala 50:{70,70}]
  wire  _GEN_227 = 7'h63 == idx ? valid_99_0 : _GEN_226; // @[icache.scala 50:{70,70}]
  wire  _GEN_228 = 7'h64 == idx ? valid_100_0 : _GEN_227; // @[icache.scala 50:{70,70}]
  wire  _GEN_229 = 7'h65 == idx ? valid_101_0 : _GEN_228; // @[icache.scala 50:{70,70}]
  wire  _GEN_230 = 7'h66 == idx ? valid_102_0 : _GEN_229; // @[icache.scala 50:{70,70}]
  wire  _GEN_231 = 7'h67 == idx ? valid_103_0 : _GEN_230; // @[icache.scala 50:{70,70}]
  wire  _GEN_232 = 7'h68 == idx ? valid_104_0 : _GEN_231; // @[icache.scala 50:{70,70}]
  wire  _GEN_233 = 7'h69 == idx ? valid_105_0 : _GEN_232; // @[icache.scala 50:{70,70}]
  wire  _GEN_234 = 7'h6a == idx ? valid_106_0 : _GEN_233; // @[icache.scala 50:{70,70}]
  wire  _GEN_235 = 7'h6b == idx ? valid_107_0 : _GEN_234; // @[icache.scala 50:{70,70}]
  wire  _GEN_236 = 7'h6c == idx ? valid_108_0 : _GEN_235; // @[icache.scala 50:{70,70}]
  wire  _GEN_237 = 7'h6d == idx ? valid_109_0 : _GEN_236; // @[icache.scala 50:{70,70}]
  wire  _GEN_238 = 7'h6e == idx ? valid_110_0 : _GEN_237; // @[icache.scala 50:{70,70}]
  wire  _GEN_239 = 7'h6f == idx ? valid_111_0 : _GEN_238; // @[icache.scala 50:{70,70}]
  wire  _GEN_240 = 7'h70 == idx ? valid_112_0 : _GEN_239; // @[icache.scala 50:{70,70}]
  wire  _GEN_241 = 7'h71 == idx ? valid_113_0 : _GEN_240; // @[icache.scala 50:{70,70}]
  wire  _GEN_242 = 7'h72 == idx ? valid_114_0 : _GEN_241; // @[icache.scala 50:{70,70}]
  wire  _GEN_243 = 7'h73 == idx ? valid_115_0 : _GEN_242; // @[icache.scala 50:{70,70}]
  wire  _GEN_244 = 7'h74 == idx ? valid_116_0 : _GEN_243; // @[icache.scala 50:{70,70}]
  wire  _GEN_245 = 7'h75 == idx ? valid_117_0 : _GEN_244; // @[icache.scala 50:{70,70}]
  wire  _GEN_246 = 7'h76 == idx ? valid_118_0 : _GEN_245; // @[icache.scala 50:{70,70}]
  wire  _GEN_247 = 7'h77 == idx ? valid_119_0 : _GEN_246; // @[icache.scala 50:{70,70}]
  wire  _GEN_248 = 7'h78 == idx ? valid_120_0 : _GEN_247; // @[icache.scala 50:{70,70}]
  wire  _GEN_249 = 7'h79 == idx ? valid_121_0 : _GEN_248; // @[icache.scala 50:{70,70}]
  wire  _GEN_250 = 7'h7a == idx ? valid_122_0 : _GEN_249; // @[icache.scala 50:{70,70}]
  wire  _GEN_251 = 7'h7b == idx ? valid_123_0 : _GEN_250; // @[icache.scala 50:{70,70}]
  wire  _GEN_252 = 7'h7c == idx ? valid_124_0 : _GEN_251; // @[icache.scala 50:{70,70}]
  wire  _GEN_253 = 7'h7d == idx ? valid_125_0 : _GEN_252; // @[icache.scala 50:{70,70}]
  wire  _GEN_254 = 7'h7e == idx ? valid_126_0 : _GEN_253; // @[icache.scala 50:{70,70}]
  wire  _GEN_255 = 7'h7f == idx ? valid_127_0 : _GEN_254; // @[icache.scala 50:{70,70}]
  wire  _GEN_257 = 7'h1 == idx ? valid_1_1 : valid_0_1; // @[icache.scala 51:{70,70}]
  wire  _GEN_258 = 7'h2 == idx ? valid_2_1 : _GEN_257; // @[icache.scala 51:{70,70}]
  wire  _GEN_259 = 7'h3 == idx ? valid_3_1 : _GEN_258; // @[icache.scala 51:{70,70}]
  wire  _GEN_260 = 7'h4 == idx ? valid_4_1 : _GEN_259; // @[icache.scala 51:{70,70}]
  wire  _GEN_261 = 7'h5 == idx ? valid_5_1 : _GEN_260; // @[icache.scala 51:{70,70}]
  wire  _GEN_262 = 7'h6 == idx ? valid_6_1 : _GEN_261; // @[icache.scala 51:{70,70}]
  wire  _GEN_263 = 7'h7 == idx ? valid_7_1 : _GEN_262; // @[icache.scala 51:{70,70}]
  wire  _GEN_264 = 7'h8 == idx ? valid_8_1 : _GEN_263; // @[icache.scala 51:{70,70}]
  wire  _GEN_265 = 7'h9 == idx ? valid_9_1 : _GEN_264; // @[icache.scala 51:{70,70}]
  wire  _GEN_266 = 7'ha == idx ? valid_10_1 : _GEN_265; // @[icache.scala 51:{70,70}]
  wire  _GEN_267 = 7'hb == idx ? valid_11_1 : _GEN_266; // @[icache.scala 51:{70,70}]
  wire  _GEN_268 = 7'hc == idx ? valid_12_1 : _GEN_267; // @[icache.scala 51:{70,70}]
  wire  _GEN_269 = 7'hd == idx ? valid_13_1 : _GEN_268; // @[icache.scala 51:{70,70}]
  wire  _GEN_270 = 7'he == idx ? valid_14_1 : _GEN_269; // @[icache.scala 51:{70,70}]
  wire  _GEN_271 = 7'hf == idx ? valid_15_1 : _GEN_270; // @[icache.scala 51:{70,70}]
  wire  _GEN_272 = 7'h10 == idx ? valid_16_1 : _GEN_271; // @[icache.scala 51:{70,70}]
  wire  _GEN_273 = 7'h11 == idx ? valid_17_1 : _GEN_272; // @[icache.scala 51:{70,70}]
  wire  _GEN_274 = 7'h12 == idx ? valid_18_1 : _GEN_273; // @[icache.scala 51:{70,70}]
  wire  _GEN_275 = 7'h13 == idx ? valid_19_1 : _GEN_274; // @[icache.scala 51:{70,70}]
  wire  _GEN_276 = 7'h14 == idx ? valid_20_1 : _GEN_275; // @[icache.scala 51:{70,70}]
  wire  _GEN_277 = 7'h15 == idx ? valid_21_1 : _GEN_276; // @[icache.scala 51:{70,70}]
  wire  _GEN_278 = 7'h16 == idx ? valid_22_1 : _GEN_277; // @[icache.scala 51:{70,70}]
  wire  _GEN_279 = 7'h17 == idx ? valid_23_1 : _GEN_278; // @[icache.scala 51:{70,70}]
  wire  _GEN_280 = 7'h18 == idx ? valid_24_1 : _GEN_279; // @[icache.scala 51:{70,70}]
  wire  _GEN_281 = 7'h19 == idx ? valid_25_1 : _GEN_280; // @[icache.scala 51:{70,70}]
  wire  _GEN_282 = 7'h1a == idx ? valid_26_1 : _GEN_281; // @[icache.scala 51:{70,70}]
  wire  _GEN_283 = 7'h1b == idx ? valid_27_1 : _GEN_282; // @[icache.scala 51:{70,70}]
  wire  _GEN_284 = 7'h1c == idx ? valid_28_1 : _GEN_283; // @[icache.scala 51:{70,70}]
  wire  _GEN_285 = 7'h1d == idx ? valid_29_1 : _GEN_284; // @[icache.scala 51:{70,70}]
  wire  _GEN_286 = 7'h1e == idx ? valid_30_1 : _GEN_285; // @[icache.scala 51:{70,70}]
  wire  _GEN_287 = 7'h1f == idx ? valid_31_1 : _GEN_286; // @[icache.scala 51:{70,70}]
  wire  _GEN_288 = 7'h20 == idx ? valid_32_1 : _GEN_287; // @[icache.scala 51:{70,70}]
  wire  _GEN_289 = 7'h21 == idx ? valid_33_1 : _GEN_288; // @[icache.scala 51:{70,70}]
  wire  _GEN_290 = 7'h22 == idx ? valid_34_1 : _GEN_289; // @[icache.scala 51:{70,70}]
  wire  _GEN_291 = 7'h23 == idx ? valid_35_1 : _GEN_290; // @[icache.scala 51:{70,70}]
  wire  _GEN_292 = 7'h24 == idx ? valid_36_1 : _GEN_291; // @[icache.scala 51:{70,70}]
  wire  _GEN_293 = 7'h25 == idx ? valid_37_1 : _GEN_292; // @[icache.scala 51:{70,70}]
  wire  _GEN_294 = 7'h26 == idx ? valid_38_1 : _GEN_293; // @[icache.scala 51:{70,70}]
  wire  _GEN_295 = 7'h27 == idx ? valid_39_1 : _GEN_294; // @[icache.scala 51:{70,70}]
  wire  _GEN_296 = 7'h28 == idx ? valid_40_1 : _GEN_295; // @[icache.scala 51:{70,70}]
  wire  _GEN_297 = 7'h29 == idx ? valid_41_1 : _GEN_296; // @[icache.scala 51:{70,70}]
  wire  _GEN_298 = 7'h2a == idx ? valid_42_1 : _GEN_297; // @[icache.scala 51:{70,70}]
  wire  _GEN_299 = 7'h2b == idx ? valid_43_1 : _GEN_298; // @[icache.scala 51:{70,70}]
  wire  _GEN_300 = 7'h2c == idx ? valid_44_1 : _GEN_299; // @[icache.scala 51:{70,70}]
  wire  _GEN_301 = 7'h2d == idx ? valid_45_1 : _GEN_300; // @[icache.scala 51:{70,70}]
  wire  _GEN_302 = 7'h2e == idx ? valid_46_1 : _GEN_301; // @[icache.scala 51:{70,70}]
  wire  _GEN_303 = 7'h2f == idx ? valid_47_1 : _GEN_302; // @[icache.scala 51:{70,70}]
  wire  _GEN_304 = 7'h30 == idx ? valid_48_1 : _GEN_303; // @[icache.scala 51:{70,70}]
  wire  _GEN_305 = 7'h31 == idx ? valid_49_1 : _GEN_304; // @[icache.scala 51:{70,70}]
  wire  _GEN_306 = 7'h32 == idx ? valid_50_1 : _GEN_305; // @[icache.scala 51:{70,70}]
  wire  _GEN_307 = 7'h33 == idx ? valid_51_1 : _GEN_306; // @[icache.scala 51:{70,70}]
  wire  _GEN_308 = 7'h34 == idx ? valid_52_1 : _GEN_307; // @[icache.scala 51:{70,70}]
  wire  _GEN_309 = 7'h35 == idx ? valid_53_1 : _GEN_308; // @[icache.scala 51:{70,70}]
  wire  _GEN_310 = 7'h36 == idx ? valid_54_1 : _GEN_309; // @[icache.scala 51:{70,70}]
  wire  _GEN_311 = 7'h37 == idx ? valid_55_1 : _GEN_310; // @[icache.scala 51:{70,70}]
  wire  _GEN_312 = 7'h38 == idx ? valid_56_1 : _GEN_311; // @[icache.scala 51:{70,70}]
  wire  _GEN_313 = 7'h39 == idx ? valid_57_1 : _GEN_312; // @[icache.scala 51:{70,70}]
  wire  _GEN_314 = 7'h3a == idx ? valid_58_1 : _GEN_313; // @[icache.scala 51:{70,70}]
  wire  _GEN_315 = 7'h3b == idx ? valid_59_1 : _GEN_314; // @[icache.scala 51:{70,70}]
  wire  _GEN_316 = 7'h3c == idx ? valid_60_1 : _GEN_315; // @[icache.scala 51:{70,70}]
  wire  _GEN_317 = 7'h3d == idx ? valid_61_1 : _GEN_316; // @[icache.scala 51:{70,70}]
  wire  _GEN_318 = 7'h3e == idx ? valid_62_1 : _GEN_317; // @[icache.scala 51:{70,70}]
  wire  _GEN_319 = 7'h3f == idx ? valid_63_1 : _GEN_318; // @[icache.scala 51:{70,70}]
  wire  _GEN_320 = 7'h40 == idx ? valid_64_1 : _GEN_319; // @[icache.scala 51:{70,70}]
  wire  _GEN_321 = 7'h41 == idx ? valid_65_1 : _GEN_320; // @[icache.scala 51:{70,70}]
  wire  _GEN_322 = 7'h42 == idx ? valid_66_1 : _GEN_321; // @[icache.scala 51:{70,70}]
  wire  _GEN_323 = 7'h43 == idx ? valid_67_1 : _GEN_322; // @[icache.scala 51:{70,70}]
  wire  _GEN_324 = 7'h44 == idx ? valid_68_1 : _GEN_323; // @[icache.scala 51:{70,70}]
  wire  _GEN_325 = 7'h45 == idx ? valid_69_1 : _GEN_324; // @[icache.scala 51:{70,70}]
  wire  _GEN_326 = 7'h46 == idx ? valid_70_1 : _GEN_325; // @[icache.scala 51:{70,70}]
  wire  _GEN_327 = 7'h47 == idx ? valid_71_1 : _GEN_326; // @[icache.scala 51:{70,70}]
  wire  _GEN_328 = 7'h48 == idx ? valid_72_1 : _GEN_327; // @[icache.scala 51:{70,70}]
  wire  _GEN_329 = 7'h49 == idx ? valid_73_1 : _GEN_328; // @[icache.scala 51:{70,70}]
  wire  _GEN_330 = 7'h4a == idx ? valid_74_1 : _GEN_329; // @[icache.scala 51:{70,70}]
  wire  _GEN_331 = 7'h4b == idx ? valid_75_1 : _GEN_330; // @[icache.scala 51:{70,70}]
  wire  _GEN_332 = 7'h4c == idx ? valid_76_1 : _GEN_331; // @[icache.scala 51:{70,70}]
  wire  _GEN_333 = 7'h4d == idx ? valid_77_1 : _GEN_332; // @[icache.scala 51:{70,70}]
  wire  _GEN_334 = 7'h4e == idx ? valid_78_1 : _GEN_333; // @[icache.scala 51:{70,70}]
  wire  _GEN_335 = 7'h4f == idx ? valid_79_1 : _GEN_334; // @[icache.scala 51:{70,70}]
  wire  _GEN_336 = 7'h50 == idx ? valid_80_1 : _GEN_335; // @[icache.scala 51:{70,70}]
  wire  _GEN_337 = 7'h51 == idx ? valid_81_1 : _GEN_336; // @[icache.scala 51:{70,70}]
  wire  _GEN_338 = 7'h52 == idx ? valid_82_1 : _GEN_337; // @[icache.scala 51:{70,70}]
  wire  _GEN_339 = 7'h53 == idx ? valid_83_1 : _GEN_338; // @[icache.scala 51:{70,70}]
  wire  _GEN_340 = 7'h54 == idx ? valid_84_1 : _GEN_339; // @[icache.scala 51:{70,70}]
  wire  _GEN_341 = 7'h55 == idx ? valid_85_1 : _GEN_340; // @[icache.scala 51:{70,70}]
  wire  _GEN_342 = 7'h56 == idx ? valid_86_1 : _GEN_341; // @[icache.scala 51:{70,70}]
  wire  _GEN_343 = 7'h57 == idx ? valid_87_1 : _GEN_342; // @[icache.scala 51:{70,70}]
  wire  _GEN_344 = 7'h58 == idx ? valid_88_1 : _GEN_343; // @[icache.scala 51:{70,70}]
  wire  _GEN_345 = 7'h59 == idx ? valid_89_1 : _GEN_344; // @[icache.scala 51:{70,70}]
  wire  _GEN_346 = 7'h5a == idx ? valid_90_1 : _GEN_345; // @[icache.scala 51:{70,70}]
  wire  _GEN_347 = 7'h5b == idx ? valid_91_1 : _GEN_346; // @[icache.scala 51:{70,70}]
  wire  _GEN_348 = 7'h5c == idx ? valid_92_1 : _GEN_347; // @[icache.scala 51:{70,70}]
  wire  _GEN_349 = 7'h5d == idx ? valid_93_1 : _GEN_348; // @[icache.scala 51:{70,70}]
  wire  _GEN_350 = 7'h5e == idx ? valid_94_1 : _GEN_349; // @[icache.scala 51:{70,70}]
  wire  _GEN_351 = 7'h5f == idx ? valid_95_1 : _GEN_350; // @[icache.scala 51:{70,70}]
  wire  _GEN_352 = 7'h60 == idx ? valid_96_1 : _GEN_351; // @[icache.scala 51:{70,70}]
  wire  _GEN_353 = 7'h61 == idx ? valid_97_1 : _GEN_352; // @[icache.scala 51:{70,70}]
  wire  _GEN_354 = 7'h62 == idx ? valid_98_1 : _GEN_353; // @[icache.scala 51:{70,70}]
  wire  _GEN_355 = 7'h63 == idx ? valid_99_1 : _GEN_354; // @[icache.scala 51:{70,70}]
  wire  _GEN_356 = 7'h64 == idx ? valid_100_1 : _GEN_355; // @[icache.scala 51:{70,70}]
  wire  _GEN_357 = 7'h65 == idx ? valid_101_1 : _GEN_356; // @[icache.scala 51:{70,70}]
  wire  _GEN_358 = 7'h66 == idx ? valid_102_1 : _GEN_357; // @[icache.scala 51:{70,70}]
  wire  _GEN_359 = 7'h67 == idx ? valid_103_1 : _GEN_358; // @[icache.scala 51:{70,70}]
  wire  _GEN_360 = 7'h68 == idx ? valid_104_1 : _GEN_359; // @[icache.scala 51:{70,70}]
  wire  _GEN_361 = 7'h69 == idx ? valid_105_1 : _GEN_360; // @[icache.scala 51:{70,70}]
  wire  _GEN_362 = 7'h6a == idx ? valid_106_1 : _GEN_361; // @[icache.scala 51:{70,70}]
  wire  _GEN_363 = 7'h6b == idx ? valid_107_1 : _GEN_362; // @[icache.scala 51:{70,70}]
  wire  _GEN_364 = 7'h6c == idx ? valid_108_1 : _GEN_363; // @[icache.scala 51:{70,70}]
  wire  _GEN_365 = 7'h6d == idx ? valid_109_1 : _GEN_364; // @[icache.scala 51:{70,70}]
  wire  _GEN_366 = 7'h6e == idx ? valid_110_1 : _GEN_365; // @[icache.scala 51:{70,70}]
  wire  _GEN_367 = 7'h6f == idx ? valid_111_1 : _GEN_366; // @[icache.scala 51:{70,70}]
  wire  _GEN_368 = 7'h70 == idx ? valid_112_1 : _GEN_367; // @[icache.scala 51:{70,70}]
  wire  _GEN_369 = 7'h71 == idx ? valid_113_1 : _GEN_368; // @[icache.scala 51:{70,70}]
  wire  _GEN_370 = 7'h72 == idx ? valid_114_1 : _GEN_369; // @[icache.scala 51:{70,70}]
  wire  _GEN_371 = 7'h73 == idx ? valid_115_1 : _GEN_370; // @[icache.scala 51:{70,70}]
  wire  _GEN_372 = 7'h74 == idx ? valid_116_1 : _GEN_371; // @[icache.scala 51:{70,70}]
  wire  _GEN_373 = 7'h75 == idx ? valid_117_1 : _GEN_372; // @[icache.scala 51:{70,70}]
  wire  _GEN_374 = 7'h76 == idx ? valid_118_1 : _GEN_373; // @[icache.scala 51:{70,70}]
  wire  _GEN_375 = 7'h77 == idx ? valid_119_1 : _GEN_374; // @[icache.scala 51:{70,70}]
  wire  _GEN_376 = 7'h78 == idx ? valid_120_1 : _GEN_375; // @[icache.scala 51:{70,70}]
  wire  _GEN_377 = 7'h79 == idx ? valid_121_1 : _GEN_376; // @[icache.scala 51:{70,70}]
  wire  _GEN_378 = 7'h7a == idx ? valid_122_1 : _GEN_377; // @[icache.scala 51:{70,70}]
  wire  _GEN_379 = 7'h7b == idx ? valid_123_1 : _GEN_378; // @[icache.scala 51:{70,70}]
  wire  _GEN_380 = 7'h7c == idx ? valid_124_1 : _GEN_379; // @[icache.scala 51:{70,70}]
  wire  _GEN_381 = 7'h7d == idx ? valid_125_1 : _GEN_380; // @[icache.scala 51:{70,70}]
  wire  _GEN_382 = 7'h7e == idx ? valid_126_1 : _GEN_381; // @[icache.scala 51:{70,70}]
  wire  _GEN_383 = 7'h7f == idx ? valid_127_1 : _GEN_382; // @[icache.scala 51:{70,70}]
  wire [1:0] _hit_T_8 = _GEN_127[41:21] == tag & _GEN_383 ? 2'h1 : 2'h3; // @[icache.scala 51:16]
  wire [1:0] hit = _GEN_127[20:0] == tag & _GEN_255 ? 2'h0 : _hit_T_8; // @[icache.scala 50:16]
  wire  hit_way = hit[0]; // @[icache.scala 52:21]
  wire  miss = hit[1] | uncache; // @[icache.scala 53:29]
  wire  _lfsr8_io_en_T = state == 2'h2; // @[icache.scala 55:25]
  reg  way; // @[Reg.scala 35:20]
  reg  cnt; // @[icache.scala 58:20]
  wire [1:0] _state_T_1 = req ? 2'h1 : 2'h0; // @[icache.scala 61:49]
  wire [1:0] _state_T_2 = io_flush ? 2'h0 : _state_T_1; // @[icache.scala 61:22]
  wire [1:0] _state_T_5 = miss ? 2'h2 : _state_T_1; // @[icache.scala 62:49]
  wire [1:0] _state_T_6 = io_flush ? 2'h0 : _state_T_5; // @[icache.scala 62:22]
  wire  _state_T_8 = io_mem_ar_ready & io_mem_ar_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _state_T_9 = _state_T_8 ? 2'h3 : 2'h2; // @[icache.scala 64:49]
  wire  _state_T_12 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 52:35]
  wire  _state_T_14 = _state_T_12 & io_mem_r_bits_last; // @[icache.scala 65:64]
  wire  _valid_T_2 = _lfsr8_io_en_T & ~uncache; // @[icache.scala 68:43]
  wire  _GEN_386 = 7'h0 == idx & way ? valid_0_1 : valid_0_0; // @[icache.scala 68:{25,25}]
  wire  _GEN_1027 = ~way; // @[icache.scala 68:{25,25}]
  wire  _GEN_387 = 7'h1 == idx & ~way ? valid_1_0 : _GEN_386; // @[icache.scala 68:{25,25}]
  wire  _GEN_388 = 7'h1 == idx & way ? valid_1_1 : _GEN_387; // @[icache.scala 68:{25,25}]
  wire  _GEN_389 = 7'h2 == idx & ~way ? valid_2_0 : _GEN_388; // @[icache.scala 68:{25,25}]
  wire  _GEN_390 = 7'h2 == idx & way ? valid_2_1 : _GEN_389; // @[icache.scala 68:{25,25}]
  wire  _GEN_391 = 7'h3 == idx & ~way ? valid_3_0 : _GEN_390; // @[icache.scala 68:{25,25}]
  wire  _GEN_392 = 7'h3 == idx & way ? valid_3_1 : _GEN_391; // @[icache.scala 68:{25,25}]
  wire  _GEN_393 = 7'h4 == idx & ~way ? valid_4_0 : _GEN_392; // @[icache.scala 68:{25,25}]
  wire  _GEN_394 = 7'h4 == idx & way ? valid_4_1 : _GEN_393; // @[icache.scala 68:{25,25}]
  wire  _GEN_395 = 7'h5 == idx & ~way ? valid_5_0 : _GEN_394; // @[icache.scala 68:{25,25}]
  wire  _GEN_396 = 7'h5 == idx & way ? valid_5_1 : _GEN_395; // @[icache.scala 68:{25,25}]
  wire  _GEN_397 = 7'h6 == idx & ~way ? valid_6_0 : _GEN_396; // @[icache.scala 68:{25,25}]
  wire  _GEN_398 = 7'h6 == idx & way ? valid_6_1 : _GEN_397; // @[icache.scala 68:{25,25}]
  wire  _GEN_399 = 7'h7 == idx & ~way ? valid_7_0 : _GEN_398; // @[icache.scala 68:{25,25}]
  wire  _GEN_400 = 7'h7 == idx & way ? valid_7_1 : _GEN_399; // @[icache.scala 68:{25,25}]
  wire  _GEN_401 = 7'h8 == idx & ~way ? valid_8_0 : _GEN_400; // @[icache.scala 68:{25,25}]
  wire  _GEN_402 = 7'h8 == idx & way ? valid_8_1 : _GEN_401; // @[icache.scala 68:{25,25}]
  wire  _GEN_403 = 7'h9 == idx & ~way ? valid_9_0 : _GEN_402; // @[icache.scala 68:{25,25}]
  wire  _GEN_404 = 7'h9 == idx & way ? valid_9_1 : _GEN_403; // @[icache.scala 68:{25,25}]
  wire  _GEN_405 = 7'ha == idx & ~way ? valid_10_0 : _GEN_404; // @[icache.scala 68:{25,25}]
  wire  _GEN_406 = 7'ha == idx & way ? valid_10_1 : _GEN_405; // @[icache.scala 68:{25,25}]
  wire  _GEN_407 = 7'hb == idx & ~way ? valid_11_0 : _GEN_406; // @[icache.scala 68:{25,25}]
  wire  _GEN_408 = 7'hb == idx & way ? valid_11_1 : _GEN_407; // @[icache.scala 68:{25,25}]
  wire  _GEN_409 = 7'hc == idx & ~way ? valid_12_0 : _GEN_408; // @[icache.scala 68:{25,25}]
  wire  _GEN_410 = 7'hc == idx & way ? valid_12_1 : _GEN_409; // @[icache.scala 68:{25,25}]
  wire  _GEN_411 = 7'hd == idx & ~way ? valid_13_0 : _GEN_410; // @[icache.scala 68:{25,25}]
  wire  _GEN_412 = 7'hd == idx & way ? valid_13_1 : _GEN_411; // @[icache.scala 68:{25,25}]
  wire  _GEN_413 = 7'he == idx & ~way ? valid_14_0 : _GEN_412; // @[icache.scala 68:{25,25}]
  wire  _GEN_414 = 7'he == idx & way ? valid_14_1 : _GEN_413; // @[icache.scala 68:{25,25}]
  wire  _GEN_415 = 7'hf == idx & ~way ? valid_15_0 : _GEN_414; // @[icache.scala 68:{25,25}]
  wire  _GEN_416 = 7'hf == idx & way ? valid_15_1 : _GEN_415; // @[icache.scala 68:{25,25}]
  wire  _GEN_417 = 7'h10 == idx & ~way ? valid_16_0 : _GEN_416; // @[icache.scala 68:{25,25}]
  wire  _GEN_418 = 7'h10 == idx & way ? valid_16_1 : _GEN_417; // @[icache.scala 68:{25,25}]
  wire  _GEN_419 = 7'h11 == idx & ~way ? valid_17_0 : _GEN_418; // @[icache.scala 68:{25,25}]
  wire  _GEN_420 = 7'h11 == idx & way ? valid_17_1 : _GEN_419; // @[icache.scala 68:{25,25}]
  wire  _GEN_421 = 7'h12 == idx & ~way ? valid_18_0 : _GEN_420; // @[icache.scala 68:{25,25}]
  wire  _GEN_422 = 7'h12 == idx & way ? valid_18_1 : _GEN_421; // @[icache.scala 68:{25,25}]
  wire  _GEN_423 = 7'h13 == idx & ~way ? valid_19_0 : _GEN_422; // @[icache.scala 68:{25,25}]
  wire  _GEN_424 = 7'h13 == idx & way ? valid_19_1 : _GEN_423; // @[icache.scala 68:{25,25}]
  wire  _GEN_425 = 7'h14 == idx & ~way ? valid_20_0 : _GEN_424; // @[icache.scala 68:{25,25}]
  wire  _GEN_426 = 7'h14 == idx & way ? valid_20_1 : _GEN_425; // @[icache.scala 68:{25,25}]
  wire  _GEN_427 = 7'h15 == idx & ~way ? valid_21_0 : _GEN_426; // @[icache.scala 68:{25,25}]
  wire  _GEN_428 = 7'h15 == idx & way ? valid_21_1 : _GEN_427; // @[icache.scala 68:{25,25}]
  wire  _GEN_429 = 7'h16 == idx & ~way ? valid_22_0 : _GEN_428; // @[icache.scala 68:{25,25}]
  wire  _GEN_430 = 7'h16 == idx & way ? valid_22_1 : _GEN_429; // @[icache.scala 68:{25,25}]
  wire  _GEN_431 = 7'h17 == idx & ~way ? valid_23_0 : _GEN_430; // @[icache.scala 68:{25,25}]
  wire  _GEN_432 = 7'h17 == idx & way ? valid_23_1 : _GEN_431; // @[icache.scala 68:{25,25}]
  wire  _GEN_433 = 7'h18 == idx & ~way ? valid_24_0 : _GEN_432; // @[icache.scala 68:{25,25}]
  wire  _GEN_434 = 7'h18 == idx & way ? valid_24_1 : _GEN_433; // @[icache.scala 68:{25,25}]
  wire  _GEN_435 = 7'h19 == idx & ~way ? valid_25_0 : _GEN_434; // @[icache.scala 68:{25,25}]
  wire  _GEN_436 = 7'h19 == idx & way ? valid_25_1 : _GEN_435; // @[icache.scala 68:{25,25}]
  wire  _GEN_437 = 7'h1a == idx & ~way ? valid_26_0 : _GEN_436; // @[icache.scala 68:{25,25}]
  wire  _GEN_438 = 7'h1a == idx & way ? valid_26_1 : _GEN_437; // @[icache.scala 68:{25,25}]
  wire  _GEN_439 = 7'h1b == idx & ~way ? valid_27_0 : _GEN_438; // @[icache.scala 68:{25,25}]
  wire  _GEN_440 = 7'h1b == idx & way ? valid_27_1 : _GEN_439; // @[icache.scala 68:{25,25}]
  wire  _GEN_441 = 7'h1c == idx & ~way ? valid_28_0 : _GEN_440; // @[icache.scala 68:{25,25}]
  wire  _GEN_442 = 7'h1c == idx & way ? valid_28_1 : _GEN_441; // @[icache.scala 68:{25,25}]
  wire  _GEN_443 = 7'h1d == idx & ~way ? valid_29_0 : _GEN_442; // @[icache.scala 68:{25,25}]
  wire  _GEN_444 = 7'h1d == idx & way ? valid_29_1 : _GEN_443; // @[icache.scala 68:{25,25}]
  wire  _GEN_445 = 7'h1e == idx & ~way ? valid_30_0 : _GEN_444; // @[icache.scala 68:{25,25}]
  wire  _GEN_446 = 7'h1e == idx & way ? valid_30_1 : _GEN_445; // @[icache.scala 68:{25,25}]
  wire  _GEN_447 = 7'h1f == idx & ~way ? valid_31_0 : _GEN_446; // @[icache.scala 68:{25,25}]
  wire  _GEN_448 = 7'h1f == idx & way ? valid_31_1 : _GEN_447; // @[icache.scala 68:{25,25}]
  wire  _GEN_449 = 7'h20 == idx & ~way ? valid_32_0 : _GEN_448; // @[icache.scala 68:{25,25}]
  wire  _GEN_450 = 7'h20 == idx & way ? valid_32_1 : _GEN_449; // @[icache.scala 68:{25,25}]
  wire  _GEN_451 = 7'h21 == idx & ~way ? valid_33_0 : _GEN_450; // @[icache.scala 68:{25,25}]
  wire  _GEN_452 = 7'h21 == idx & way ? valid_33_1 : _GEN_451; // @[icache.scala 68:{25,25}]
  wire  _GEN_453 = 7'h22 == idx & ~way ? valid_34_0 : _GEN_452; // @[icache.scala 68:{25,25}]
  wire  _GEN_454 = 7'h22 == idx & way ? valid_34_1 : _GEN_453; // @[icache.scala 68:{25,25}]
  wire  _GEN_455 = 7'h23 == idx & ~way ? valid_35_0 : _GEN_454; // @[icache.scala 68:{25,25}]
  wire  _GEN_456 = 7'h23 == idx & way ? valid_35_1 : _GEN_455; // @[icache.scala 68:{25,25}]
  wire  _GEN_457 = 7'h24 == idx & ~way ? valid_36_0 : _GEN_456; // @[icache.scala 68:{25,25}]
  wire  _GEN_458 = 7'h24 == idx & way ? valid_36_1 : _GEN_457; // @[icache.scala 68:{25,25}]
  wire  _GEN_459 = 7'h25 == idx & ~way ? valid_37_0 : _GEN_458; // @[icache.scala 68:{25,25}]
  wire  _GEN_460 = 7'h25 == idx & way ? valid_37_1 : _GEN_459; // @[icache.scala 68:{25,25}]
  wire  _GEN_461 = 7'h26 == idx & ~way ? valid_38_0 : _GEN_460; // @[icache.scala 68:{25,25}]
  wire  _GEN_462 = 7'h26 == idx & way ? valid_38_1 : _GEN_461; // @[icache.scala 68:{25,25}]
  wire  _GEN_463 = 7'h27 == idx & ~way ? valid_39_0 : _GEN_462; // @[icache.scala 68:{25,25}]
  wire  _GEN_464 = 7'h27 == idx & way ? valid_39_1 : _GEN_463; // @[icache.scala 68:{25,25}]
  wire  _GEN_465 = 7'h28 == idx & ~way ? valid_40_0 : _GEN_464; // @[icache.scala 68:{25,25}]
  wire  _GEN_466 = 7'h28 == idx & way ? valid_40_1 : _GEN_465; // @[icache.scala 68:{25,25}]
  wire  _GEN_467 = 7'h29 == idx & ~way ? valid_41_0 : _GEN_466; // @[icache.scala 68:{25,25}]
  wire  _GEN_468 = 7'h29 == idx & way ? valid_41_1 : _GEN_467; // @[icache.scala 68:{25,25}]
  wire  _GEN_469 = 7'h2a == idx & ~way ? valid_42_0 : _GEN_468; // @[icache.scala 68:{25,25}]
  wire  _GEN_470 = 7'h2a == idx & way ? valid_42_1 : _GEN_469; // @[icache.scala 68:{25,25}]
  wire  _GEN_471 = 7'h2b == idx & ~way ? valid_43_0 : _GEN_470; // @[icache.scala 68:{25,25}]
  wire  _GEN_472 = 7'h2b == idx & way ? valid_43_1 : _GEN_471; // @[icache.scala 68:{25,25}]
  wire  _GEN_473 = 7'h2c == idx & ~way ? valid_44_0 : _GEN_472; // @[icache.scala 68:{25,25}]
  wire  _GEN_474 = 7'h2c == idx & way ? valid_44_1 : _GEN_473; // @[icache.scala 68:{25,25}]
  wire  _GEN_475 = 7'h2d == idx & ~way ? valid_45_0 : _GEN_474; // @[icache.scala 68:{25,25}]
  wire  _GEN_476 = 7'h2d == idx & way ? valid_45_1 : _GEN_475; // @[icache.scala 68:{25,25}]
  wire  _GEN_477 = 7'h2e == idx & ~way ? valid_46_0 : _GEN_476; // @[icache.scala 68:{25,25}]
  wire  _GEN_478 = 7'h2e == idx & way ? valid_46_1 : _GEN_477; // @[icache.scala 68:{25,25}]
  wire  _GEN_479 = 7'h2f == idx & ~way ? valid_47_0 : _GEN_478; // @[icache.scala 68:{25,25}]
  wire  _GEN_480 = 7'h2f == idx & way ? valid_47_1 : _GEN_479; // @[icache.scala 68:{25,25}]
  wire  _GEN_481 = 7'h30 == idx & ~way ? valid_48_0 : _GEN_480; // @[icache.scala 68:{25,25}]
  wire  _GEN_482 = 7'h30 == idx & way ? valid_48_1 : _GEN_481; // @[icache.scala 68:{25,25}]
  wire  _GEN_483 = 7'h31 == idx & ~way ? valid_49_0 : _GEN_482; // @[icache.scala 68:{25,25}]
  wire  _GEN_484 = 7'h31 == idx & way ? valid_49_1 : _GEN_483; // @[icache.scala 68:{25,25}]
  wire  _GEN_485 = 7'h32 == idx & ~way ? valid_50_0 : _GEN_484; // @[icache.scala 68:{25,25}]
  wire  _GEN_486 = 7'h32 == idx & way ? valid_50_1 : _GEN_485; // @[icache.scala 68:{25,25}]
  wire  _GEN_487 = 7'h33 == idx & ~way ? valid_51_0 : _GEN_486; // @[icache.scala 68:{25,25}]
  wire  _GEN_488 = 7'h33 == idx & way ? valid_51_1 : _GEN_487; // @[icache.scala 68:{25,25}]
  wire  _GEN_489 = 7'h34 == idx & ~way ? valid_52_0 : _GEN_488; // @[icache.scala 68:{25,25}]
  wire  _GEN_490 = 7'h34 == idx & way ? valid_52_1 : _GEN_489; // @[icache.scala 68:{25,25}]
  wire  _GEN_491 = 7'h35 == idx & ~way ? valid_53_0 : _GEN_490; // @[icache.scala 68:{25,25}]
  wire  _GEN_492 = 7'h35 == idx & way ? valid_53_1 : _GEN_491; // @[icache.scala 68:{25,25}]
  wire  _GEN_493 = 7'h36 == idx & ~way ? valid_54_0 : _GEN_492; // @[icache.scala 68:{25,25}]
  wire  _GEN_494 = 7'h36 == idx & way ? valid_54_1 : _GEN_493; // @[icache.scala 68:{25,25}]
  wire  _GEN_495 = 7'h37 == idx & ~way ? valid_55_0 : _GEN_494; // @[icache.scala 68:{25,25}]
  wire  _GEN_496 = 7'h37 == idx & way ? valid_55_1 : _GEN_495; // @[icache.scala 68:{25,25}]
  wire  _GEN_497 = 7'h38 == idx & ~way ? valid_56_0 : _GEN_496; // @[icache.scala 68:{25,25}]
  wire  _GEN_498 = 7'h38 == idx & way ? valid_56_1 : _GEN_497; // @[icache.scala 68:{25,25}]
  wire  _GEN_499 = 7'h39 == idx & ~way ? valid_57_0 : _GEN_498; // @[icache.scala 68:{25,25}]
  wire  _GEN_500 = 7'h39 == idx & way ? valid_57_1 : _GEN_499; // @[icache.scala 68:{25,25}]
  wire  _GEN_501 = 7'h3a == idx & ~way ? valid_58_0 : _GEN_500; // @[icache.scala 68:{25,25}]
  wire  _GEN_502 = 7'h3a == idx & way ? valid_58_1 : _GEN_501; // @[icache.scala 68:{25,25}]
  wire  _GEN_503 = 7'h3b == idx & ~way ? valid_59_0 : _GEN_502; // @[icache.scala 68:{25,25}]
  wire  _GEN_504 = 7'h3b == idx & way ? valid_59_1 : _GEN_503; // @[icache.scala 68:{25,25}]
  wire  _GEN_505 = 7'h3c == idx & ~way ? valid_60_0 : _GEN_504; // @[icache.scala 68:{25,25}]
  wire  _GEN_506 = 7'h3c == idx & way ? valid_60_1 : _GEN_505; // @[icache.scala 68:{25,25}]
  wire  _GEN_507 = 7'h3d == idx & ~way ? valid_61_0 : _GEN_506; // @[icache.scala 68:{25,25}]
  wire  _GEN_508 = 7'h3d == idx & way ? valid_61_1 : _GEN_507; // @[icache.scala 68:{25,25}]
  wire  _GEN_509 = 7'h3e == idx & ~way ? valid_62_0 : _GEN_508; // @[icache.scala 68:{25,25}]
  wire  _GEN_510 = 7'h3e == idx & way ? valid_62_1 : _GEN_509; // @[icache.scala 68:{25,25}]
  wire  _GEN_511 = 7'h3f == idx & ~way ? valid_63_0 : _GEN_510; // @[icache.scala 68:{25,25}]
  wire  _GEN_512 = 7'h3f == idx & way ? valid_63_1 : _GEN_511; // @[icache.scala 68:{25,25}]
  wire  _GEN_513 = 7'h40 == idx & ~way ? valid_64_0 : _GEN_512; // @[icache.scala 68:{25,25}]
  wire  _GEN_514 = 7'h40 == idx & way ? valid_64_1 : _GEN_513; // @[icache.scala 68:{25,25}]
  wire  _GEN_515 = 7'h41 == idx & ~way ? valid_65_0 : _GEN_514; // @[icache.scala 68:{25,25}]
  wire  _GEN_516 = 7'h41 == idx & way ? valid_65_1 : _GEN_515; // @[icache.scala 68:{25,25}]
  wire  _GEN_517 = 7'h42 == idx & ~way ? valid_66_0 : _GEN_516; // @[icache.scala 68:{25,25}]
  wire  _GEN_518 = 7'h42 == idx & way ? valid_66_1 : _GEN_517; // @[icache.scala 68:{25,25}]
  wire  _GEN_519 = 7'h43 == idx & ~way ? valid_67_0 : _GEN_518; // @[icache.scala 68:{25,25}]
  wire  _GEN_520 = 7'h43 == idx & way ? valid_67_1 : _GEN_519; // @[icache.scala 68:{25,25}]
  wire  _GEN_521 = 7'h44 == idx & ~way ? valid_68_0 : _GEN_520; // @[icache.scala 68:{25,25}]
  wire  _GEN_522 = 7'h44 == idx & way ? valid_68_1 : _GEN_521; // @[icache.scala 68:{25,25}]
  wire  _GEN_523 = 7'h45 == idx & ~way ? valid_69_0 : _GEN_522; // @[icache.scala 68:{25,25}]
  wire  _GEN_524 = 7'h45 == idx & way ? valid_69_1 : _GEN_523; // @[icache.scala 68:{25,25}]
  wire  _GEN_525 = 7'h46 == idx & ~way ? valid_70_0 : _GEN_524; // @[icache.scala 68:{25,25}]
  wire  _GEN_526 = 7'h46 == idx & way ? valid_70_1 : _GEN_525; // @[icache.scala 68:{25,25}]
  wire  _GEN_527 = 7'h47 == idx & ~way ? valid_71_0 : _GEN_526; // @[icache.scala 68:{25,25}]
  wire  _GEN_528 = 7'h47 == idx & way ? valid_71_1 : _GEN_527; // @[icache.scala 68:{25,25}]
  wire  _GEN_529 = 7'h48 == idx & ~way ? valid_72_0 : _GEN_528; // @[icache.scala 68:{25,25}]
  wire  _GEN_530 = 7'h48 == idx & way ? valid_72_1 : _GEN_529; // @[icache.scala 68:{25,25}]
  wire  _GEN_531 = 7'h49 == idx & ~way ? valid_73_0 : _GEN_530; // @[icache.scala 68:{25,25}]
  wire  _GEN_532 = 7'h49 == idx & way ? valid_73_1 : _GEN_531; // @[icache.scala 68:{25,25}]
  wire  _GEN_533 = 7'h4a == idx & ~way ? valid_74_0 : _GEN_532; // @[icache.scala 68:{25,25}]
  wire  _GEN_534 = 7'h4a == idx & way ? valid_74_1 : _GEN_533; // @[icache.scala 68:{25,25}]
  wire  _GEN_535 = 7'h4b == idx & ~way ? valid_75_0 : _GEN_534; // @[icache.scala 68:{25,25}]
  wire  _GEN_536 = 7'h4b == idx & way ? valid_75_1 : _GEN_535; // @[icache.scala 68:{25,25}]
  wire  _GEN_537 = 7'h4c == idx & ~way ? valid_76_0 : _GEN_536; // @[icache.scala 68:{25,25}]
  wire  _GEN_538 = 7'h4c == idx & way ? valid_76_1 : _GEN_537; // @[icache.scala 68:{25,25}]
  wire  _GEN_539 = 7'h4d == idx & ~way ? valid_77_0 : _GEN_538; // @[icache.scala 68:{25,25}]
  wire  _GEN_540 = 7'h4d == idx & way ? valid_77_1 : _GEN_539; // @[icache.scala 68:{25,25}]
  wire  _GEN_541 = 7'h4e == idx & ~way ? valid_78_0 : _GEN_540; // @[icache.scala 68:{25,25}]
  wire  _GEN_542 = 7'h4e == idx & way ? valid_78_1 : _GEN_541; // @[icache.scala 68:{25,25}]
  wire  _GEN_543 = 7'h4f == idx & ~way ? valid_79_0 : _GEN_542; // @[icache.scala 68:{25,25}]
  wire  _GEN_544 = 7'h4f == idx & way ? valid_79_1 : _GEN_543; // @[icache.scala 68:{25,25}]
  wire  _GEN_545 = 7'h50 == idx & ~way ? valid_80_0 : _GEN_544; // @[icache.scala 68:{25,25}]
  wire  _GEN_546 = 7'h50 == idx & way ? valid_80_1 : _GEN_545; // @[icache.scala 68:{25,25}]
  wire  _GEN_547 = 7'h51 == idx & ~way ? valid_81_0 : _GEN_546; // @[icache.scala 68:{25,25}]
  wire  _GEN_548 = 7'h51 == idx & way ? valid_81_1 : _GEN_547; // @[icache.scala 68:{25,25}]
  wire  _GEN_549 = 7'h52 == idx & ~way ? valid_82_0 : _GEN_548; // @[icache.scala 68:{25,25}]
  wire  _GEN_550 = 7'h52 == idx & way ? valid_82_1 : _GEN_549; // @[icache.scala 68:{25,25}]
  wire  _GEN_551 = 7'h53 == idx & ~way ? valid_83_0 : _GEN_550; // @[icache.scala 68:{25,25}]
  wire  _GEN_552 = 7'h53 == idx & way ? valid_83_1 : _GEN_551; // @[icache.scala 68:{25,25}]
  wire  _GEN_553 = 7'h54 == idx & ~way ? valid_84_0 : _GEN_552; // @[icache.scala 68:{25,25}]
  wire  _GEN_554 = 7'h54 == idx & way ? valid_84_1 : _GEN_553; // @[icache.scala 68:{25,25}]
  wire  _GEN_555 = 7'h55 == idx & ~way ? valid_85_0 : _GEN_554; // @[icache.scala 68:{25,25}]
  wire  _GEN_556 = 7'h55 == idx & way ? valid_85_1 : _GEN_555; // @[icache.scala 68:{25,25}]
  wire  _GEN_557 = 7'h56 == idx & ~way ? valid_86_0 : _GEN_556; // @[icache.scala 68:{25,25}]
  wire  _GEN_558 = 7'h56 == idx & way ? valid_86_1 : _GEN_557; // @[icache.scala 68:{25,25}]
  wire  _GEN_559 = 7'h57 == idx & ~way ? valid_87_0 : _GEN_558; // @[icache.scala 68:{25,25}]
  wire  _GEN_560 = 7'h57 == idx & way ? valid_87_1 : _GEN_559; // @[icache.scala 68:{25,25}]
  wire  _GEN_561 = 7'h58 == idx & ~way ? valid_88_0 : _GEN_560; // @[icache.scala 68:{25,25}]
  wire  _GEN_562 = 7'h58 == idx & way ? valid_88_1 : _GEN_561; // @[icache.scala 68:{25,25}]
  wire  _GEN_563 = 7'h59 == idx & ~way ? valid_89_0 : _GEN_562; // @[icache.scala 68:{25,25}]
  wire  _GEN_564 = 7'h59 == idx & way ? valid_89_1 : _GEN_563; // @[icache.scala 68:{25,25}]
  wire  _GEN_565 = 7'h5a == idx & ~way ? valid_90_0 : _GEN_564; // @[icache.scala 68:{25,25}]
  wire  _GEN_566 = 7'h5a == idx & way ? valid_90_1 : _GEN_565; // @[icache.scala 68:{25,25}]
  wire  _GEN_567 = 7'h5b == idx & ~way ? valid_91_0 : _GEN_566; // @[icache.scala 68:{25,25}]
  wire  _GEN_568 = 7'h5b == idx & way ? valid_91_1 : _GEN_567; // @[icache.scala 68:{25,25}]
  wire  _GEN_569 = 7'h5c == idx & ~way ? valid_92_0 : _GEN_568; // @[icache.scala 68:{25,25}]
  wire  _GEN_570 = 7'h5c == idx & way ? valid_92_1 : _GEN_569; // @[icache.scala 68:{25,25}]
  wire  _GEN_571 = 7'h5d == idx & ~way ? valid_93_0 : _GEN_570; // @[icache.scala 68:{25,25}]
  wire  _GEN_572 = 7'h5d == idx & way ? valid_93_1 : _GEN_571; // @[icache.scala 68:{25,25}]
  wire  _GEN_573 = 7'h5e == idx & ~way ? valid_94_0 : _GEN_572; // @[icache.scala 68:{25,25}]
  wire  _GEN_574 = 7'h5e == idx & way ? valid_94_1 : _GEN_573; // @[icache.scala 68:{25,25}]
  wire  _GEN_575 = 7'h5f == idx & ~way ? valid_95_0 : _GEN_574; // @[icache.scala 68:{25,25}]
  wire  _GEN_576 = 7'h5f == idx & way ? valid_95_1 : _GEN_575; // @[icache.scala 68:{25,25}]
  wire  _GEN_577 = 7'h60 == idx & ~way ? valid_96_0 : _GEN_576; // @[icache.scala 68:{25,25}]
  wire  _GEN_578 = 7'h60 == idx & way ? valid_96_1 : _GEN_577; // @[icache.scala 68:{25,25}]
  wire  _GEN_579 = 7'h61 == idx & ~way ? valid_97_0 : _GEN_578; // @[icache.scala 68:{25,25}]
  wire  _GEN_580 = 7'h61 == idx & way ? valid_97_1 : _GEN_579; // @[icache.scala 68:{25,25}]
  wire  _GEN_581 = 7'h62 == idx & ~way ? valid_98_0 : _GEN_580; // @[icache.scala 68:{25,25}]
  wire  _GEN_582 = 7'h62 == idx & way ? valid_98_1 : _GEN_581; // @[icache.scala 68:{25,25}]
  wire  _GEN_583 = 7'h63 == idx & ~way ? valid_99_0 : _GEN_582; // @[icache.scala 68:{25,25}]
  wire  _GEN_584 = 7'h63 == idx & way ? valid_99_1 : _GEN_583; // @[icache.scala 68:{25,25}]
  wire  _GEN_585 = 7'h64 == idx & ~way ? valid_100_0 : _GEN_584; // @[icache.scala 68:{25,25}]
  wire  _GEN_586 = 7'h64 == idx & way ? valid_100_1 : _GEN_585; // @[icache.scala 68:{25,25}]
  wire  _GEN_587 = 7'h65 == idx & ~way ? valid_101_0 : _GEN_586; // @[icache.scala 68:{25,25}]
  wire  _GEN_588 = 7'h65 == idx & way ? valid_101_1 : _GEN_587; // @[icache.scala 68:{25,25}]
  wire  _GEN_589 = 7'h66 == idx & ~way ? valid_102_0 : _GEN_588; // @[icache.scala 68:{25,25}]
  wire  _GEN_590 = 7'h66 == idx & way ? valid_102_1 : _GEN_589; // @[icache.scala 68:{25,25}]
  wire  _GEN_591 = 7'h67 == idx & ~way ? valid_103_0 : _GEN_590; // @[icache.scala 68:{25,25}]
  wire  _GEN_592 = 7'h67 == idx & way ? valid_103_1 : _GEN_591; // @[icache.scala 68:{25,25}]
  wire  _GEN_593 = 7'h68 == idx & ~way ? valid_104_0 : _GEN_592; // @[icache.scala 68:{25,25}]
  wire  _GEN_594 = 7'h68 == idx & way ? valid_104_1 : _GEN_593; // @[icache.scala 68:{25,25}]
  wire  _GEN_595 = 7'h69 == idx & ~way ? valid_105_0 : _GEN_594; // @[icache.scala 68:{25,25}]
  wire  _GEN_596 = 7'h69 == idx & way ? valid_105_1 : _GEN_595; // @[icache.scala 68:{25,25}]
  wire  _GEN_597 = 7'h6a == idx & ~way ? valid_106_0 : _GEN_596; // @[icache.scala 68:{25,25}]
  wire  _GEN_598 = 7'h6a == idx & way ? valid_106_1 : _GEN_597; // @[icache.scala 68:{25,25}]
  wire  _GEN_599 = 7'h6b == idx & ~way ? valid_107_0 : _GEN_598; // @[icache.scala 68:{25,25}]
  wire  _GEN_600 = 7'h6b == idx & way ? valid_107_1 : _GEN_599; // @[icache.scala 68:{25,25}]
  wire  _GEN_601 = 7'h6c == idx & ~way ? valid_108_0 : _GEN_600; // @[icache.scala 68:{25,25}]
  wire  _GEN_602 = 7'h6c == idx & way ? valid_108_1 : _GEN_601; // @[icache.scala 68:{25,25}]
  wire  _GEN_603 = 7'h6d == idx & ~way ? valid_109_0 : _GEN_602; // @[icache.scala 68:{25,25}]
  wire  _GEN_604 = 7'h6d == idx & way ? valid_109_1 : _GEN_603; // @[icache.scala 68:{25,25}]
  wire  _GEN_605 = 7'h6e == idx & ~way ? valid_110_0 : _GEN_604; // @[icache.scala 68:{25,25}]
  wire  _GEN_606 = 7'h6e == idx & way ? valid_110_1 : _GEN_605; // @[icache.scala 68:{25,25}]
  wire  _GEN_607 = 7'h6f == idx & ~way ? valid_111_0 : _GEN_606; // @[icache.scala 68:{25,25}]
  wire  _GEN_608 = 7'h6f == idx & way ? valid_111_1 : _GEN_607; // @[icache.scala 68:{25,25}]
  wire  _GEN_609 = 7'h70 == idx & ~way ? valid_112_0 : _GEN_608; // @[icache.scala 68:{25,25}]
  wire  _GEN_610 = 7'h70 == idx & way ? valid_112_1 : _GEN_609; // @[icache.scala 68:{25,25}]
  wire  _GEN_611 = 7'h71 == idx & ~way ? valid_113_0 : _GEN_610; // @[icache.scala 68:{25,25}]
  wire  _GEN_612 = 7'h71 == idx & way ? valid_113_1 : _GEN_611; // @[icache.scala 68:{25,25}]
  wire  _GEN_613 = 7'h72 == idx & ~way ? valid_114_0 : _GEN_612; // @[icache.scala 68:{25,25}]
  wire  _GEN_614 = 7'h72 == idx & way ? valid_114_1 : _GEN_613; // @[icache.scala 68:{25,25}]
  wire  _GEN_615 = 7'h73 == idx & ~way ? valid_115_0 : _GEN_614; // @[icache.scala 68:{25,25}]
  wire  _GEN_616 = 7'h73 == idx & way ? valid_115_1 : _GEN_615; // @[icache.scala 68:{25,25}]
  wire  _GEN_617 = 7'h74 == idx & ~way ? valid_116_0 : _GEN_616; // @[icache.scala 68:{25,25}]
  wire  _GEN_618 = 7'h74 == idx & way ? valid_116_1 : _GEN_617; // @[icache.scala 68:{25,25}]
  wire  _GEN_619 = 7'h75 == idx & ~way ? valid_117_0 : _GEN_618; // @[icache.scala 68:{25,25}]
  wire  _GEN_620 = 7'h75 == idx & way ? valid_117_1 : _GEN_619; // @[icache.scala 68:{25,25}]
  wire  _GEN_621 = 7'h76 == idx & ~way ? valid_118_0 : _GEN_620; // @[icache.scala 68:{25,25}]
  wire  _GEN_622 = 7'h76 == idx & way ? valid_118_1 : _GEN_621; // @[icache.scala 68:{25,25}]
  wire  _GEN_623 = 7'h77 == idx & ~way ? valid_119_0 : _GEN_622; // @[icache.scala 68:{25,25}]
  wire  _GEN_624 = 7'h77 == idx & way ? valid_119_1 : _GEN_623; // @[icache.scala 68:{25,25}]
  wire  _GEN_625 = 7'h78 == idx & ~way ? valid_120_0 : _GEN_624; // @[icache.scala 68:{25,25}]
  wire  _GEN_626 = 7'h78 == idx & way ? valid_120_1 : _GEN_625; // @[icache.scala 68:{25,25}]
  wire  _GEN_627 = 7'h79 == idx & ~way ? valid_121_0 : _GEN_626; // @[icache.scala 68:{25,25}]
  wire  _GEN_628 = 7'h79 == idx & way ? valid_121_1 : _GEN_627; // @[icache.scala 68:{25,25}]
  wire  _GEN_629 = 7'h7a == idx & ~way ? valid_122_0 : _GEN_628; // @[icache.scala 68:{25,25}]
  wire  _GEN_630 = 7'h7a == idx & way ? valid_122_1 : _GEN_629; // @[icache.scala 68:{25,25}]
  wire  _GEN_631 = 7'h7b == idx & ~way ? valid_123_0 : _GEN_630; // @[icache.scala 68:{25,25}]
  wire  _GEN_632 = 7'h7b == idx & way ? valid_123_1 : _GEN_631; // @[icache.scala 68:{25,25}]
  wire  _GEN_633 = 7'h7c == idx & ~way ? valid_124_0 : _GEN_632; // @[icache.scala 68:{25,25}]
  wire  _GEN_634 = 7'h7c == idx & way ? valid_124_1 : _GEN_633; // @[icache.scala 68:{25,25}]
  wire  _GEN_635 = 7'h7d == idx & ~way ? valid_125_0 : _GEN_634; // @[icache.scala 68:{25,25}]
  wire  _GEN_636 = 7'h7d == idx & way ? valid_125_1 : _GEN_635; // @[icache.scala 68:{25,25}]
  wire  _GEN_637 = 7'h7e == idx & ~way ? valid_126_0 : _GEN_636; // @[icache.scala 68:{25,25}]
  wire  _GEN_638 = 7'h7e == idx & way ? valid_126_1 : _GEN_637; // @[icache.scala 68:{25,25}]
  wire  _GEN_639 = 7'h7f == idx & ~way ? valid_127_0 : _GEN_638; // @[icache.scala 68:{25,25}]
  wire  _GEN_640 = 7'h7f == idx & way ? valid_127_1 : _GEN_639; // @[icache.scala 68:{25,25}]
  wire [41:0] _cache_tag_T_5 = {_GEN_127[41:21],tag}; // @[Cat.scala 33:92]
  wire [41:0] _cache_tag_T_7 = {tag,_GEN_127[20:0]}; // @[Cat.scala 33:92]
  wire  _addr_T = state == 2'h0; // @[icache.scala 71:26]
  wire  _addr_T_2 = state == 2'h1; // @[icache.scala 71:57]
  wire  _addr_T_3 = state == 2'h1 & req; // @[icache.scala 71:71]
  wire  _addr_T_4 = ~miss; // @[icache.scala 71:82]
  wire  _addr_T_6 = state == 2'h0 & req | state == 2'h1 & req & ~miss; // @[icache.scala 71:46]
  wire  _en_w_T = state == 2'h3; // @[icache.scala 81:20]
  wire  en_w = state == 2'h3 & _state_T_12; // @[icache.scala 81:35]
  wire [6:0] _GEN_1791 = {cnt, 6'h0}; // @[icache.scala 84:90]
  wire [7:0] _io_ram_bits_BWEN_T = {{1'd0}, _GEN_1791}; // @[icache.scala 84:90]
  wire [382:0] _io_ram_bits_BWEN_T_1 = 383'hffffffffffffffff << _io_ram_bits_BWEN_T; // @[icache.scala 84:82]
  wire [382:0] _io_ram_bits_BWEN_T_2 = ~_io_ram_bits_BWEN_T_1; // @[icache.scala 84:32]
  wire [382:0] _io_ram_bits_BWEN_T_4 = en_w ? _io_ram_bits_BWEN_T_2 : 383'hffffffffffffffffffffffffffffffff; // @[icache.scala 84:25]
  wire [127:0] _io_ram_bits_D_T = {64'h0,io_mem_r_bits_data}; // @[Cat.scala 33:92]
  wire [382:0] _GEN_0 = {{255'd0}, _io_ram_bits_D_T}; // @[icache.scala 86:62]
  wire [382:0] _io_ram_bits_D_T_2 = _GEN_0 << _io_ram_bits_BWEN_T; // @[icache.scala 86:62]
  wire [382:0] _io_ram_bits_D_T_3 = en_w ? _io_ram_bits_D_T_2 : 383'h0; // @[icache.scala 86:22]
  reg  flag; // @[icache.scala 89:20]
  reg [63:0] rdata; // @[icache.scala 90:21]
  wire  _flag_T_4 = en_w ? 1'h0 : flag; // @[icache.scala 92:14]
  wire [34:0] _GEN_1793 = {{3'd0}, addr}; // @[icache.scala 95:31]
  wire [34:0] _io_mem_ar_bits_addr_T_2 = _GEN_1793 & 35'h7fffffff8; // @[icache.scala 95:31]
  wire  _io_mem_ar_bits_len_T = uncache ? 1'h0 : 1'h1; // @[icache.scala 97:28]
  wire  _io_in_r_bits_data_T_2 = _addr_T_2 & _addr_T_4; // @[icache.scala 118:50]
  wire [127:0] _io_in_r_bits_data_T_3 = io_ram_bits_Q1 >> offset; // @[icache.scala 120:44]
  wire [127:0] _io_in_r_bits_data_T_5 = io_ram_bits_Q0 >> offset; // @[icache.scala 121:44]
  wire [63:0] _io_in_r_bits_data_T_7 = hit_way ? _io_in_r_bits_data_T_3[63:0] : _io_in_r_bits_data_T_5[63:0]; // @[icache.scala 119:30]
  wire [63:0] _io_in_r_bits_data_T_14 = rdata >> offset[5:0]; // @[icache.scala 125:37]
  wire [63:0] _io_in_r_bits_data_T_15 = uncache ? io_mem_r_bits_data : _io_in_r_bits_data_T_14; // @[icache.scala 123:32]
  wire [63:0] _io_in_r_bits_data_T_16 = en_w & io_mem_r_bits_last ? _io_in_r_bits_data_T_15 : 64'h0; // @[icache.scala 122:30]
  reg [31:0] hit_num; // @[icache.scala 135:22]
  reg [31:0] inst_num; // @[icache.scala 136:23]
  wire [31:0] _hit_num_T_4 = hit_num + 32'h1; // @[icache.scala 138:58]
  wire [31:0] _inst_num_T_4 = inst_num + 32'h1; // @[icache.scala 139:59]
  LFSR_8 lfsr8 ( // @[icache.scala 54:21]
    .clock(lfsr8_clock),
    .reset(lfsr8_reset),
    .io_en(lfsr8_io_en),
    .io_out(lfsr8_io_out)
  );
  assign io_in_ar_ready = _addr_T | _addr_T_2; // @[icache.scala 127:40]
  assign io_in_r_valid = _io_in_r_bits_data_T_2 | _state_T_14; // @[icache.scala 128:55]
  assign io_in_r_bits_data = _addr_T_2 & _addr_T_4 ? _io_in_r_bits_data_T_7 : _io_in_r_bits_data_T_16; // @[icache.scala 118:28]
  assign io_mem_ar_valid = state == 2'h2; // @[icache.scala 96:28]
  assign io_mem_ar_bits_addr = _io_mem_ar_bits_addr_T_2[31:0]; // @[icache.scala 95:23]
  assign io_mem_ar_bits_len = {{7'd0}, _io_mem_ar_bits_len_T}; // @[icache.scala 97:22]
  assign io_mem_r_ready = 1'h1; // @[icache.scala 102:18]
  assign io_ram_bits_CEN = ~(_addr_T | _addr_T_3 | _en_w_T); // @[icache.scala 82:21]
  assign io_ram_bits_WEN = ~en_w; // @[icache.scala 83:21]
  assign io_ram_bits_BWEN = _io_ram_bits_BWEN_T_4[127:0]; // @[icache.scala 84:19]
  assign io_ram_bits_A = en_w ? idx : io_in_ar_bits_addr[10:4]; // @[icache.scala 85:22]
  assign io_ram_bits_D = _io_ram_bits_D_T_3[127:0]; // @[icache.scala 86:16]
  assign io_ram_bits_WAY = way; // @[icache.scala 87:18]
  assign io_hitrate = {inst_num,hit_num}; // @[Cat.scala 33:92]
  assign lfsr8_clock = clock;
  assign lfsr8_reset = reset;
  assign lfsr8_io_en = state == 2'h2; // @[icache.scala 55:25]
  always @(posedge clock) begin
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_0 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h0 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_0 <= _cache_tag_T_5;
        end else begin
          cache_tag_0 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_0 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_0 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_1 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_1 <= _cache_tag_T_5;
        end else begin
          cache_tag_1 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_1 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_1 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_2 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_2 <= _cache_tag_T_5;
        end else begin
          cache_tag_2 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_2 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_2 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_3 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_3 <= _cache_tag_T_5;
        end else begin
          cache_tag_3 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_3 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_3 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_4 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_4 <= _cache_tag_T_5;
        end else begin
          cache_tag_4 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_4 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_4 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_5 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_5 <= _cache_tag_T_5;
        end else begin
          cache_tag_5 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_5 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_5 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_6 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_6 <= _cache_tag_T_5;
        end else begin
          cache_tag_6 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_6 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_6 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_7 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_7 <= _cache_tag_T_5;
        end else begin
          cache_tag_7 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_7 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_7 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_8 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h8 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_8 <= _cache_tag_T_5;
        end else begin
          cache_tag_8 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_8 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_8 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_9 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h9 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_9 <= _cache_tag_T_5;
        end else begin
          cache_tag_9 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_9 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_9 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_10 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'ha == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_10 <= _cache_tag_T_5;
        end else begin
          cache_tag_10 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_10 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_10 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_11 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'hb == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_11 <= _cache_tag_T_5;
        end else begin
          cache_tag_11 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_11 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_11 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_12 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'hc == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_12 <= _cache_tag_T_5;
        end else begin
          cache_tag_12 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_12 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_12 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_13 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'hd == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_13 <= _cache_tag_T_5;
        end else begin
          cache_tag_13 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_13 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_13 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_14 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'he == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_14 <= _cache_tag_T_5;
        end else begin
          cache_tag_14 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_14 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_14 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_15 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'hf == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_15 <= _cache_tag_T_5;
        end else begin
          cache_tag_15 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_15 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_15 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_16 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h10 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_16 <= _cache_tag_T_5;
        end else begin
          cache_tag_16 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_16 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_16 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_17 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h11 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_17 <= _cache_tag_T_5;
        end else begin
          cache_tag_17 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_17 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_17 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_18 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h12 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_18 <= _cache_tag_T_5;
        end else begin
          cache_tag_18 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_18 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_18 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_19 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h13 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_19 <= _cache_tag_T_5;
        end else begin
          cache_tag_19 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_19 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_19 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_20 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h14 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_20 <= _cache_tag_T_5;
        end else begin
          cache_tag_20 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_20 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_20 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_21 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h15 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_21 <= _cache_tag_T_5;
        end else begin
          cache_tag_21 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_21 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_21 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_22 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h16 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_22 <= _cache_tag_T_5;
        end else begin
          cache_tag_22 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_22 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_22 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_23 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h17 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_23 <= _cache_tag_T_5;
        end else begin
          cache_tag_23 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_23 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_23 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_24 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h18 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_24 <= _cache_tag_T_5;
        end else begin
          cache_tag_24 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_24 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_24 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_25 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h19 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_25 <= _cache_tag_T_5;
        end else begin
          cache_tag_25 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_25 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_25 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_26 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_26 <= _cache_tag_T_5;
        end else begin
          cache_tag_26 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_26 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_26 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_27 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_27 <= _cache_tag_T_5;
        end else begin
          cache_tag_27 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_27 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_27 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_28 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_28 <= _cache_tag_T_5;
        end else begin
          cache_tag_28 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_28 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_28 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_29 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_29 <= _cache_tag_T_5;
        end else begin
          cache_tag_29 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_29 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_29 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_30 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_30 <= _cache_tag_T_5;
        end else begin
          cache_tag_30 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_30 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_30 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_31 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h1f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_31 <= _cache_tag_T_5;
        end else begin
          cache_tag_31 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_31 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_31 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_32 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h20 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_32 <= _cache_tag_T_5;
        end else begin
          cache_tag_32 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_32 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_32 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_33 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h21 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_33 <= _cache_tag_T_5;
        end else begin
          cache_tag_33 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_33 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_33 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_34 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h22 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_34 <= _cache_tag_T_5;
        end else begin
          cache_tag_34 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_34 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_34 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_35 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h23 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_35 <= _cache_tag_T_5;
        end else begin
          cache_tag_35 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_35 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_35 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_36 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h24 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_36 <= _cache_tag_T_5;
        end else begin
          cache_tag_36 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_36 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_36 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_37 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h25 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_37 <= _cache_tag_T_5;
        end else begin
          cache_tag_37 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_37 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_37 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_38 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h26 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_38 <= _cache_tag_T_5;
        end else begin
          cache_tag_38 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_38 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_38 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_39 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h27 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_39 <= _cache_tag_T_5;
        end else begin
          cache_tag_39 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_39 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_39 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_40 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h28 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_40 <= _cache_tag_T_5;
        end else begin
          cache_tag_40 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_40 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_40 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_41 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h29 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_41 <= _cache_tag_T_5;
        end else begin
          cache_tag_41 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_41 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_41 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_42 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_42 <= _cache_tag_T_5;
        end else begin
          cache_tag_42 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_42 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_42 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_43 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_43 <= _cache_tag_T_5;
        end else begin
          cache_tag_43 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_43 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_43 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_44 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_44 <= _cache_tag_T_5;
        end else begin
          cache_tag_44 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_44 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_44 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_45 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_45 <= _cache_tag_T_5;
        end else begin
          cache_tag_45 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_45 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_45 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_46 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_46 <= _cache_tag_T_5;
        end else begin
          cache_tag_46 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_46 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_46 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_47 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h2f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_47 <= _cache_tag_T_5;
        end else begin
          cache_tag_47 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_47 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_47 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_48 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h30 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_48 <= _cache_tag_T_5;
        end else begin
          cache_tag_48 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_48 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_48 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_49 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h31 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_49 <= _cache_tag_T_5;
        end else begin
          cache_tag_49 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_49 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_49 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_50 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h32 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_50 <= _cache_tag_T_5;
        end else begin
          cache_tag_50 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_50 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_50 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_51 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h33 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_51 <= _cache_tag_T_5;
        end else begin
          cache_tag_51 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_51 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_51 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_52 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h34 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_52 <= _cache_tag_T_5;
        end else begin
          cache_tag_52 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_52 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_52 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_53 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h35 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_53 <= _cache_tag_T_5;
        end else begin
          cache_tag_53 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_53 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_53 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_54 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h36 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_54 <= _cache_tag_T_5;
        end else begin
          cache_tag_54 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_54 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_54 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_55 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h37 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_55 <= _cache_tag_T_5;
        end else begin
          cache_tag_55 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_55 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_55 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_56 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h38 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_56 <= _cache_tag_T_5;
        end else begin
          cache_tag_56 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_56 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_56 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_57 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h39 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_57 <= _cache_tag_T_5;
        end else begin
          cache_tag_57 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_57 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_57 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_58 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_58 <= _cache_tag_T_5;
        end else begin
          cache_tag_58 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_58 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_58 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_59 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_59 <= _cache_tag_T_5;
        end else begin
          cache_tag_59 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_59 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_59 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_60 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_60 <= _cache_tag_T_5;
        end else begin
          cache_tag_60 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_60 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_60 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_61 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_61 <= _cache_tag_T_5;
        end else begin
          cache_tag_61 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_61 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_61 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_62 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_62 <= _cache_tag_T_5;
        end else begin
          cache_tag_62 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_62 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_62 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_63 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h3f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_63 <= _cache_tag_T_5;
        end else begin
          cache_tag_63 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_63 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_63 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_64 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h40 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_64 <= _cache_tag_T_5;
        end else begin
          cache_tag_64 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_64 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_64 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_65 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h41 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_65 <= _cache_tag_T_5;
        end else begin
          cache_tag_65 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_65 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_65 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_66 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h42 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_66 <= _cache_tag_T_5;
        end else begin
          cache_tag_66 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_66 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_66 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_67 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h43 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_67 <= _cache_tag_T_5;
        end else begin
          cache_tag_67 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_67 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_67 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_68 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h44 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_68 <= _cache_tag_T_5;
        end else begin
          cache_tag_68 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_68 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_68 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_69 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h45 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_69 <= _cache_tag_T_5;
        end else begin
          cache_tag_69 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_69 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_69 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_70 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h46 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_70 <= _cache_tag_T_5;
        end else begin
          cache_tag_70 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_70 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_70 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_71 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h47 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_71 <= _cache_tag_T_5;
        end else begin
          cache_tag_71 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_71 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_71 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_72 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h48 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_72 <= _cache_tag_T_5;
        end else begin
          cache_tag_72 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_72 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_72 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_73 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h49 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_73 <= _cache_tag_T_5;
        end else begin
          cache_tag_73 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_73 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_73 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_74 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_74 <= _cache_tag_T_5;
        end else begin
          cache_tag_74 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_74 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_74 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_75 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_75 <= _cache_tag_T_5;
        end else begin
          cache_tag_75 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_75 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_75 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_76 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_76 <= _cache_tag_T_5;
        end else begin
          cache_tag_76 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_76 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_76 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_77 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_77 <= _cache_tag_T_5;
        end else begin
          cache_tag_77 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_77 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_77 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_78 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_78 <= _cache_tag_T_5;
        end else begin
          cache_tag_78 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_78 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_78 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_79 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h4f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_79 <= _cache_tag_T_5;
        end else begin
          cache_tag_79 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_79 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_79 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_80 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h50 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_80 <= _cache_tag_T_5;
        end else begin
          cache_tag_80 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_80 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_80 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_81 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h51 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_81 <= _cache_tag_T_5;
        end else begin
          cache_tag_81 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_81 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_81 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_82 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h52 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_82 <= _cache_tag_T_5;
        end else begin
          cache_tag_82 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_82 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_82 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_83 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h53 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_83 <= _cache_tag_T_5;
        end else begin
          cache_tag_83 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_83 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_83 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_84 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h54 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_84 <= _cache_tag_T_5;
        end else begin
          cache_tag_84 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_84 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_84 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_85 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h55 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_85 <= _cache_tag_T_5;
        end else begin
          cache_tag_85 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_85 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_85 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_86 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h56 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_86 <= _cache_tag_T_5;
        end else begin
          cache_tag_86 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_86 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_86 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_87 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h57 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_87 <= _cache_tag_T_5;
        end else begin
          cache_tag_87 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_87 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_87 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_88 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h58 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_88 <= _cache_tag_T_5;
        end else begin
          cache_tag_88 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_88 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_88 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_89 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h59 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_89 <= _cache_tag_T_5;
        end else begin
          cache_tag_89 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_89 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_89 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_90 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_90 <= _cache_tag_T_5;
        end else begin
          cache_tag_90 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_90 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_90 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_91 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_91 <= _cache_tag_T_5;
        end else begin
          cache_tag_91 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_91 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_91 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_92 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_92 <= _cache_tag_T_5;
        end else begin
          cache_tag_92 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_92 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_92 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_93 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_93 <= _cache_tag_T_5;
        end else begin
          cache_tag_93 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_93 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_93 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_94 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_94 <= _cache_tag_T_5;
        end else begin
          cache_tag_94 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_94 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_94 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_95 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h5f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_95 <= _cache_tag_T_5;
        end else begin
          cache_tag_95 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_95 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_95 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_96 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h60 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_96 <= _cache_tag_T_5;
        end else begin
          cache_tag_96 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_96 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_96 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_97 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h61 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_97 <= _cache_tag_T_5;
        end else begin
          cache_tag_97 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_97 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_97 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_98 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h62 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_98 <= _cache_tag_T_5;
        end else begin
          cache_tag_98 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_98 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_98 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_99 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h63 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_99 <= _cache_tag_T_5;
        end else begin
          cache_tag_99 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_99 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_99 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_100 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h64 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_100 <= _cache_tag_T_5;
        end else begin
          cache_tag_100 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_100 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_100 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_101 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h65 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_101 <= _cache_tag_T_5;
        end else begin
          cache_tag_101 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_101 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_101 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_102 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h66 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_102 <= _cache_tag_T_5;
        end else begin
          cache_tag_102 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_102 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_102 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_103 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h67 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_103 <= _cache_tag_T_5;
        end else begin
          cache_tag_103 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_103 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_103 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_104 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h68 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_104 <= _cache_tag_T_5;
        end else begin
          cache_tag_104 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_104 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_104 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_105 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h69 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_105 <= _cache_tag_T_5;
        end else begin
          cache_tag_105 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_105 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_105 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_106 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_106 <= _cache_tag_T_5;
        end else begin
          cache_tag_106 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_106 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_106 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_107 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_107 <= _cache_tag_T_5;
        end else begin
          cache_tag_107 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_107 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_107 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_108 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_108 <= _cache_tag_T_5;
        end else begin
          cache_tag_108 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_108 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_108 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_109 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_109 <= _cache_tag_T_5;
        end else begin
          cache_tag_109 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_109 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_109 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_110 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_110 <= _cache_tag_T_5;
        end else begin
          cache_tag_110 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_110 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_110 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_111 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h6f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_111 <= _cache_tag_T_5;
        end else begin
          cache_tag_111 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_111 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_111 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_112 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h70 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_112 <= _cache_tag_T_5;
        end else begin
          cache_tag_112 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_112 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_112 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_113 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h71 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_113 <= _cache_tag_T_5;
        end else begin
          cache_tag_113 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_113 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_113 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_114 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h72 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_114 <= _cache_tag_T_5;
        end else begin
          cache_tag_114 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_114 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_114 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_115 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h73 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_115 <= _cache_tag_T_5;
        end else begin
          cache_tag_115 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_115 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_115 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_116 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h74 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_116 <= _cache_tag_T_5;
        end else begin
          cache_tag_116 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_116 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_116 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_117 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h75 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_117 <= _cache_tag_T_5;
        end else begin
          cache_tag_117 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_117 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_117 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_118 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h76 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_118 <= _cache_tag_T_5;
        end else begin
          cache_tag_118 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_118 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_118 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_119 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h77 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_119 <= _cache_tag_T_5;
        end else begin
          cache_tag_119 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_119 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_119 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_120 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h78 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_120 <= _cache_tag_T_5;
        end else begin
          cache_tag_120 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_120 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_120 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_121 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h79 == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_121 <= _cache_tag_T_5;
        end else begin
          cache_tag_121 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_121 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_121 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_122 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7a == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_122 <= _cache_tag_T_5;
        end else begin
          cache_tag_122 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_122 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_122 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_123 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7b == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_123 <= _cache_tag_T_5;
        end else begin
          cache_tag_123 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_123 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_123 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_124 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7c == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_124 <= _cache_tag_T_5;
        end else begin
          cache_tag_124 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_124 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_124 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_125 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7d == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_125 <= _cache_tag_T_5;
        end else begin
          cache_tag_125 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_125 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_125 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_126 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7e == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_126 <= _cache_tag_T_5;
        end else begin
          cache_tag_126 <= _cache_tag_T_7;
        end
      end else if (7'h7f == idx) begin // @[icache.scala 50:33]
        cache_tag_126 <= cache_tag_127; // @[icache.scala 50:33]
      end else begin
        cache_tag_126 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 30:26]
      cache_tag_127 <= 42'h0; // @[icache.scala 30:26]
    end else if (7'h7f == idx) begin // @[icache.scala 69:18]
      if (_valid_T_2) begin // @[icache.scala 69:24]
        if (_GEN_1027) begin // @[icache.scala 69:58]
          cache_tag_127 <= _cache_tag_T_5;
        end else begin
          cache_tag_127 <= _cache_tag_T_7;
        end
      end else if (!(7'h7f == idx)) begin // @[icache.scala 50:33]
        cache_tag_127 <= _GEN_126;
      end
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_0_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h0 == idx & ~way) begin // @[icache.scala 68:19]
      valid_0_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_0_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h0 == idx & way) begin // @[icache.scala 68:19]
      valid_0_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_1_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1 == idx & ~way) begin // @[icache.scala 68:19]
      valid_1_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_1_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1 == idx & way) begin // @[icache.scala 68:19]
      valid_1_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_2_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2 == idx & ~way) begin // @[icache.scala 68:19]
      valid_2_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_2_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2 == idx & way) begin // @[icache.scala 68:19]
      valid_2_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_3_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3 == idx & ~way) begin // @[icache.scala 68:19]
      valid_3_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_3_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3 == idx & way) begin // @[icache.scala 68:19]
      valid_3_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_4_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4 == idx & ~way) begin // @[icache.scala 68:19]
      valid_4_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_4_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4 == idx & way) begin // @[icache.scala 68:19]
      valid_4_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_5_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5 == idx & ~way) begin // @[icache.scala 68:19]
      valid_5_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_5_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5 == idx & way) begin // @[icache.scala 68:19]
      valid_5_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_6_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6 == idx & ~way) begin // @[icache.scala 68:19]
      valid_6_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_6_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6 == idx & way) begin // @[icache.scala 68:19]
      valid_6_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_7_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7 == idx & ~way) begin // @[icache.scala 68:19]
      valid_7_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_7_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7 == idx & way) begin // @[icache.scala 68:19]
      valid_7_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_8_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h8 == idx & ~way) begin // @[icache.scala 68:19]
      valid_8_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_8_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h8 == idx & way) begin // @[icache.scala 68:19]
      valid_8_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_9_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h9 == idx & ~way) begin // @[icache.scala 68:19]
      valid_9_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_9_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h9 == idx & way) begin // @[icache.scala 68:19]
      valid_9_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_10_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'ha == idx & ~way) begin // @[icache.scala 68:19]
      valid_10_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_10_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'ha == idx & way) begin // @[icache.scala 68:19]
      valid_10_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_11_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hb == idx & ~way) begin // @[icache.scala 68:19]
      valid_11_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_11_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hb == idx & way) begin // @[icache.scala 68:19]
      valid_11_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_12_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hc == idx & ~way) begin // @[icache.scala 68:19]
      valid_12_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_12_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hc == idx & way) begin // @[icache.scala 68:19]
      valid_12_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_13_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hd == idx & ~way) begin // @[icache.scala 68:19]
      valid_13_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_13_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hd == idx & way) begin // @[icache.scala 68:19]
      valid_13_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_14_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'he == idx & ~way) begin // @[icache.scala 68:19]
      valid_14_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_14_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'he == idx & way) begin // @[icache.scala 68:19]
      valid_14_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_15_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hf == idx & ~way) begin // @[icache.scala 68:19]
      valid_15_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_15_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'hf == idx & way) begin // @[icache.scala 68:19]
      valid_15_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_16_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h10 == idx & ~way) begin // @[icache.scala 68:19]
      valid_16_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_16_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h10 == idx & way) begin // @[icache.scala 68:19]
      valid_16_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_17_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h11 == idx & ~way) begin // @[icache.scala 68:19]
      valid_17_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_17_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h11 == idx & way) begin // @[icache.scala 68:19]
      valid_17_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_18_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h12 == idx & ~way) begin // @[icache.scala 68:19]
      valid_18_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_18_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h12 == idx & way) begin // @[icache.scala 68:19]
      valid_18_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_19_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h13 == idx & ~way) begin // @[icache.scala 68:19]
      valid_19_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_19_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h13 == idx & way) begin // @[icache.scala 68:19]
      valid_19_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_20_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h14 == idx & ~way) begin // @[icache.scala 68:19]
      valid_20_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_20_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h14 == idx & way) begin // @[icache.scala 68:19]
      valid_20_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_21_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h15 == idx & ~way) begin // @[icache.scala 68:19]
      valid_21_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_21_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h15 == idx & way) begin // @[icache.scala 68:19]
      valid_21_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_22_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h16 == idx & ~way) begin // @[icache.scala 68:19]
      valid_22_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_22_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h16 == idx & way) begin // @[icache.scala 68:19]
      valid_22_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_23_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h17 == idx & ~way) begin // @[icache.scala 68:19]
      valid_23_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_23_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h17 == idx & way) begin // @[icache.scala 68:19]
      valid_23_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_24_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h18 == idx & ~way) begin // @[icache.scala 68:19]
      valid_24_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_24_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h18 == idx & way) begin // @[icache.scala 68:19]
      valid_24_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_25_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h19 == idx & ~way) begin // @[icache.scala 68:19]
      valid_25_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_25_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h19 == idx & way) begin // @[icache.scala 68:19]
      valid_25_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_26_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1a == idx & ~way) begin // @[icache.scala 68:19]
      valid_26_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_26_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1a == idx & way) begin // @[icache.scala 68:19]
      valid_26_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_27_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1b == idx & ~way) begin // @[icache.scala 68:19]
      valid_27_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_27_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1b == idx & way) begin // @[icache.scala 68:19]
      valid_27_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_28_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1c == idx & ~way) begin // @[icache.scala 68:19]
      valid_28_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_28_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1c == idx & way) begin // @[icache.scala 68:19]
      valid_28_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_29_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1d == idx & ~way) begin // @[icache.scala 68:19]
      valid_29_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_29_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1d == idx & way) begin // @[icache.scala 68:19]
      valid_29_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_30_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1e == idx & ~way) begin // @[icache.scala 68:19]
      valid_30_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_30_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1e == idx & way) begin // @[icache.scala 68:19]
      valid_30_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_31_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1f == idx & ~way) begin // @[icache.scala 68:19]
      valid_31_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_31_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h1f == idx & way) begin // @[icache.scala 68:19]
      valid_31_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_32_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h20 == idx & ~way) begin // @[icache.scala 68:19]
      valid_32_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_32_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h20 == idx & way) begin // @[icache.scala 68:19]
      valid_32_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_33_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h21 == idx & ~way) begin // @[icache.scala 68:19]
      valid_33_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_33_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h21 == idx & way) begin // @[icache.scala 68:19]
      valid_33_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_34_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h22 == idx & ~way) begin // @[icache.scala 68:19]
      valid_34_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_34_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h22 == idx & way) begin // @[icache.scala 68:19]
      valid_34_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_35_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h23 == idx & ~way) begin // @[icache.scala 68:19]
      valid_35_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_35_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h23 == idx & way) begin // @[icache.scala 68:19]
      valid_35_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_36_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h24 == idx & ~way) begin // @[icache.scala 68:19]
      valid_36_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_36_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h24 == idx & way) begin // @[icache.scala 68:19]
      valid_36_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_37_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h25 == idx & ~way) begin // @[icache.scala 68:19]
      valid_37_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_37_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h25 == idx & way) begin // @[icache.scala 68:19]
      valid_37_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_38_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h26 == idx & ~way) begin // @[icache.scala 68:19]
      valid_38_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_38_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h26 == idx & way) begin // @[icache.scala 68:19]
      valid_38_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_39_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h27 == idx & ~way) begin // @[icache.scala 68:19]
      valid_39_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_39_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h27 == idx & way) begin // @[icache.scala 68:19]
      valid_39_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_40_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h28 == idx & ~way) begin // @[icache.scala 68:19]
      valid_40_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_40_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h28 == idx & way) begin // @[icache.scala 68:19]
      valid_40_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_41_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h29 == idx & ~way) begin // @[icache.scala 68:19]
      valid_41_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_41_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h29 == idx & way) begin // @[icache.scala 68:19]
      valid_41_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_42_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2a == idx & ~way) begin // @[icache.scala 68:19]
      valid_42_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_42_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2a == idx & way) begin // @[icache.scala 68:19]
      valid_42_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_43_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2b == idx & ~way) begin // @[icache.scala 68:19]
      valid_43_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_43_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2b == idx & way) begin // @[icache.scala 68:19]
      valid_43_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_44_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2c == idx & ~way) begin // @[icache.scala 68:19]
      valid_44_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_44_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2c == idx & way) begin // @[icache.scala 68:19]
      valid_44_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_45_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2d == idx & ~way) begin // @[icache.scala 68:19]
      valid_45_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_45_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2d == idx & way) begin // @[icache.scala 68:19]
      valid_45_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_46_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2e == idx & ~way) begin // @[icache.scala 68:19]
      valid_46_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_46_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2e == idx & way) begin // @[icache.scala 68:19]
      valid_46_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_47_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2f == idx & ~way) begin // @[icache.scala 68:19]
      valid_47_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_47_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h2f == idx & way) begin // @[icache.scala 68:19]
      valid_47_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_48_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h30 == idx & ~way) begin // @[icache.scala 68:19]
      valid_48_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_48_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h30 == idx & way) begin // @[icache.scala 68:19]
      valid_48_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_49_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h31 == idx & ~way) begin // @[icache.scala 68:19]
      valid_49_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_49_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h31 == idx & way) begin // @[icache.scala 68:19]
      valid_49_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_50_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h32 == idx & ~way) begin // @[icache.scala 68:19]
      valid_50_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_50_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h32 == idx & way) begin // @[icache.scala 68:19]
      valid_50_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_51_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h33 == idx & ~way) begin // @[icache.scala 68:19]
      valid_51_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_51_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h33 == idx & way) begin // @[icache.scala 68:19]
      valid_51_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_52_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h34 == idx & ~way) begin // @[icache.scala 68:19]
      valid_52_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_52_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h34 == idx & way) begin // @[icache.scala 68:19]
      valid_52_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_53_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h35 == idx & ~way) begin // @[icache.scala 68:19]
      valid_53_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_53_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h35 == idx & way) begin // @[icache.scala 68:19]
      valid_53_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_54_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h36 == idx & ~way) begin // @[icache.scala 68:19]
      valid_54_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_54_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h36 == idx & way) begin // @[icache.scala 68:19]
      valid_54_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_55_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h37 == idx & ~way) begin // @[icache.scala 68:19]
      valid_55_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_55_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h37 == idx & way) begin // @[icache.scala 68:19]
      valid_55_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_56_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h38 == idx & ~way) begin // @[icache.scala 68:19]
      valid_56_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_56_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h38 == idx & way) begin // @[icache.scala 68:19]
      valid_56_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_57_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h39 == idx & ~way) begin // @[icache.scala 68:19]
      valid_57_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_57_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h39 == idx & way) begin // @[icache.scala 68:19]
      valid_57_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_58_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3a == idx & ~way) begin // @[icache.scala 68:19]
      valid_58_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_58_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3a == idx & way) begin // @[icache.scala 68:19]
      valid_58_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_59_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3b == idx & ~way) begin // @[icache.scala 68:19]
      valid_59_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_59_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3b == idx & way) begin // @[icache.scala 68:19]
      valid_59_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_60_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3c == idx & ~way) begin // @[icache.scala 68:19]
      valid_60_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_60_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3c == idx & way) begin // @[icache.scala 68:19]
      valid_60_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_61_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3d == idx & ~way) begin // @[icache.scala 68:19]
      valid_61_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_61_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3d == idx & way) begin // @[icache.scala 68:19]
      valid_61_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_62_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3e == idx & ~way) begin // @[icache.scala 68:19]
      valid_62_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_62_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3e == idx & way) begin // @[icache.scala 68:19]
      valid_62_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_63_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3f == idx & ~way) begin // @[icache.scala 68:19]
      valid_63_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_63_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h3f == idx & way) begin // @[icache.scala 68:19]
      valid_63_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_64_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h40 == idx & ~way) begin // @[icache.scala 68:19]
      valid_64_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_64_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h40 == idx & way) begin // @[icache.scala 68:19]
      valid_64_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_65_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h41 == idx & ~way) begin // @[icache.scala 68:19]
      valid_65_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_65_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h41 == idx & way) begin // @[icache.scala 68:19]
      valid_65_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_66_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h42 == idx & ~way) begin // @[icache.scala 68:19]
      valid_66_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_66_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h42 == idx & way) begin // @[icache.scala 68:19]
      valid_66_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_67_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h43 == idx & ~way) begin // @[icache.scala 68:19]
      valid_67_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_67_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h43 == idx & way) begin // @[icache.scala 68:19]
      valid_67_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_68_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h44 == idx & ~way) begin // @[icache.scala 68:19]
      valid_68_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_68_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h44 == idx & way) begin // @[icache.scala 68:19]
      valid_68_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_69_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h45 == idx & ~way) begin // @[icache.scala 68:19]
      valid_69_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_69_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h45 == idx & way) begin // @[icache.scala 68:19]
      valid_69_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_70_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h46 == idx & ~way) begin // @[icache.scala 68:19]
      valid_70_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_70_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h46 == idx & way) begin // @[icache.scala 68:19]
      valid_70_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_71_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h47 == idx & ~way) begin // @[icache.scala 68:19]
      valid_71_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_71_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h47 == idx & way) begin // @[icache.scala 68:19]
      valid_71_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_72_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h48 == idx & ~way) begin // @[icache.scala 68:19]
      valid_72_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_72_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h48 == idx & way) begin // @[icache.scala 68:19]
      valid_72_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_73_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h49 == idx & ~way) begin // @[icache.scala 68:19]
      valid_73_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_73_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h49 == idx & way) begin // @[icache.scala 68:19]
      valid_73_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_74_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4a == idx & ~way) begin // @[icache.scala 68:19]
      valid_74_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_74_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4a == idx & way) begin // @[icache.scala 68:19]
      valid_74_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_75_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4b == idx & ~way) begin // @[icache.scala 68:19]
      valid_75_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_75_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4b == idx & way) begin // @[icache.scala 68:19]
      valid_75_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_76_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4c == idx & ~way) begin // @[icache.scala 68:19]
      valid_76_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_76_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4c == idx & way) begin // @[icache.scala 68:19]
      valid_76_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_77_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4d == idx & ~way) begin // @[icache.scala 68:19]
      valid_77_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_77_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4d == idx & way) begin // @[icache.scala 68:19]
      valid_77_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_78_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4e == idx & ~way) begin // @[icache.scala 68:19]
      valid_78_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_78_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4e == idx & way) begin // @[icache.scala 68:19]
      valid_78_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_79_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4f == idx & ~way) begin // @[icache.scala 68:19]
      valid_79_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_79_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h4f == idx & way) begin // @[icache.scala 68:19]
      valid_79_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_80_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h50 == idx & ~way) begin // @[icache.scala 68:19]
      valid_80_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_80_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h50 == idx & way) begin // @[icache.scala 68:19]
      valid_80_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_81_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h51 == idx & ~way) begin // @[icache.scala 68:19]
      valid_81_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_81_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h51 == idx & way) begin // @[icache.scala 68:19]
      valid_81_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_82_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h52 == idx & ~way) begin // @[icache.scala 68:19]
      valid_82_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_82_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h52 == idx & way) begin // @[icache.scala 68:19]
      valid_82_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_83_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h53 == idx & ~way) begin // @[icache.scala 68:19]
      valid_83_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_83_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h53 == idx & way) begin // @[icache.scala 68:19]
      valid_83_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_84_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h54 == idx & ~way) begin // @[icache.scala 68:19]
      valid_84_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_84_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h54 == idx & way) begin // @[icache.scala 68:19]
      valid_84_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_85_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h55 == idx & ~way) begin // @[icache.scala 68:19]
      valid_85_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_85_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h55 == idx & way) begin // @[icache.scala 68:19]
      valid_85_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_86_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h56 == idx & ~way) begin // @[icache.scala 68:19]
      valid_86_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_86_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h56 == idx & way) begin // @[icache.scala 68:19]
      valid_86_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_87_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h57 == idx & ~way) begin // @[icache.scala 68:19]
      valid_87_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_87_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h57 == idx & way) begin // @[icache.scala 68:19]
      valid_87_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_88_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h58 == idx & ~way) begin // @[icache.scala 68:19]
      valid_88_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_88_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h58 == idx & way) begin // @[icache.scala 68:19]
      valid_88_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_89_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h59 == idx & ~way) begin // @[icache.scala 68:19]
      valid_89_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_89_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h59 == idx & way) begin // @[icache.scala 68:19]
      valid_89_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_90_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5a == idx & ~way) begin // @[icache.scala 68:19]
      valid_90_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_90_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5a == idx & way) begin // @[icache.scala 68:19]
      valid_90_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_91_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5b == idx & ~way) begin // @[icache.scala 68:19]
      valid_91_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_91_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5b == idx & way) begin // @[icache.scala 68:19]
      valid_91_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_92_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5c == idx & ~way) begin // @[icache.scala 68:19]
      valid_92_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_92_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5c == idx & way) begin // @[icache.scala 68:19]
      valid_92_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_93_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5d == idx & ~way) begin // @[icache.scala 68:19]
      valid_93_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_93_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5d == idx & way) begin // @[icache.scala 68:19]
      valid_93_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_94_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5e == idx & ~way) begin // @[icache.scala 68:19]
      valid_94_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_94_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5e == idx & way) begin // @[icache.scala 68:19]
      valid_94_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_95_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5f == idx & ~way) begin // @[icache.scala 68:19]
      valid_95_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_95_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h5f == idx & way) begin // @[icache.scala 68:19]
      valid_95_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_96_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h60 == idx & ~way) begin // @[icache.scala 68:19]
      valid_96_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_96_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h60 == idx & way) begin // @[icache.scala 68:19]
      valid_96_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_97_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h61 == idx & ~way) begin // @[icache.scala 68:19]
      valid_97_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_97_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h61 == idx & way) begin // @[icache.scala 68:19]
      valid_97_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_98_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h62 == idx & ~way) begin // @[icache.scala 68:19]
      valid_98_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_98_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h62 == idx & way) begin // @[icache.scala 68:19]
      valid_98_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_99_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h63 == idx & ~way) begin // @[icache.scala 68:19]
      valid_99_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_99_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h63 == idx & way) begin // @[icache.scala 68:19]
      valid_99_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_100_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h64 == idx & ~way) begin // @[icache.scala 68:19]
      valid_100_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_100_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h64 == idx & way) begin // @[icache.scala 68:19]
      valid_100_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_101_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h65 == idx & ~way) begin // @[icache.scala 68:19]
      valid_101_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_101_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h65 == idx & way) begin // @[icache.scala 68:19]
      valid_101_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_102_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h66 == idx & ~way) begin // @[icache.scala 68:19]
      valid_102_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_102_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h66 == idx & way) begin // @[icache.scala 68:19]
      valid_102_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_103_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h67 == idx & ~way) begin // @[icache.scala 68:19]
      valid_103_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_103_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h67 == idx & way) begin // @[icache.scala 68:19]
      valid_103_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_104_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h68 == idx & ~way) begin // @[icache.scala 68:19]
      valid_104_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_104_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h68 == idx & way) begin // @[icache.scala 68:19]
      valid_104_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_105_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h69 == idx & ~way) begin // @[icache.scala 68:19]
      valid_105_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_105_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h69 == idx & way) begin // @[icache.scala 68:19]
      valid_105_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_106_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6a == idx & ~way) begin // @[icache.scala 68:19]
      valid_106_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_106_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6a == idx & way) begin // @[icache.scala 68:19]
      valid_106_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_107_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6b == idx & ~way) begin // @[icache.scala 68:19]
      valid_107_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_107_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6b == idx & way) begin // @[icache.scala 68:19]
      valid_107_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_108_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6c == idx & ~way) begin // @[icache.scala 68:19]
      valid_108_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_108_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6c == idx & way) begin // @[icache.scala 68:19]
      valid_108_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_109_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6d == idx & ~way) begin // @[icache.scala 68:19]
      valid_109_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_109_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6d == idx & way) begin // @[icache.scala 68:19]
      valid_109_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_110_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6e == idx & ~way) begin // @[icache.scala 68:19]
      valid_110_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_110_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6e == idx & way) begin // @[icache.scala 68:19]
      valid_110_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_111_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6f == idx & ~way) begin // @[icache.scala 68:19]
      valid_111_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_111_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h6f == idx & way) begin // @[icache.scala 68:19]
      valid_111_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_112_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h70 == idx & ~way) begin // @[icache.scala 68:19]
      valid_112_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_112_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h70 == idx & way) begin // @[icache.scala 68:19]
      valid_112_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_113_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h71 == idx & ~way) begin // @[icache.scala 68:19]
      valid_113_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_113_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h71 == idx & way) begin // @[icache.scala 68:19]
      valid_113_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_114_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h72 == idx & ~way) begin // @[icache.scala 68:19]
      valid_114_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_114_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h72 == idx & way) begin // @[icache.scala 68:19]
      valid_114_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_115_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h73 == idx & ~way) begin // @[icache.scala 68:19]
      valid_115_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_115_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h73 == idx & way) begin // @[icache.scala 68:19]
      valid_115_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_116_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h74 == idx & ~way) begin // @[icache.scala 68:19]
      valid_116_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_116_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h74 == idx & way) begin // @[icache.scala 68:19]
      valid_116_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_117_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h75 == idx & ~way) begin // @[icache.scala 68:19]
      valid_117_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_117_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h75 == idx & way) begin // @[icache.scala 68:19]
      valid_117_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_118_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h76 == idx & ~way) begin // @[icache.scala 68:19]
      valid_118_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_118_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h76 == idx & way) begin // @[icache.scala 68:19]
      valid_118_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_119_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h77 == idx & ~way) begin // @[icache.scala 68:19]
      valid_119_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_119_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h77 == idx & way) begin // @[icache.scala 68:19]
      valid_119_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_120_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h78 == idx & ~way) begin // @[icache.scala 68:19]
      valid_120_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_120_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h78 == idx & way) begin // @[icache.scala 68:19]
      valid_120_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_121_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h79 == idx & ~way) begin // @[icache.scala 68:19]
      valid_121_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_121_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h79 == idx & way) begin // @[icache.scala 68:19]
      valid_121_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_122_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7a == idx & ~way) begin // @[icache.scala 68:19]
      valid_122_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_122_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7a == idx & way) begin // @[icache.scala 68:19]
      valid_122_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_123_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7b == idx & ~way) begin // @[icache.scala 68:19]
      valid_123_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_123_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7b == idx & way) begin // @[icache.scala 68:19]
      valid_123_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_124_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7c == idx & ~way) begin // @[icache.scala 68:19]
      valid_124_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_124_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7c == idx & way) begin // @[icache.scala 68:19]
      valid_124_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_125_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7d == idx & ~way) begin // @[icache.scala 68:19]
      valid_125_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_125_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7d == idx & way) begin // @[icache.scala 68:19]
      valid_125_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_126_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7e == idx & ~way) begin // @[icache.scala 68:19]
      valid_126_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_126_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7e == idx & way) begin // @[icache.scala 68:19]
      valid_126_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_127_0 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7f == idx & ~way) begin // @[icache.scala 68:19]
      valid_127_0 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 31:22]
      valid_127_1 <= 1'h0; // @[icache.scala 31:22]
    end else if (7'h7f == idx & way) begin // @[icache.scala 68:19]
      valid_127_1 <= _lfsr8_io_en_T & ~uncache | _GEN_640; // @[icache.scala 68:19]
    end
    if (reset) begin // @[icache.scala 36:22]
      state <= 2'h0; // @[icache.scala 36:22]
    end else if (2'h3 == state) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[icache.scala 65:22]
        state <= 2'h0;
      end else if (_state_T_12 & io_mem_r_bits_last) begin // @[icache.scala 65:49]
        state <= 2'h0;
      end else begin
        state <= 2'h3;
      end
    end else if (2'h2 == state) begin // @[Mux.scala 81:58]
      if (io_flush) begin // @[icache.scala 64:22]
        state <= 2'h0;
      end else begin
        state <= _state_T_9;
      end
    end else if (2'h1 == state) begin // @[Mux.scala 81:58]
      state <= _state_T_6;
    end else begin
      state <= _state_T_2;
    end
    if (reset) begin // @[icache.scala 39:21]
      addr <= 32'h0; // @[icache.scala 39:21]
    end else if (state == 2'h0 & req | state == 2'h1 & req & ~miss) begin // @[icache.scala 71:17]
      addr <= io_in_ar_bits_addr;
    end
    if (reset) begin // @[icache.scala 40:24]
      uncache <= 1'h0; // @[icache.scala 40:24]
    end else if (_addr_T_6) begin // @[icache.scala 72:17]
      uncache <= io_in_ar_bits_addr >= 32'ha0000000;
    end
    if (reset) begin // @[Reg.scala 35:20]
      way <= 1'h0; // @[Reg.scala 35:20]
    end else if (miss) begin // @[Reg.scala 36:18]
      way <= lfsr8_io_out[0]; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[icache.scala 58:20]
      cnt <= 1'h0; // @[icache.scala 58:20]
    end else if (_lfsr8_io_en_T) begin // @[icache.scala 76:13]
      cnt <= addr[3];
    end else if (_state_T_12) begin // @[icache.scala 77:13]
      cnt <= ~cnt;
    end
    if (reset) begin // @[icache.scala 89:20]
      flag <= 1'h0; // @[icache.scala 89:20]
    end else begin
      flag <= _addr_T | _flag_T_4; // @[icache.scala 91:8]
    end
    if (reset) begin // @[icache.scala 90:21]
      rdata <= 64'h0; // @[icache.scala 90:21]
    end else if (en_w & flag) begin // @[icache.scala 93:14]
      rdata <= io_mem_r_bits_data;
    end
    if (reset) begin // @[icache.scala 135:22]
      hit_num <= 32'h0; // @[icache.scala 135:22]
    end else if (_io_in_r_bits_data_T_2) begin // @[icache.scala 138:17]
      hit_num <= _hit_num_T_4;
    end
    if (reset) begin // @[icache.scala 136:23]
      inst_num <= 32'h0; // @[icache.scala 136:23]
    end else if (req) begin // @[icache.scala 139:18]
      inst_num <= _inst_num_T_4;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cache_tag_0 = _RAND_0[41:0];
  _RAND_1 = {2{`RANDOM}};
  cache_tag_1 = _RAND_1[41:0];
  _RAND_2 = {2{`RANDOM}};
  cache_tag_2 = _RAND_2[41:0];
  _RAND_3 = {2{`RANDOM}};
  cache_tag_3 = _RAND_3[41:0];
  _RAND_4 = {2{`RANDOM}};
  cache_tag_4 = _RAND_4[41:0];
  _RAND_5 = {2{`RANDOM}};
  cache_tag_5 = _RAND_5[41:0];
  _RAND_6 = {2{`RANDOM}};
  cache_tag_6 = _RAND_6[41:0];
  _RAND_7 = {2{`RANDOM}};
  cache_tag_7 = _RAND_7[41:0];
  _RAND_8 = {2{`RANDOM}};
  cache_tag_8 = _RAND_8[41:0];
  _RAND_9 = {2{`RANDOM}};
  cache_tag_9 = _RAND_9[41:0];
  _RAND_10 = {2{`RANDOM}};
  cache_tag_10 = _RAND_10[41:0];
  _RAND_11 = {2{`RANDOM}};
  cache_tag_11 = _RAND_11[41:0];
  _RAND_12 = {2{`RANDOM}};
  cache_tag_12 = _RAND_12[41:0];
  _RAND_13 = {2{`RANDOM}};
  cache_tag_13 = _RAND_13[41:0];
  _RAND_14 = {2{`RANDOM}};
  cache_tag_14 = _RAND_14[41:0];
  _RAND_15 = {2{`RANDOM}};
  cache_tag_15 = _RAND_15[41:0];
  _RAND_16 = {2{`RANDOM}};
  cache_tag_16 = _RAND_16[41:0];
  _RAND_17 = {2{`RANDOM}};
  cache_tag_17 = _RAND_17[41:0];
  _RAND_18 = {2{`RANDOM}};
  cache_tag_18 = _RAND_18[41:0];
  _RAND_19 = {2{`RANDOM}};
  cache_tag_19 = _RAND_19[41:0];
  _RAND_20 = {2{`RANDOM}};
  cache_tag_20 = _RAND_20[41:0];
  _RAND_21 = {2{`RANDOM}};
  cache_tag_21 = _RAND_21[41:0];
  _RAND_22 = {2{`RANDOM}};
  cache_tag_22 = _RAND_22[41:0];
  _RAND_23 = {2{`RANDOM}};
  cache_tag_23 = _RAND_23[41:0];
  _RAND_24 = {2{`RANDOM}};
  cache_tag_24 = _RAND_24[41:0];
  _RAND_25 = {2{`RANDOM}};
  cache_tag_25 = _RAND_25[41:0];
  _RAND_26 = {2{`RANDOM}};
  cache_tag_26 = _RAND_26[41:0];
  _RAND_27 = {2{`RANDOM}};
  cache_tag_27 = _RAND_27[41:0];
  _RAND_28 = {2{`RANDOM}};
  cache_tag_28 = _RAND_28[41:0];
  _RAND_29 = {2{`RANDOM}};
  cache_tag_29 = _RAND_29[41:0];
  _RAND_30 = {2{`RANDOM}};
  cache_tag_30 = _RAND_30[41:0];
  _RAND_31 = {2{`RANDOM}};
  cache_tag_31 = _RAND_31[41:0];
  _RAND_32 = {2{`RANDOM}};
  cache_tag_32 = _RAND_32[41:0];
  _RAND_33 = {2{`RANDOM}};
  cache_tag_33 = _RAND_33[41:0];
  _RAND_34 = {2{`RANDOM}};
  cache_tag_34 = _RAND_34[41:0];
  _RAND_35 = {2{`RANDOM}};
  cache_tag_35 = _RAND_35[41:0];
  _RAND_36 = {2{`RANDOM}};
  cache_tag_36 = _RAND_36[41:0];
  _RAND_37 = {2{`RANDOM}};
  cache_tag_37 = _RAND_37[41:0];
  _RAND_38 = {2{`RANDOM}};
  cache_tag_38 = _RAND_38[41:0];
  _RAND_39 = {2{`RANDOM}};
  cache_tag_39 = _RAND_39[41:0];
  _RAND_40 = {2{`RANDOM}};
  cache_tag_40 = _RAND_40[41:0];
  _RAND_41 = {2{`RANDOM}};
  cache_tag_41 = _RAND_41[41:0];
  _RAND_42 = {2{`RANDOM}};
  cache_tag_42 = _RAND_42[41:0];
  _RAND_43 = {2{`RANDOM}};
  cache_tag_43 = _RAND_43[41:0];
  _RAND_44 = {2{`RANDOM}};
  cache_tag_44 = _RAND_44[41:0];
  _RAND_45 = {2{`RANDOM}};
  cache_tag_45 = _RAND_45[41:0];
  _RAND_46 = {2{`RANDOM}};
  cache_tag_46 = _RAND_46[41:0];
  _RAND_47 = {2{`RANDOM}};
  cache_tag_47 = _RAND_47[41:0];
  _RAND_48 = {2{`RANDOM}};
  cache_tag_48 = _RAND_48[41:0];
  _RAND_49 = {2{`RANDOM}};
  cache_tag_49 = _RAND_49[41:0];
  _RAND_50 = {2{`RANDOM}};
  cache_tag_50 = _RAND_50[41:0];
  _RAND_51 = {2{`RANDOM}};
  cache_tag_51 = _RAND_51[41:0];
  _RAND_52 = {2{`RANDOM}};
  cache_tag_52 = _RAND_52[41:0];
  _RAND_53 = {2{`RANDOM}};
  cache_tag_53 = _RAND_53[41:0];
  _RAND_54 = {2{`RANDOM}};
  cache_tag_54 = _RAND_54[41:0];
  _RAND_55 = {2{`RANDOM}};
  cache_tag_55 = _RAND_55[41:0];
  _RAND_56 = {2{`RANDOM}};
  cache_tag_56 = _RAND_56[41:0];
  _RAND_57 = {2{`RANDOM}};
  cache_tag_57 = _RAND_57[41:0];
  _RAND_58 = {2{`RANDOM}};
  cache_tag_58 = _RAND_58[41:0];
  _RAND_59 = {2{`RANDOM}};
  cache_tag_59 = _RAND_59[41:0];
  _RAND_60 = {2{`RANDOM}};
  cache_tag_60 = _RAND_60[41:0];
  _RAND_61 = {2{`RANDOM}};
  cache_tag_61 = _RAND_61[41:0];
  _RAND_62 = {2{`RANDOM}};
  cache_tag_62 = _RAND_62[41:0];
  _RAND_63 = {2{`RANDOM}};
  cache_tag_63 = _RAND_63[41:0];
  _RAND_64 = {2{`RANDOM}};
  cache_tag_64 = _RAND_64[41:0];
  _RAND_65 = {2{`RANDOM}};
  cache_tag_65 = _RAND_65[41:0];
  _RAND_66 = {2{`RANDOM}};
  cache_tag_66 = _RAND_66[41:0];
  _RAND_67 = {2{`RANDOM}};
  cache_tag_67 = _RAND_67[41:0];
  _RAND_68 = {2{`RANDOM}};
  cache_tag_68 = _RAND_68[41:0];
  _RAND_69 = {2{`RANDOM}};
  cache_tag_69 = _RAND_69[41:0];
  _RAND_70 = {2{`RANDOM}};
  cache_tag_70 = _RAND_70[41:0];
  _RAND_71 = {2{`RANDOM}};
  cache_tag_71 = _RAND_71[41:0];
  _RAND_72 = {2{`RANDOM}};
  cache_tag_72 = _RAND_72[41:0];
  _RAND_73 = {2{`RANDOM}};
  cache_tag_73 = _RAND_73[41:0];
  _RAND_74 = {2{`RANDOM}};
  cache_tag_74 = _RAND_74[41:0];
  _RAND_75 = {2{`RANDOM}};
  cache_tag_75 = _RAND_75[41:0];
  _RAND_76 = {2{`RANDOM}};
  cache_tag_76 = _RAND_76[41:0];
  _RAND_77 = {2{`RANDOM}};
  cache_tag_77 = _RAND_77[41:0];
  _RAND_78 = {2{`RANDOM}};
  cache_tag_78 = _RAND_78[41:0];
  _RAND_79 = {2{`RANDOM}};
  cache_tag_79 = _RAND_79[41:0];
  _RAND_80 = {2{`RANDOM}};
  cache_tag_80 = _RAND_80[41:0];
  _RAND_81 = {2{`RANDOM}};
  cache_tag_81 = _RAND_81[41:0];
  _RAND_82 = {2{`RANDOM}};
  cache_tag_82 = _RAND_82[41:0];
  _RAND_83 = {2{`RANDOM}};
  cache_tag_83 = _RAND_83[41:0];
  _RAND_84 = {2{`RANDOM}};
  cache_tag_84 = _RAND_84[41:0];
  _RAND_85 = {2{`RANDOM}};
  cache_tag_85 = _RAND_85[41:0];
  _RAND_86 = {2{`RANDOM}};
  cache_tag_86 = _RAND_86[41:0];
  _RAND_87 = {2{`RANDOM}};
  cache_tag_87 = _RAND_87[41:0];
  _RAND_88 = {2{`RANDOM}};
  cache_tag_88 = _RAND_88[41:0];
  _RAND_89 = {2{`RANDOM}};
  cache_tag_89 = _RAND_89[41:0];
  _RAND_90 = {2{`RANDOM}};
  cache_tag_90 = _RAND_90[41:0];
  _RAND_91 = {2{`RANDOM}};
  cache_tag_91 = _RAND_91[41:0];
  _RAND_92 = {2{`RANDOM}};
  cache_tag_92 = _RAND_92[41:0];
  _RAND_93 = {2{`RANDOM}};
  cache_tag_93 = _RAND_93[41:0];
  _RAND_94 = {2{`RANDOM}};
  cache_tag_94 = _RAND_94[41:0];
  _RAND_95 = {2{`RANDOM}};
  cache_tag_95 = _RAND_95[41:0];
  _RAND_96 = {2{`RANDOM}};
  cache_tag_96 = _RAND_96[41:0];
  _RAND_97 = {2{`RANDOM}};
  cache_tag_97 = _RAND_97[41:0];
  _RAND_98 = {2{`RANDOM}};
  cache_tag_98 = _RAND_98[41:0];
  _RAND_99 = {2{`RANDOM}};
  cache_tag_99 = _RAND_99[41:0];
  _RAND_100 = {2{`RANDOM}};
  cache_tag_100 = _RAND_100[41:0];
  _RAND_101 = {2{`RANDOM}};
  cache_tag_101 = _RAND_101[41:0];
  _RAND_102 = {2{`RANDOM}};
  cache_tag_102 = _RAND_102[41:0];
  _RAND_103 = {2{`RANDOM}};
  cache_tag_103 = _RAND_103[41:0];
  _RAND_104 = {2{`RANDOM}};
  cache_tag_104 = _RAND_104[41:0];
  _RAND_105 = {2{`RANDOM}};
  cache_tag_105 = _RAND_105[41:0];
  _RAND_106 = {2{`RANDOM}};
  cache_tag_106 = _RAND_106[41:0];
  _RAND_107 = {2{`RANDOM}};
  cache_tag_107 = _RAND_107[41:0];
  _RAND_108 = {2{`RANDOM}};
  cache_tag_108 = _RAND_108[41:0];
  _RAND_109 = {2{`RANDOM}};
  cache_tag_109 = _RAND_109[41:0];
  _RAND_110 = {2{`RANDOM}};
  cache_tag_110 = _RAND_110[41:0];
  _RAND_111 = {2{`RANDOM}};
  cache_tag_111 = _RAND_111[41:0];
  _RAND_112 = {2{`RANDOM}};
  cache_tag_112 = _RAND_112[41:0];
  _RAND_113 = {2{`RANDOM}};
  cache_tag_113 = _RAND_113[41:0];
  _RAND_114 = {2{`RANDOM}};
  cache_tag_114 = _RAND_114[41:0];
  _RAND_115 = {2{`RANDOM}};
  cache_tag_115 = _RAND_115[41:0];
  _RAND_116 = {2{`RANDOM}};
  cache_tag_116 = _RAND_116[41:0];
  _RAND_117 = {2{`RANDOM}};
  cache_tag_117 = _RAND_117[41:0];
  _RAND_118 = {2{`RANDOM}};
  cache_tag_118 = _RAND_118[41:0];
  _RAND_119 = {2{`RANDOM}};
  cache_tag_119 = _RAND_119[41:0];
  _RAND_120 = {2{`RANDOM}};
  cache_tag_120 = _RAND_120[41:0];
  _RAND_121 = {2{`RANDOM}};
  cache_tag_121 = _RAND_121[41:0];
  _RAND_122 = {2{`RANDOM}};
  cache_tag_122 = _RAND_122[41:0];
  _RAND_123 = {2{`RANDOM}};
  cache_tag_123 = _RAND_123[41:0];
  _RAND_124 = {2{`RANDOM}};
  cache_tag_124 = _RAND_124[41:0];
  _RAND_125 = {2{`RANDOM}};
  cache_tag_125 = _RAND_125[41:0];
  _RAND_126 = {2{`RANDOM}};
  cache_tag_126 = _RAND_126[41:0];
  _RAND_127 = {2{`RANDOM}};
  cache_tag_127 = _RAND_127[41:0];
  _RAND_128 = {1{`RANDOM}};
  valid_0_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_0_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_1_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_1_1 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_2_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_2_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_3_0 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_3_1 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_4_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_4_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_5_0 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_5_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_6_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_6_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_7_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_7_1 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_8_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_8_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_9_0 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_9_1 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_10_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_10_1 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_11_0 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_11_1 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_12_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_12_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_13_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_13_1 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_14_0 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_14_1 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_15_0 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_15_1 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_16_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_16_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_17_0 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_17_1 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_18_0 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_18_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_19_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_19_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_20_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_20_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_21_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_21_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_22_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_22_1 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_23_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_23_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_24_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_24_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_25_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_25_1 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_26_0 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_26_1 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_27_0 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_27_1 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_28_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_28_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_29_0 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_29_1 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_30_0 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_30_1 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_31_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_31_1 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_32_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_32_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_33_0 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_33_1 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_34_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_34_1 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_35_0 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_35_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_36_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_36_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_37_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_37_1 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_38_0 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_38_1 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_39_0 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_39_1 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_40_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_40_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_41_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_41_1 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_42_0 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_42_1 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_43_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_43_1 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_44_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_44_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_45_0 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_45_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_46_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_46_1 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_47_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_47_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_48_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_48_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_49_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_49_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_50_0 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_50_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_51_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_51_1 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_52_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_52_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_53_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_53_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_54_0 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_54_1 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_55_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_55_1 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_56_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_56_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_57_0 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_57_1 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_58_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_58_1 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_59_0 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_59_1 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_60_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_60_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_61_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_61_1 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_62_0 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_62_1 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_63_0 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_63_1 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_64_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_64_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_65_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_65_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_66_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_66_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_67_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_67_1 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_68_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_68_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_69_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_69_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_70_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_70_1 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_71_0 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_71_1 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_72_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_72_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_73_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_73_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_74_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_74_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_75_0 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_75_1 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_76_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_76_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_77_0 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_77_1 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_78_0 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_78_1 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_79_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_79_1 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_80_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_80_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_81_0 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_81_1 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_82_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_82_1 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_83_0 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_83_1 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_84_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_84_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_85_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_85_1 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_86_0 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_86_1 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_87_0 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_87_1 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_88_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_88_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_89_0 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_89_1 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_90_0 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_90_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_91_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_91_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_92_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_92_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_93_0 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_93_1 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_94_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_94_1 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_95_0 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_95_1 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_96_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_96_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_97_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_97_1 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_98_0 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_98_1 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_99_0 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_99_1 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_100_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_100_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_101_0 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_101_1 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_102_0 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_102_1 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_103_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_103_1 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_104_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_104_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_105_0 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_105_1 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_106_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_106_1 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_107_0 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_107_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_108_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_108_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_109_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_109_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_110_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_110_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_111_0 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_111_1 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_112_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_112_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_113_0 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_113_1 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_114_0 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_114_1 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_115_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_115_1 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_116_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_116_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_117_0 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_117_1 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_118_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_118_1 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_119_0 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_119_1 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_120_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_120_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_121_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_121_1 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_122_0 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_122_1 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_123_0 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_123_1 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_124_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_124_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_125_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_125_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_126_0 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_126_1 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_127_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_127_1 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  state = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  addr = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  uncache = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  cnt = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  flag = _RAND_389[0:0];
  _RAND_390 = {2{`RANDOM}};
  rdata = _RAND_390[63:0];
  _RAND_391 = {1{`RANDOM}};
  hit_num = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  inst_num = _RAND_392[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
