/* verilator lint_off WIDTH */
module AXI4SRAM(
  input         clock,
  input         reset,
  output        io_ar_ready,
  input         io_ar_valid,
  input  [31:0] io_ar_bits_addr,
  input  [7:0]  io_ar_bits_len,
  input  [2:0]  io_ar_bits_size,
  input         io_r_ready,
  output        io_r_valid,
  output [63:0] io_r_bits_data,
  output        io_aw_ready,
  input         io_aw_valid,
  input  [31:0] io_aw_bits_addr,
  input  [2:0]  io_aw_bits_size,
  output        io_w_ready,
  input         io_w_valid,
  input  [63:0] io_w_bits_data,
  input  [7:0]  io_w_bits_strb,
  input         io_w_bits_last,
  output        io_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] pmem_raddr; // @[SRAM.scala 134:19]
  wire [63:0] pmem_rdata; // @[SRAM.scala 134:19]
  wire [31:0] pmem_waddr; // @[SRAM.scala 134:19]
  wire [63:0] pmem_wdata; // @[SRAM.scala 134:19]
  wire [7:0] pmem_wmask; // @[SRAM.scala 134:19]
  reg  rstate; // @[SRAM.scala 78:23]
  wire  _rstate_T = io_ar_ready & io_ar_valid; // @[Decoupled.scala 52:35]
  reg [7:0] rcnt; // @[SRAM.scala 96:21]
  reg [7:0] rlen; // @[SRAM.scala 92:19]
  wire  _rlast_T_1 = io_r_ready & io_r_valid; // @[Decoupled.scala 52:35]
  wire  rlast = rcnt == rlen & _rlast_T_1; // @[SRAM.scala 115:25]
  reg  wstate; // @[SRAM.scala 84:23]
  wire  _wstate_T = io_aw_ready & io_aw_valid; // @[Decoupled.scala 52:35]
  reg [31:0] raddr; // @[SRAM.scala 91:20]
  reg [2:0] rsize; // @[SRAM.scala 93:20]
  reg [31:0] lower_bound_addr; // @[SRAM.scala 95:31]
  reg [7:0] beatcnt; // @[SRAM.scala 97:24]
  wire [31:0] _lower_bound_addr_WIRE = {{24'd0}, io_ar_bits_len}; // @[SRAM.scala 100:{81,81}]
  wire [31:0] _lower_bound_addr_T_1 = ~_lower_bound_addr_WIRE; // @[SRAM.scala 100:57]
  wire [38:0] _GEN_2 = {{7'd0}, _lower_bound_addr_T_1}; // @[SRAM.scala 100:95]
  wire [38:0] _lower_bound_addr_T_2 = _GEN_2 << io_ar_bits_size; // @[SRAM.scala 100:95]
  wire [38:0] _GEN_0 = {{7'd0}, io_ar_bits_addr}; // @[SRAM.scala 100:52]
  wire [38:0] _lower_bound_addr_T_3 = _GEN_0 & _lower_bound_addr_T_2; // @[SRAM.scala 100:52]
  wire [38:0] _lower_bound_addr_T_4 = _rstate_T ? _lower_bound_addr_T_3 : {{7'd0}, lower_bound_addr}; // @[SRAM.scala 100:24]
  wire  _raddr_T_7 = beatcnt == 8'hff | beatcnt == rlen; // @[SRAM.scala 104:47]
  wire [38:0] _raddr_T_10 = 39'h1 << rsize; // @[SRAM.scala 105:45]
  wire [38:0] _GEN_1 = {{7'd0}, raddr}; // @[SRAM.scala 105:33]
  wire [38:0] _raddr_T_12 = _GEN_1 + _raddr_T_10; // @[SRAM.scala 105:33]
  wire [38:0] _raddr_T_13 = _rlast_T_1 ? _raddr_T_12 : {{7'd0}, raddr}; // @[SRAM.scala 105:15]
  wire [38:0] _raddr_T_14 = _rlast_T_1 & (beatcnt == 8'hff | beatcnt == rlen) ? {{7'd0}, lower_bound_addr} : _raddr_T_13
    ; // @[SRAM.scala 104:15]
  wire [38:0] _raddr_T_15 = rlast ? 39'h0 : _raddr_T_14; // @[SRAM.scala 103:15]
  wire [38:0] _raddr_T_16 = _rstate_T & ~rstate ? {{7'd0}, io_ar_bits_addr} : _raddr_T_15; // @[SRAM.scala 102:15]
  wire [7:0] _rcnt_T_7 = rcnt + 8'h1; // @[SRAM.scala 110:28]
  wire [31:0] _beatcnt_T_1 = io_ar_bits_addr >> io_ar_bits_size; // @[SRAM.scala 111:44]
  wire [31:0] _beatcnt_T_2 = _beatcnt_T_1 & _lower_bound_addr_WIRE; // @[SRAM.scala 111:64]
  wire [7:0] _beatcnt_T_8 = beatcnt + 8'h1; // @[SRAM.scala 113:41]
  wire [7:0] _beatcnt_T_9 = rstate ? _beatcnt_T_8 : 8'h0; // @[SRAM.scala 113:15]
  wire [7:0] _beatcnt_T_10 = _raddr_T_7 ? 8'h0 : _beatcnt_T_9; // @[SRAM.scala 112:15]
  wire [31:0] _beatcnt_T_11 = _rstate_T ? _beatcnt_T_2 : {{24'd0}, _beatcnt_T_10}; // @[SRAM.scala 111:15]
  reg [31:0] waddr; // @[SRAM.scala 121:22]
  reg [2:0] wsize; // @[SRAM.scala 124:22]
  wire  _waddr_T_4 = io_w_ready & io_w_valid; // @[Decoupled.scala 52:35]
  wire [38:0] _waddr_T_5 = 39'h1 << wsize; // @[SRAM.scala 130:41]
  wire [38:0] _GEN_3 = {{7'd0}, waddr}; // @[SRAM.scala 130:30]
  wire [38:0] _waddr_T_7 = _GEN_3 + _waddr_T_5; // @[SRAM.scala 130:30]
  wire [38:0] _waddr_T_8 = _waddr_T_4 ? _waddr_T_7 : {{7'd0}, waddr}; // @[SRAM.scala 130:13]
  wire [38:0] _waddr_T_9 = io_w_bits_last ? 39'h0 : _waddr_T_8; // @[SRAM.scala 129:13]
  wire [38:0] _waddr_T_10 = _wstate_T & ~wstate ? {{7'd0}, io_aw_bits_addr} : _waddr_T_9; // @[SRAM.scala 128:13]
  reg  b; // @[SRAM.scala 148:16]
  wire [7:0] _T_1 = rlen + 8'h1; // @[SRAM.scala 156:45]
  wire [7:0] _T_2 = 8'h1 << rsize; // @[SRAM.scala 156:55]
  wire [15:0] _T_3 = _T_1 * _T_2; // @[SRAM.scala 156:50]
  wire [31:0] _GEN_4 = {{16'd0}, _T_3}; // @[SRAM.scala 156:38]
  wire [31:0] _T_5 = lower_bound_addr + _GEN_4; // @[SRAM.scala 156:38]
  wire [38:0] _GEN_5 = reset ? 39'h0 : _raddr_T_16; // @[SRAM.scala 91:{20,20} 102:9]
  wire [38:0] _GEN_6 = reset ? 39'h0 : _lower_bound_addr_T_4; // @[SRAM.scala 100:19 95:{31,31}]
  wire [31:0] _GEN_7 = reset ? 32'h0 : _beatcnt_T_11; // @[SRAM.scala 111:10 97:{24,24}]
  wire [38:0] _GEN_8 = reset ? 39'h0 : _waddr_T_10; // @[SRAM.scala 121:{22,22} 128:8]
  memory pmem ( // @[SRAM.scala 134:19]
    .raddr(pmem_raddr),
    .rdata(pmem_rdata),
    .waddr(pmem_waddr),
    .wdata(pmem_wdata),
    .wmask(pmem_wmask)
  );
  assign io_ar_ready = ~rstate; // @[SRAM.scala 140:26]
  assign io_r_valid = rstate; // @[SRAM.scala 141:26]
  assign io_r_bits_data = pmem_rdata; // @[SRAM.scala 145:18]
  assign io_aw_ready = ~wstate; // @[SRAM.scala 143:26]
  assign io_w_ready = wstate; // @[SRAM.scala 144:26]
  assign io_b_valid = b; // @[SRAM.scala 150:14]
  assign pmem_raddr = raddr; // @[SRAM.scala 135:16]
  assign pmem_waddr = waddr; // @[SRAM.scala 136:16]
  assign pmem_wdata = io_w_bits_data; // @[SRAM.scala 137:16]
  assign pmem_wmask = _waddr_T_4 ? io_w_bits_strb : 8'h0; // @[SRAM.scala 138:22]
  always @(posedge clock) begin
    if (reset) begin // @[SRAM.scala 78:23]
      rstate <= 1'h0; // @[SRAM.scala 78:23]
    end else if (rstate) begin // @[Mux.scala 81:58]
      if (rlast) begin // @[SRAM.scala 82:25]
        rstate <= 1'h0;
      end else begin
        rstate <= 1'h1;
      end
    end else begin
      rstate <= _rstate_T;
    end
    if (reset) begin // @[SRAM.scala 96:21]
      rcnt <= 8'h0; // @[SRAM.scala 96:21]
    end else if (rcnt == 8'hff | rlast | _rstate_T) begin // @[SRAM.scala 109:12]
      rcnt <= 8'h0;
    end else if (_rlast_T_1) begin // @[SRAM.scala 110:12]
      rcnt <= _rcnt_T_7;
    end
    if (reset) begin // @[SRAM.scala 92:19]
      rlen <= 8'h0; // @[SRAM.scala 92:19]
    end else if (_rstate_T) begin // @[SRAM.scala 106:14]
      rlen <= io_ar_bits_len;
    end
    if (reset) begin // @[SRAM.scala 84:23]
      wstate <= 1'h0; // @[SRAM.scala 84:23]
    end else if (wstate) begin // @[Mux.scala 81:58]
      if (io_w_bits_last) begin // @[SRAM.scala 87:25]
        wstate <= 1'h0;
      end else begin
        wstate <= 1'h1;
      end
    end else begin
      wstate <= _wstate_T;
    end
    raddr <= _GEN_5[31:0]; // @[SRAM.scala 91:{20,20} 102:9]
    if (reset) begin // @[SRAM.scala 93:20]
      rsize <= 3'h0; // @[SRAM.scala 93:20]
    end else if (_rstate_T) begin // @[SRAM.scala 107:15]
      rsize <= io_ar_bits_size;
    end
    lower_bound_addr <= _GEN_6[31:0]; // @[SRAM.scala 100:19 95:{31,31}]
    beatcnt <= _GEN_7[7:0]; // @[SRAM.scala 111:10 97:{24,24}]
    waddr <= _GEN_8[31:0]; // @[SRAM.scala 121:{22,22} 128:8]
    if (reset) begin // @[SRAM.scala 124:22]
      wsize <= 3'h0; // @[SRAM.scala 124:22]
    end else if (_wstate_T) begin // @[SRAM.scala 127:13]
      wsize <= io_aw_bits_size;
    end
    if (reset) begin // @[SRAM.scala 148:16]
      b <= 1'h0; // @[SRAM.scala 148:16]
    end else begin
      b <= io_w_bits_last; // @[SRAM.scala 149:4]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(raddr < _T_5 & raddr >= lower_bound_addr | raddr == 32'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SRAM.scala:156 assert(((raddr <  lower_bound_addr + (rlen+1.U)*(1.U<<rsize )) && (raddr >= lower_bound_addr)) || (raddr === 0.U))\n"
            ); // @[SRAM.scala 156:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(raddr < _T_5 & raddr >= lower_bound_addr | raddr == 32'h0)) begin
          $fatal; // @[SRAM.scala 156:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rstate = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rcnt = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  rlen = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  wstate = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  raddr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rsize = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  lower_bound_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  beatcnt = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  waddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  wsize = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  b = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pre_Decode(
  input  [31:0] io_inst,
  output        io_jump
);
  wire  _io_jump_T_5 = io_inst[14:12] == 3'h0; // @[IFU.scala 83:51]
  wire  _io_jump_T_6 = io_inst[6:0] == 7'h67 & io_inst[14:12] == 3'h0; // @[IFU.scala 83:38]
  wire  _io_jump_T_7 = io_inst[6:0] == 7'h6f | _io_jump_T_6; // @[IFU.scala 82:64]
  wire  _io_jump_T_9 = io_inst[6:0] == 7'h63; // @[IFU.scala 84:22]
  wire  _io_jump_T_12 = io_inst[6:0] == 7'h63 & _io_jump_T_5; // @[IFU.scala 84:38]
  wire  _io_jump_T_13 = _io_jump_T_7 | _io_jump_T_12; // @[IFU.scala 83:64]
  wire  _io_jump_T_18 = _io_jump_T_9 & io_inst[14:12] == 3'h1; // @[IFU.scala 85:38]
  wire  _io_jump_T_19 = _io_jump_T_13 | _io_jump_T_18; // @[IFU.scala 84:64]
  wire  _io_jump_T_24 = _io_jump_T_9 & io_inst[14:12] == 3'h5; // @[IFU.scala 86:38]
  wire  _io_jump_T_25 = _io_jump_T_19 | _io_jump_T_24; // @[IFU.scala 85:64]
  wire  _io_jump_T_30 = _io_jump_T_9 & io_inst[14:12] == 3'h7; // @[IFU.scala 87:38]
  wire  _io_jump_T_31 = _io_jump_T_25 | _io_jump_T_30; // @[IFU.scala 86:64]
  wire  _io_jump_T_36 = _io_jump_T_9 & io_inst[14:12] == 3'h4; // @[IFU.scala 88:38]
  wire  _io_jump_T_37 = _io_jump_T_31 | _io_jump_T_36; // @[IFU.scala 87:64]
  wire  _io_jump_T_42 = _io_jump_T_9 & io_inst[14:12] == 3'h6; // @[IFU.scala 89:38]
  wire  _io_jump_T_43 = _io_jump_T_37 | _io_jump_T_42; // @[IFU.scala 88:64]
  wire  _io_jump_T_44 = io_inst == 32'h73; // @[IFU.scala 90:17]
  wire  _io_jump_T_45 = _io_jump_T_43 | _io_jump_T_44; // @[IFU.scala 89:64]
  wire  _io_jump_T_46 = io_inst == 32'h30200073; // @[IFU.scala 91:17]
  wire  _io_jump_T_47 = _io_jump_T_45 | _io_jump_T_46; // @[IFU.scala 90:64]
  wire  _io_jump_T_48 = io_inst == 32'h100073; // @[IFU.scala 92:17]
  assign io_jump = _io_jump_T_47 | _io_jump_T_48; // @[IFU.scala 91:64]
endmodule
module IFU(
  input         clock,
  input         reset,
  input  [63:0] io_pc_dnpc,
  input         io_clearJump,
  input         io_lm_ar_ready,
  output        io_lm_ar_valid,
  output [31:0] io_lm_ar_bits_addr,
  output        io_lm_r_ready,
  input         io_lm_r_valid,
  input  [63:0] io_lm_r_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_pc,
  output [31:0] io_out_bits_inst,
  output        io_out_bits_isJump
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] pre_decode_io_inst; // @[IFU.scala 37:25]
  wire  pre_decode_io_jump; // @[IFU.scala 37:25]
  wire [63:0] it_pc; // @[IFU.scala 68:16]
  wire  it_en; // @[IFU.scala 68:16]
  wire [31:0] it_inst; // @[IFU.scala 68:16]
  reg [1:0] state; // @[IFU.scala 29:22]
  wire  _state_T = io_lm_ar_ready & io_lm_ar_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _state_T_1 = _state_T ? 2'h1 : 2'h0; // @[IFU.scala 31:25]
  wire  _state_T_2 = io_lm_r_ready & io_lm_r_valid; // @[Decoupled.scala 52:35]
  wire  _state_T_4 = io_out_ready & io_out_valid; // @[Decoupled.scala 52:35]
  reg [31:0] IF_reg_inst; // @[Reg.scala 35:20]
  reg  IF_reg_valid; // @[Reg.scala 35:20]
  wire  _next_valid_T_4 = pre_decode_io_jump & _state_T_4 ? 1'h0 : IF_reg_valid; // @[IFU.scala 45:18]
  wire  next_valid = io_clearJump | _next_valid_T_4; // @[IFU.scala 44:18]
  reg [63:0] IF_reg_pc; // @[Reg.scala 35:20]
  wire [63:0] _next_pc_T_3 = IF_reg_pc + 64'h4; // @[IFU.scala 49:38]
  Pre_Decode pre_decode ( // @[IFU.scala 37:25]
    .io_inst(pre_decode_io_inst),
    .io_jump(pre_decode_io_jump)
  );
  itrace it ( // @[IFU.scala 68:16]
    .pc(it_pc),
    .en(it_en),
    .inst(it_inst)
  );
  assign io_lm_ar_valid = state == 2'h0 & ~reset & IF_reg_valid; // @[IFU.scala 53:53]
  assign io_lm_ar_bits_addr = IF_reg_pc[31:0]; // @[IFU.scala 52:32]
  assign io_lm_r_ready = 1'h1; // @[IFU.scala 54:16]
  assign io_out_valid = state == 2'h2; // @[IFU.scala 66:26]
  assign io_out_bits_pc = IF_reg_pc[31:0]; // @[IFU.scala 64:28]
  assign io_out_bits_inst = IF_reg_inst; // @[IFU.scala 63:19]
  assign io_out_bits_isJump = pre_decode_io_jump; // @[IFU.scala 65:21]
  assign pre_decode_io_inst = IF_reg_inst; // @[IFU.scala 38:21]
  assign it_pc = {{32'd0}, io_lm_ar_bits_addr}; // @[IFU.scala 71:11]
  assign it_en = io_lm_r_ready & io_lm_r_valid; // @[Decoupled.scala 52:35]
  assign it_inst = io_lm_r_bits_data[31:0]; // @[IFU.scala 70:32]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 29:22]
      state <= 2'h0; // @[IFU.scala 29:22]
    end else if (2'h2 == state) begin // @[Mux.scala 81:58]
      if (_state_T_4) begin // @[IFU.scala 33:25]
        state <= 2'h0;
      end else begin
        state <= 2'h2;
      end
    end else if (2'h1 == state) begin // @[Mux.scala 81:58]
      if (_state_T_2) begin // @[IFU.scala 32:25]
        state <= 2'h2;
      end else begin
        state <= 2'h1;
      end
    end else if (2'h0 == state) begin // @[Mux.scala 81:58]
      state <= _state_T_1;
    end else begin
      state <= 2'h0;
    end
    if (reset) begin // @[Reg.scala 35:20]
      IF_reg_inst <= 32'h0; // @[Reg.scala 35:20]
    end else if (_state_T_2) begin // @[Reg.scala 36:18]
      IF_reg_inst <= io_lm_r_bits_data[31:0]; // @[Reg.scala 36:22]
    end
    IF_reg_valid <= reset | next_valid; // @[Reg.scala 35:{20,20}]
    if (reset) begin // @[Reg.scala 35:20]
      IF_reg_pc <= 64'h80000000; // @[Reg.scala 35:20]
    end else if (next_valid) begin // @[Reg.scala 36:18]
      if (io_clearJump) begin // @[IFU.scala 48:16]
        IF_reg_pc <= io_pc_dnpc;
      end else if (_state_T_4) begin // @[IFU.scala 49:16]
        IF_reg_pc <= _next_pc_T_3;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  IF_reg_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  IF_reg_valid = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  IF_reg_pc = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [31:0] io_in_bits_inst,
  input         io_in_bits_isJump,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_pc,
  output [31:0] io_out_bits_inst,
  output [4:0]  io_out_bits_rs1,
  output [4:0]  io_out_bits_rs2,
  output [4:0]  io_out_bits_rd,
  output [63:0] io_out_bits_imm,
  output [79:0] io_out_bits_op,
  output [5:0]  io_out_bits_typ,
  output        io_out_bits_isJump,
  output [4:0]  io_out_bits_clearidx,
  output [4:0]  io_sb_lookidx1,
  output [4:0]  io_sb_lookidx2,
  output [4:0]  io_sb_setidx,
  input         io_sb_isBusy
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  _ID_reg_inst_T = io_in_ready & io_in_valid; // @[Decoupled.scala 52:35]
  reg [31:0] ID_reg_inst; // @[Reg.scala 35:20]
  reg [31:0] ID_reg_pc; // @[Reg.scala 35:20]
  reg  ID_reg_isJump; // @[Reg.scala 35:20]
  reg  state; // @[IDU.scala 34:23]
  wire  _state_T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 52:35]
  wire  _io_in_ready_T_1 = ~io_sb_isBusy; // @[IDU.scala 41:39]
  wire  _op_t_0_T_1 = ID_reg_inst[6:0] == 7'h33; // @[IDU.scala 50:31]
  wire  _op_t_0_T_3 = ID_reg_inst[14:12] == 3'h0; // @[IDU.scala 50:67]
  wire  _op_t_0_T_4 = ID_reg_inst[6:0] == 7'h33 & ID_reg_inst[14:12] == 3'h0; // @[IDU.scala 50:47]
  wire  _op_t_0_T_6 = ID_reg_inst[31:25] == 7'h0; // @[IDU.scala 50:99]
  wire  op_t_0 = ID_reg_inst[6:0] == 7'h33 & ID_reg_inst[14:12] == 3'h0 & ID_reg_inst[31:25] == 7'h0; // @[IDU.scala 50:79]
  wire  _op_t_1_T_1 = ID_reg_inst[6:0] == 7'h3b; // @[IDU.scala 51:31]
  wire  _op_t_1_T_4 = ID_reg_inst[6:0] == 7'h3b & _op_t_0_T_3; // @[IDU.scala 51:47]
  wire  op_t_1 = ID_reg_inst[6:0] == 7'h3b & _op_t_0_T_3 & _op_t_0_T_6; // @[IDU.scala 51:79]
  wire  _op_t_2_T_1 = ID_reg_inst[6:0] == 7'h13; // @[IDU.scala 52:31]
  wire  op_t_2 = ID_reg_inst[6:0] == 7'h13 & _op_t_0_T_3; // @[IDU.scala 52:47]
  wire  _op_t_3_T_1 = ID_reg_inst[6:0] == 7'h1b; // @[IDU.scala 53:31]
  wire  op_t_3 = ID_reg_inst[6:0] == 7'h1b & _op_t_0_T_3; // @[IDU.scala 53:47]
  wire  _op_t_4_T_6 = ID_reg_inst[31:25] == 7'h20; // @[IDU.scala 54:99]
  wire  op_t_4 = _op_t_0_T_4 & ID_reg_inst[31:25] == 7'h20; // @[IDU.scala 54:79]
  wire  op_t_5 = _op_t_1_T_4 & _op_t_4_T_6; // @[IDU.scala 55:79]
  wire  _op_t_6_T_3 = ID_reg_inst[14:12] == 3'h7; // @[IDU.scala 56:67]
  wire  _op_t_6_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h7; // @[IDU.scala 56:47]
  wire  op_t_6 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h7 & _op_t_0_T_6; // @[IDU.scala 56:79]
  wire  op_t_7 = _op_t_2_T_1 & _op_t_6_T_3; // @[IDU.scala 57:47]
  wire  _op_t_8_T_3 = ID_reg_inst[14:12] == 3'h6; // @[IDU.scala 58:67]
  wire  _op_t_8_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h6; // @[IDU.scala 58:47]
  wire  op_t_8 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h6 & _op_t_0_T_6; // @[IDU.scala 58:79]
  wire  op_t_9 = _op_t_2_T_1 & _op_t_8_T_3; // @[IDU.scala 59:47]
  wire  _op_t_10_T_3 = ID_reg_inst[14:12] == 3'h4; // @[IDU.scala 60:67]
  wire  _op_t_10_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h4; // @[IDU.scala 60:47]
  wire  op_t_10 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h4 & _op_t_0_T_6; // @[IDU.scala 60:79]
  wire  op_t_11 = _op_t_2_T_1 & _op_t_10_T_3; // @[IDU.scala 61:47]
  wire  _op_t_12_T_3 = ID_reg_inst[14:12] == 3'h1; // @[IDU.scala 62:67]
  wire  _op_t_12_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h1; // @[IDU.scala 62:47]
  wire  op_t_12 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h1 & _op_t_0_T_6; // @[IDU.scala 62:79]
  wire  op_t_13 = _op_t_1_T_1 & _op_t_12_T_3 & _op_t_0_T_6; // @[IDU.scala 63:79]
  wire  _op_t_14_T_6 = ID_reg_inst[31:26] == 6'h0; // @[IDU.scala 64:99]
  wire  op_t_14 = _op_t_2_T_1 & _op_t_12_T_3 & ID_reg_inst[31:26] == 6'h0; // @[IDU.scala 64:79]
  wire  op_t_15 = _op_t_3_T_1 & _op_t_12_T_3 & _op_t_14_T_6; // @[IDU.scala 65:79]
  wire  _op_t_16_T_3 = ID_reg_inst[14:12] == 3'h5; // @[IDU.scala 66:67]
  wire  _op_t_16_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h5; // @[IDU.scala 66:47]
  wire  op_t_16 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h5 & _op_t_4_T_6; // @[IDU.scala 66:79]
  wire  _op_t_17_T_4 = _op_t_1_T_1 & _op_t_16_T_3; // @[IDU.scala 67:47]
  wire  op_t_17 = _op_t_1_T_1 & _op_t_16_T_3 & _op_t_4_T_6; // @[IDU.scala 67:79]
  wire  _op_t_18_T_4 = _op_t_2_T_1 & _op_t_16_T_3; // @[IDU.scala 68:47]
  wire  _op_t_18_T_6 = ID_reg_inst[31:26] == 6'h10; // @[IDU.scala 68:99]
  wire  op_t_18 = _op_t_2_T_1 & _op_t_16_T_3 & ID_reg_inst[31:26] == 6'h10; // @[IDU.scala 68:79]
  wire  _op_t_19_T_4 = _op_t_3_T_1 & _op_t_16_T_3; // @[IDU.scala 69:47]
  wire  op_t_19 = _op_t_3_T_1 & _op_t_16_T_3 & _op_t_18_T_6; // @[IDU.scala 69:79]
  wire  op_t_20 = _op_t_16_T_4 & _op_t_0_T_6; // @[IDU.scala 70:79]
  wire  op_t_21 = _op_t_17_T_4 & _op_t_0_T_6; // @[IDU.scala 71:79]
  wire  op_t_22 = _op_t_18_T_4 & _op_t_14_T_6; // @[IDU.scala 72:79]
  wire  op_t_23 = _op_t_19_T_4 & _op_t_14_T_6; // @[IDU.scala 73:79]
  wire  op_t_24 = ID_reg_inst[6:0] == 7'h37; // @[IDU.scala 74:31]
  wire  op_t_25 = ID_reg_inst[6:0] == 7'h17; // @[IDU.scala 75:31]
  wire  _op_t_26_T_3 = ID_reg_inst[14:12] == 3'h2; // @[IDU.scala 76:67]
  wire  _op_t_26_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h2; // @[IDU.scala 76:47]
  wire  op_t_26 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h2 & _op_t_0_T_6; // @[IDU.scala 76:79]
  wire  _op_t_27_T_3 = ID_reg_inst[14:12] == 3'h3; // @[IDU.scala 77:67]
  wire  _op_t_27_T_4 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h3; // @[IDU.scala 77:47]
  wire  op_t_27 = _op_t_0_T_1 & ID_reg_inst[14:12] == 3'h3 & _op_t_0_T_6; // @[IDU.scala 77:79]
  wire  op_t_28 = _op_t_2_T_1 & _op_t_26_T_3; // @[IDU.scala 78:47]
  wire  op_t_29 = _op_t_2_T_1 & _op_t_27_T_3; // @[IDU.scala 79:47]
  wire  _op_t_30_T_1 = ID_reg_inst[6:0] == 7'h63; // @[IDU.scala 80:31]
  wire  op_t_30 = ID_reg_inst[6:0] == 7'h63 & _op_t_0_T_3; // @[IDU.scala 80:47]
  wire  op_t_31 = _op_t_30_T_1 & _op_t_12_T_3; // @[IDU.scala 81:47]
  wire  op_t_32 = _op_t_30_T_1 & _op_t_16_T_3; // @[IDU.scala 82:47]
  wire  op_t_33 = _op_t_30_T_1 & _op_t_6_T_3; // @[IDU.scala 83:47]
  wire  op_t_34 = _op_t_30_T_1 & _op_t_10_T_3; // @[IDU.scala 84:47]
  wire  op_t_35 = _op_t_30_T_1 & _op_t_8_T_3; // @[IDU.scala 85:47]
  wire  op_t_36 = ID_reg_inst[6:0] == 7'h6f; // @[IDU.scala 86:31]
  wire  op_t_37 = ID_reg_inst[6:0] == 7'h67 & _op_t_0_T_3; // @[IDU.scala 87:47]
  wire  _op_t_38_T_1 = ID_reg_inst[6:0] == 7'h3; // @[IDU.scala 88:31]
  wire  op_t_38 = ID_reg_inst[6:0] == 7'h3 & _op_t_0_T_3; // @[IDU.scala 88:47]
  wire  op_t_39 = _op_t_38_T_1 & _op_t_12_T_3; // @[IDU.scala 89:47]
  wire  op_t_40 = _op_t_38_T_1 & _op_t_26_T_3; // @[IDU.scala 90:47]
  wire  op_t_41 = _op_t_38_T_1 & _op_t_27_T_3; // @[IDU.scala 91:47]
  wire  _op_t_42_T_1 = ID_reg_inst[6:0] == 7'h23; // @[IDU.scala 92:31]
  wire  op_t_42 = ID_reg_inst[6:0] == 7'h23 & _op_t_0_T_3; // @[IDU.scala 92:47]
  wire  op_t_43 = _op_t_42_T_1 & _op_t_12_T_3; // @[IDU.scala 93:47]
  wire  op_t_44 = _op_t_42_T_1 & _op_t_26_T_3; // @[IDU.scala 94:47]
  wire  op_t_45 = _op_t_42_T_1 & _op_t_27_T_3; // @[IDU.scala 95:47]
  wire  op_t_46 = _op_t_38_T_1 & _op_t_10_T_3; // @[IDU.scala 96:47]
  wire  op_t_47 = _op_t_38_T_1 & _op_t_16_T_3; // @[IDU.scala 97:47]
  wire  op_t_48 = _op_t_38_T_1 & _op_t_8_T_3; // @[IDU.scala 98:47]
  wire  op_t_49 = ID_reg_inst == 32'h100073; // @[IDU.scala 99:26]
  wire  _op_t_50_T_6 = ID_reg_inst[31:25] == 7'h1; // @[IDU.scala 102:99]
  wire  op_t_50 = _op_t_0_T_4 & ID_reg_inst[31:25] == 7'h1; // @[IDU.scala 102:79]
  wire  op_t_51 = _op_t_1_T_4 & _op_t_50_T_6; // @[IDU.scala 103:79]
  wire  op_t_52 = _op_t_12_T_4 & _op_t_50_T_6; // @[IDU.scala 104:79]
  wire  op_t_53 = _op_t_27_T_4 & _op_t_50_T_6; // @[IDU.scala 105:79]
  wire  op_t_54 = _op_t_26_T_4 & _op_t_50_T_6; // @[IDU.scala 106:79]
  wire  op_t_55 = _op_t_10_T_4 & _op_t_50_T_6; // @[IDU.scala 107:79]
  wire  op_t_56 = _op_t_1_T_1 & _op_t_10_T_3 & _op_t_50_T_6; // @[IDU.scala 108:79]
  wire  op_t_57 = _op_t_16_T_4 & _op_t_50_T_6; // @[IDU.scala 109:79]
  wire  op_t_58 = _op_t_17_T_4 & _op_t_50_T_6; // @[IDU.scala 110:79]
  wire  op_t_59 = _op_t_8_T_4 & _op_t_50_T_6; // @[IDU.scala 111:79]
  wire  op_t_60 = _op_t_1_T_1 & _op_t_8_T_3 & _op_t_50_T_6; // @[IDU.scala 112:79]
  wire  op_t_61 = _op_t_6_T_4 & _op_t_50_T_6; // @[IDU.scala 113:79]
  wire  op_t_62 = _op_t_1_T_1 & _op_t_6_T_3 & _op_t_50_T_6; // @[IDU.scala 114:79]
  wire  _op_t_63_T_1 = ID_reg_inst[6:0] == 7'h73; // @[IDU.scala 117:31]
  wire  op_t_63 = ID_reg_inst[6:0] == 7'h73 & _op_t_12_T_3; // @[IDU.scala 117:47]
  wire  op_t_64 = _op_t_63_T_1 & _op_t_26_T_3; // @[IDU.scala 118:47]
  wire  op_t_65 = ID_reg_inst == 32'h73; // @[IDU.scala 119:26]
  wire  op_t_66 = ID_reg_inst == 32'h30200073; // @[IDU.scala 120:26]
  wire [9:0] op_lo_lo_lo = {op_t_9,op_t_8,op_t_7,op_t_6,op_t_5,op_t_4,op_t_3,op_t_2,op_t_1,op_t_0}; // @[IDU.scala 123:13]
  wire [9:0] op_lo_lo_hi = {op_t_19,op_t_18,op_t_17,op_t_16,op_t_15,op_t_14,op_t_13,op_t_12,op_t_11,op_t_10}; // @[IDU.scala 123:13]
  wire [9:0] op_lo_hi_lo = {op_t_29,op_t_28,op_t_27,op_t_26,op_t_25,op_t_24,op_t_23,op_t_22,op_t_21,op_t_20}; // @[IDU.scala 123:13]
  wire [9:0] op_lo_hi_hi = {op_t_39,op_t_38,op_t_37,op_t_36,op_t_35,op_t_34,op_t_33,op_t_32,op_t_31,op_t_30}; // @[IDU.scala 123:13]
  wire [39:0] op_lo = {op_lo_hi_hi,op_lo_hi_lo,op_lo_lo_hi,op_lo_lo_lo}; // @[IDU.scala 123:13]
  wire [9:0] op_hi_lo_lo = {op_t_49,op_t_48,op_t_47,op_t_46,op_t_45,op_t_44,op_t_43,op_t_42,op_t_41,op_t_40}; // @[IDU.scala 123:13]
  wire [9:0] op_hi_lo_hi = {op_t_59,op_t_58,op_t_57,op_t_56,op_t_55,op_t_54,op_t_53,op_t_52,op_t_51,op_t_50}; // @[IDU.scala 123:13]
  wire [19:0] op_hi_lo = {op_hi_lo_hi,op_hi_lo_lo}; // @[IDU.scala 123:13]
  wire [39:0] op_hi = {10'h0,3'h0,op_t_66,op_t_65,op_t_64,op_t_63,op_t_62,op_t_61,op_t_60,op_hi_lo}; // @[IDU.scala 123:13]
  wire [79:0] op = {op_hi,op_lo_hi_hi,op_lo_hi_lo,op_lo_lo_hi,op_lo_lo_lo}; // @[IDU.scala 123:13]
  wire  _typ_t_0_T_30 = op[2] | op[3] | op[7] | op[9] | op[11] | op[14] | op[15] | op[18] | op[19] | op[22] | op[23] |
    op[28] | op[29] | op[37] | op[38] | op[39]; // @[IDU.scala 137:116]
  wire  typ_t_0 = _typ_t_0_T_30 | op[40] | op[41] | op[46] | op[47] | op[48] | op[63] | op[64]; // @[IDU.scala 137:165]
  wire  typ_t_1 = op[24] | op[25]; // @[IDU.scala 138:22]
  wire  typ_t_2 = op[42] | op[43] | op[44] | op[45]; // @[IDU.scala 139:36]
  wire  typ_t_3 = op[36]; // @[IDU.scala 140:18]
  wire  typ_t_4 = op[30] | op[31] | op[32] | op[33] | op[34] | op[35]; // @[IDU.scala 141:50]
  wire  _typ_t_5_T_30 = op[0] | op[1] | op[4] | op[5] | op[6] | op[8] | op[10] | op[12] | op[13] | op[16] | op[17] | op[
    20] | op[21] | op[26] | op[27] | op[50]; // @[IDU.scala 142:114]
  wire  typ_t_5 = _typ_t_5_T_30 | op[51] | op[52] | op[53] | op[54] | op[55] | op[56] | op[57] | op[58] | op[59] | op[60
    ] | op[61] | op[62]; // @[IDU.scala 142:198]
  wire [2:0] typ_lo = {typ_t_2,typ_t_1,typ_t_0}; // @[IDU.scala 144:15]
  wire [2:0] typ_hi = {typ_t_5,typ_t_4,typ_t_3}; // @[IDU.scala 144:15]
  wire [5:0] typ = {typ_t_5,typ_t_4,typ_t_3,typ_t_2,typ_t_1,typ_t_0}; // @[IDU.scala 144:15]
  wire [51:0] _io_out_bits_imm_T_3 = ID_reg_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_imm_T_5 = {_io_out_bits_imm_T_3,ID_reg_inst[31:20]}; // @[Cat.scala 33:92]
  wire [31:0] _io_out_bits_imm_T_9 = ID_reg_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_imm_T_13 = {_io_out_bits_imm_T_9,ID_reg_inst[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_imm_T_21 = {_io_out_bits_imm_T_3,ID_reg_inst[31:25],ID_reg_inst[11:7]}; // @[Cat.scala 33:92]
  wire [42:0] _io_out_bits_imm_T_25 = ID_reg_inst[31] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_imm_T_34 = {_io_out_bits_imm_T_25,ID_reg_inst[31],ID_reg_inst[19:12],ID_reg_inst[20],
    ID_reg_inst[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [50:0] _io_out_bits_imm_T_38 = ID_reg_inst[31] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_imm_T_47 = {_io_out_bits_imm_T_38,ID_reg_inst[31],ID_reg_inst[7],ID_reg_inst[30:25],
    ID_reg_inst[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_imm_T_48 = typ[4] ? _io_out_bits_imm_T_47 : 64'h0; // @[IDU.scala 153:25]
  wire [63:0] _io_out_bits_imm_T_49 = typ[3] ? _io_out_bits_imm_T_34 : _io_out_bits_imm_T_48; // @[IDU.scala 152:25]
  wire [63:0] _io_out_bits_imm_T_50 = typ[2] ? _io_out_bits_imm_T_21 : _io_out_bits_imm_T_49; // @[IDU.scala 151:25]
  wire [63:0] _io_out_bits_imm_T_51 = typ[1] ? _io_out_bits_imm_T_13 : _io_out_bits_imm_T_50; // @[IDU.scala 150:25]
  assign io_in_ready = ~state & ~io_sb_isBusy; // @[IDU.scala 41:36]
  assign io_out_valid = state & _io_in_ready_T_1; // @[IDU.scala 42:43]
  assign io_out_bits_pc = ID_reg_pc; // @[IDU.scala 43:18]
  assign io_out_bits_inst = ID_reg_inst; // @[IDU.scala 44:20]
  assign io_out_bits_rs1 = ID_reg_inst[19:15]; // @[IDU.scala 127:32]
  assign io_out_bits_rs2 = ID_reg_inst[24:20]; // @[IDU.scala 128:32]
  assign io_out_bits_rd = ID_reg_inst[11:7]; // @[IDU.scala 126:31]
  assign io_out_bits_imm = typ[0] ? _io_out_bits_imm_T_5 : _io_out_bits_imm_T_51; // @[IDU.scala 149:25]
  assign io_out_bits_op = {op_hi,op_lo}; // @[IDU.scala 123:13]
  assign io_out_bits_typ = {typ_hi,typ_lo}; // @[IDU.scala 144:15]
  assign io_out_bits_isJump = ID_reg_isJump; // @[IDU.scala 29:22]
  assign io_out_bits_clearidx = io_sb_setidx; // @[IDU.scala 160:24]
  assign io_sb_lookidx1 = typ[0] | typ[2] | typ[4] | typ[5] ? ID_reg_inst[19:15] : 5'h0; // @[IDU.scala 157:23]
  assign io_sb_lookidx2 = typ[2] | typ[4] | typ[5] ? ID_reg_inst[24:20] : 5'h0; // @[IDU.scala 158:23]
  assign io_sb_setidx = (typ[0] | typ[1] | typ[3] | typ[5]) & _state_T_2 ? ID_reg_inst[11:7] : 5'h0; // @[IDU.scala 159:21]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      ID_reg_inst <= 32'h0; // @[Reg.scala 35:20]
    end else if (_ID_reg_inst_T) begin // @[Reg.scala 36:18]
      ID_reg_inst <= io_in_bits_inst; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ID_reg_pc <= 32'h0; // @[Reg.scala 35:20]
    end else if (_ID_reg_inst_T) begin // @[Reg.scala 36:18]
      ID_reg_pc <= io_in_bits_pc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ID_reg_isJump <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ID_reg_inst_T) begin // @[Reg.scala 36:18]
      ID_reg_isJump <= io_in_bits_isJump; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[IDU.scala 34:23]
      state <= 1'h0; // @[IDU.scala 34:23]
    end else if (state) begin // @[Mux.scala 81:58]
      if (_state_T_2) begin // @[IDU.scala 39:25]
        state <= 1'h0;
      end else begin
        state <= 1'h1;
      end
    end else begin
      state <= _ID_reg_inst_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID_reg_inst = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ID_reg_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ID_reg_isJump = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_ls_in_valid,
  input  [31:0] io_ls_in_bits_raddr,
  input  [31:0] io_ls_in_bits_waddr,
  input  [63:0] io_ls_in_bits_wdata,
  input  [7:0]  io_ls_in_bits_wmask,
  input         io_ls_out_ready,
  output        io_ls_out_valid,
  output [63:0] io_ls_out_bits_rdata,
  input         io_en_r,
  input         io_en_w,
  input         io_lm_ar_ready,
  output        io_lm_ar_valid,
  output [31:0] io_lm_ar_bits_addr,
  output        io_lm_r_ready,
  input         io_lm_r_valid,
  input  [63:0] io_lm_r_bits_data,
  input         io_lm_aw_ready,
  output        io_lm_aw_valid,
  output [31:0] io_lm_aw_bits_addr,
  input         io_lm_w_ready,
  output        io_lm_w_valid,
  output [63:0] io_lm_w_bits_data,
  output [7:0]  io_lm_w_bits_strb,
  output        io_lm_b_ready,
  input         io_lm_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rstate; // @[LSU.scala 14:23]
  wire  _rstate_T = io_lm_ar_ready & io_lm_ar_valid; // @[Decoupled.scala 52:35]
  wire  _rstate_T_2 = io_lm_r_ready & io_lm_r_valid; // @[Decoupled.scala 52:35]
  reg [1:0] wstate; // @[LSU.scala 19:23]
  wire  _wstate_T = io_lm_aw_ready & io_lm_aw_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _wstate_T_1 = _wstate_T ? 2'h1 : 2'h0; // @[LSU.scala 21:19]
  wire  _wstate_T_2 = io_lm_w_ready & io_lm_w_valid; // @[Decoupled.scala 52:35]
  wire  _wstate_T_4 = io_lm_b_ready & io_lm_b_valid; // @[Decoupled.scala 52:35]
  wire  _io_lm_ar_valid_T_2 = ~reset; // @[LSU.scala 27:40]
  reg [63:0] rdata; // @[Reg.scala 35:20]
  assign io_ls_out_valid = _rstate_T_2 | _wstate_T_4; // @[LSU.scala 39:33]
  assign io_ls_out_bits_rdata = _rstate_T_2 ? io_lm_r_bits_data : rdata; // @[LSU.scala 38:28]
  assign io_lm_ar_valid = rstate == 2'h0 & ~reset & io_ls_in_valid & io_en_r; // @[LSU.scala 27:71]
  assign io_lm_ar_bits_addr = io_ls_in_bits_raddr; // @[LSU.scala 26:21]
  assign io_lm_r_ready = rstate == 2'h1; // @[LSU.scala 28:26]
  assign io_lm_aw_valid = wstate == 2'h0 & _io_lm_ar_valid_T_2 & io_ls_in_valid & io_en_w; // @[LSU.scala 30:71]
  assign io_lm_aw_bits_addr = io_ls_in_bits_waddr; // @[LSU.scala 29:21]
  assign io_lm_w_valid = wstate == 2'h1 & _io_lm_ar_valid_T_2; // @[LSU.scala 33:37]
  assign io_lm_w_bits_data = io_ls_in_bits_wdata; // @[LSU.scala 31:20]
  assign io_lm_w_bits_strb = io_ls_in_bits_wmask; // @[LSU.scala 32:20]
  assign io_lm_b_ready = 1'h1; // @[LSU.scala 34:16]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 14:23]
      rstate <= 2'h0; // @[LSU.scala 14:23]
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      if (_rstate_T_2) begin // @[LSU.scala 17:19]
        rstate <= 2'h0;
      end else begin
        rstate <= 2'h1;
      end
    end else if (2'h0 == rstate) begin // @[Mux.scala 81:58]
      if (_rstate_T) begin // @[LSU.scala 16:19]
        rstate <= 2'h1;
      end else begin
        rstate <= 2'h0;
      end
    end else begin
      rstate <= 2'h0;
    end
    if (reset) begin // @[LSU.scala 19:23]
      wstate <= 2'h0; // @[LSU.scala 19:23]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      if (_wstate_T_4) begin // @[LSU.scala 23:19]
        wstate <= 2'h0;
      end else begin
        wstate <= 2'h2;
      end
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      if (_wstate_T_2) begin // @[LSU.scala 22:19]
        wstate <= 2'h2;
      end else begin
        wstate <= 2'h1;
      end
    end else if (2'h0 == wstate) begin // @[Mux.scala 81:58]
      wstate <= _wstate_T_1;
    end else begin
      wstate <= 2'h0;
    end
    if (reset) begin // @[Reg.scala 35:20]
      rdata <= 64'h0; // @[Reg.scala 35:20]
    end else if (_rstate_T_2) begin // @[Reg.scala 36:18]
      rdata <= io_lm_r_bits_data; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rstate = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  rdata = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mul_cell(
  input          clock,
  input          reset,
  input          io_flush,
  input          io_valid,
  input  [128:0] io_a_in,
  input  [128:0] io_b_in,
  input  [128:0] io_sum_in,
  input          io_last,
  output [128:0] io_a_out,
  output [128:0] io_b_out,
  output [128:0] io_sum_out,
  output         io_ready,
  input  [63:0]  io_a,
  input  [63:0]  io_b,
  output [63:0]  io_A,
  output [63:0]  io_B
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_a; // @[mul.scala 25:22]
  reg [63:0] reg_b; // @[mul.scala 26:22]
  reg [128:0] a_in; // @[mul.scala 36:22]
  reg [128:0] b_in; // @[mul.scala 37:22]
  reg [128:0] sum_in; // @[mul.scala 38:24]
  reg  valid; // @[mul.scala 39:22]
  wire [129:0] _io_a_out_T = {a_in, 1'h0}; // @[mul.scala 56:20]
  wire [128:0] _io_sum_out_T_4 = sum_in - a_in; // @[mul.scala 59:43]
  wire [128:0] _io_sum_out_T_6 = sum_in + a_in; // @[mul.scala 60:24]
  wire [128:0] _io_sum_out_T_7 = io_last ? _io_sum_out_T_4 : _io_sum_out_T_6; // @[mul.scala 59:20]
  assign io_a_out = _io_a_out_T[128:0]; // @[mul.scala 56:12]
  assign io_b_out = {{1'd0}, b_in[128:1]}; // @[mul.scala 57:20]
  assign io_sum_out = ~b_in[0] ? sum_in : _io_sum_out_T_7; // @[mul.scala 58:20]
  assign io_ready = valid; // @[mul.scala 61:12]
  assign io_A = reg_a; // @[mul.scala 33:8]
  assign io_B = reg_b; // @[mul.scala 34:8]
  always @(posedge clock) begin
    if (reset) begin // @[mul.scala 25:22]
      reg_a <= 64'h0; // @[mul.scala 25:22]
    end else if (io_flush) begin // @[mul.scala 27:16]
      reg_a <= 64'h0;
    end else if (io_valid) begin // @[mul.scala 28:15]
      reg_a <= io_a;
    end
    if (reset) begin // @[mul.scala 26:22]
      reg_b <= 64'h0; // @[mul.scala 26:22]
    end else if (io_flush) begin // @[mul.scala 30:16]
      reg_b <= 64'h0;
    end else if (io_valid) begin // @[mul.scala 31:15]
      reg_b <= io_b;
    end
    if (reset) begin // @[mul.scala 36:22]
      a_in <= 129'h0; // @[mul.scala 36:22]
    end else if (io_flush) begin // @[mul.scala 42:17]
      a_in <= 129'h0;
    end else if (io_valid) begin // @[mul.scala 43:16]
      a_in <= io_a_in;
    end
    if (reset) begin // @[mul.scala 37:22]
      b_in <= 129'h0; // @[mul.scala 37:22]
    end else if (io_flush) begin // @[mul.scala 46:17]
      b_in <= 129'h0;
    end else if (io_valid) begin // @[mul.scala 47:16]
      b_in <= io_b_in;
    end
    if (reset) begin // @[mul.scala 38:24]
      sum_in <= 129'h0; // @[mul.scala 38:24]
    end else if (io_flush) begin // @[mul.scala 50:17]
      sum_in <= 129'h0;
    end else if (io_valid) begin // @[mul.scala 51:16]
      sum_in <= io_sum_in;
    end
    if (reset) begin // @[mul.scala 39:22]
      valid <= 1'h0; // @[mul.scala 39:22]
    end else if (io_flush) begin // @[mul.scala 54:17]
      valid <= 1'h0;
    end else begin
      valid <= io_valid;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_a = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  reg_b = _RAND_1[63:0];
  _RAND_2 = {5{`RANDOM}};
  a_in = _RAND_2[128:0];
  _RAND_3 = {5{`RANDOM}};
  b_in = _RAND_3[128:0];
  _RAND_4 = {5{`RANDOM}};
  sum_in = _RAND_4[128:0];
  _RAND_5 = {1{`RANDOM}};
  valid = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mul_pipe(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [1:0]  io_mul_signed,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [63:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  cell_0_clock; // @[mul.scala 95:35]
  wire  cell_0_reset; // @[mul.scala 95:35]
  wire  cell_0_io_flush; // @[mul.scala 95:35]
  wire  cell_0_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_sum_in; // @[mul.scala 95:35]
  wire  cell_0_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_0_io_sum_out; // @[mul.scala 95:35]
  wire  cell_0_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_0_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_0_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_0_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_0_io_B; // @[mul.scala 95:35]
  wire  cell_1_clock; // @[mul.scala 95:35]
  wire  cell_1_reset; // @[mul.scala 95:35]
  wire  cell_1_io_flush; // @[mul.scala 95:35]
  wire  cell_1_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_sum_in; // @[mul.scala 95:35]
  wire  cell_1_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_1_io_sum_out; // @[mul.scala 95:35]
  wire  cell_1_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_1_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_1_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_1_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_1_io_B; // @[mul.scala 95:35]
  wire  cell_2_clock; // @[mul.scala 95:35]
  wire  cell_2_reset; // @[mul.scala 95:35]
  wire  cell_2_io_flush; // @[mul.scala 95:35]
  wire  cell_2_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_sum_in; // @[mul.scala 95:35]
  wire  cell_2_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_2_io_sum_out; // @[mul.scala 95:35]
  wire  cell_2_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_2_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_2_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_2_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_2_io_B; // @[mul.scala 95:35]
  wire  cell_3_clock; // @[mul.scala 95:35]
  wire  cell_3_reset; // @[mul.scala 95:35]
  wire  cell_3_io_flush; // @[mul.scala 95:35]
  wire  cell_3_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_sum_in; // @[mul.scala 95:35]
  wire  cell_3_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_3_io_sum_out; // @[mul.scala 95:35]
  wire  cell_3_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_3_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_3_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_3_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_3_io_B; // @[mul.scala 95:35]
  wire  cell_4_clock; // @[mul.scala 95:35]
  wire  cell_4_reset; // @[mul.scala 95:35]
  wire  cell_4_io_flush; // @[mul.scala 95:35]
  wire  cell_4_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_sum_in; // @[mul.scala 95:35]
  wire  cell_4_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_4_io_sum_out; // @[mul.scala 95:35]
  wire  cell_4_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_4_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_4_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_4_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_4_io_B; // @[mul.scala 95:35]
  wire  cell_5_clock; // @[mul.scala 95:35]
  wire  cell_5_reset; // @[mul.scala 95:35]
  wire  cell_5_io_flush; // @[mul.scala 95:35]
  wire  cell_5_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_sum_in; // @[mul.scala 95:35]
  wire  cell_5_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_5_io_sum_out; // @[mul.scala 95:35]
  wire  cell_5_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_5_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_5_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_5_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_5_io_B; // @[mul.scala 95:35]
  wire  cell_6_clock; // @[mul.scala 95:35]
  wire  cell_6_reset; // @[mul.scala 95:35]
  wire  cell_6_io_flush; // @[mul.scala 95:35]
  wire  cell_6_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_sum_in; // @[mul.scala 95:35]
  wire  cell_6_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_6_io_sum_out; // @[mul.scala 95:35]
  wire  cell_6_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_6_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_6_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_6_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_6_io_B; // @[mul.scala 95:35]
  wire  cell_7_clock; // @[mul.scala 95:35]
  wire  cell_7_reset; // @[mul.scala 95:35]
  wire  cell_7_io_flush; // @[mul.scala 95:35]
  wire  cell_7_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_sum_in; // @[mul.scala 95:35]
  wire  cell_7_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_7_io_sum_out; // @[mul.scala 95:35]
  wire  cell_7_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_7_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_7_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_7_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_7_io_B; // @[mul.scala 95:35]
  wire  cell_8_clock; // @[mul.scala 95:35]
  wire  cell_8_reset; // @[mul.scala 95:35]
  wire  cell_8_io_flush; // @[mul.scala 95:35]
  wire  cell_8_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_sum_in; // @[mul.scala 95:35]
  wire  cell_8_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_8_io_sum_out; // @[mul.scala 95:35]
  wire  cell_8_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_8_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_8_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_8_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_8_io_B; // @[mul.scala 95:35]
  wire  cell_9_clock; // @[mul.scala 95:35]
  wire  cell_9_reset; // @[mul.scala 95:35]
  wire  cell_9_io_flush; // @[mul.scala 95:35]
  wire  cell_9_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_sum_in; // @[mul.scala 95:35]
  wire  cell_9_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_9_io_sum_out; // @[mul.scala 95:35]
  wire  cell_9_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_9_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_9_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_9_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_9_io_B; // @[mul.scala 95:35]
  wire  cell_10_clock; // @[mul.scala 95:35]
  wire  cell_10_reset; // @[mul.scala 95:35]
  wire  cell_10_io_flush; // @[mul.scala 95:35]
  wire  cell_10_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_sum_in; // @[mul.scala 95:35]
  wire  cell_10_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_10_io_sum_out; // @[mul.scala 95:35]
  wire  cell_10_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_10_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_10_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_10_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_10_io_B; // @[mul.scala 95:35]
  wire  cell_11_clock; // @[mul.scala 95:35]
  wire  cell_11_reset; // @[mul.scala 95:35]
  wire  cell_11_io_flush; // @[mul.scala 95:35]
  wire  cell_11_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_sum_in; // @[mul.scala 95:35]
  wire  cell_11_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_11_io_sum_out; // @[mul.scala 95:35]
  wire  cell_11_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_11_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_11_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_11_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_11_io_B; // @[mul.scala 95:35]
  wire  cell_12_clock; // @[mul.scala 95:35]
  wire  cell_12_reset; // @[mul.scala 95:35]
  wire  cell_12_io_flush; // @[mul.scala 95:35]
  wire  cell_12_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_sum_in; // @[mul.scala 95:35]
  wire  cell_12_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_12_io_sum_out; // @[mul.scala 95:35]
  wire  cell_12_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_12_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_12_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_12_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_12_io_B; // @[mul.scala 95:35]
  wire  cell_13_clock; // @[mul.scala 95:35]
  wire  cell_13_reset; // @[mul.scala 95:35]
  wire  cell_13_io_flush; // @[mul.scala 95:35]
  wire  cell_13_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_sum_in; // @[mul.scala 95:35]
  wire  cell_13_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_13_io_sum_out; // @[mul.scala 95:35]
  wire  cell_13_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_13_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_13_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_13_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_13_io_B; // @[mul.scala 95:35]
  wire  cell_14_clock; // @[mul.scala 95:35]
  wire  cell_14_reset; // @[mul.scala 95:35]
  wire  cell_14_io_flush; // @[mul.scala 95:35]
  wire  cell_14_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_sum_in; // @[mul.scala 95:35]
  wire  cell_14_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_14_io_sum_out; // @[mul.scala 95:35]
  wire  cell_14_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_14_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_14_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_14_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_14_io_B; // @[mul.scala 95:35]
  wire  cell_15_clock; // @[mul.scala 95:35]
  wire  cell_15_reset; // @[mul.scala 95:35]
  wire  cell_15_io_flush; // @[mul.scala 95:35]
  wire  cell_15_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_sum_in; // @[mul.scala 95:35]
  wire  cell_15_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_15_io_sum_out; // @[mul.scala 95:35]
  wire  cell_15_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_15_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_15_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_15_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_15_io_B; // @[mul.scala 95:35]
  wire  cell_16_clock; // @[mul.scala 95:35]
  wire  cell_16_reset; // @[mul.scala 95:35]
  wire  cell_16_io_flush; // @[mul.scala 95:35]
  wire  cell_16_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_sum_in; // @[mul.scala 95:35]
  wire  cell_16_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_16_io_sum_out; // @[mul.scala 95:35]
  wire  cell_16_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_16_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_16_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_16_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_16_io_B; // @[mul.scala 95:35]
  wire  cell_17_clock; // @[mul.scala 95:35]
  wire  cell_17_reset; // @[mul.scala 95:35]
  wire  cell_17_io_flush; // @[mul.scala 95:35]
  wire  cell_17_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_sum_in; // @[mul.scala 95:35]
  wire  cell_17_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_17_io_sum_out; // @[mul.scala 95:35]
  wire  cell_17_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_17_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_17_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_17_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_17_io_B; // @[mul.scala 95:35]
  wire  cell_18_clock; // @[mul.scala 95:35]
  wire  cell_18_reset; // @[mul.scala 95:35]
  wire  cell_18_io_flush; // @[mul.scala 95:35]
  wire  cell_18_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_sum_in; // @[mul.scala 95:35]
  wire  cell_18_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_18_io_sum_out; // @[mul.scala 95:35]
  wire  cell_18_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_18_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_18_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_18_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_18_io_B; // @[mul.scala 95:35]
  wire  cell_19_clock; // @[mul.scala 95:35]
  wire  cell_19_reset; // @[mul.scala 95:35]
  wire  cell_19_io_flush; // @[mul.scala 95:35]
  wire  cell_19_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_sum_in; // @[mul.scala 95:35]
  wire  cell_19_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_19_io_sum_out; // @[mul.scala 95:35]
  wire  cell_19_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_19_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_19_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_19_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_19_io_B; // @[mul.scala 95:35]
  wire  cell_20_clock; // @[mul.scala 95:35]
  wire  cell_20_reset; // @[mul.scala 95:35]
  wire  cell_20_io_flush; // @[mul.scala 95:35]
  wire  cell_20_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_sum_in; // @[mul.scala 95:35]
  wire  cell_20_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_20_io_sum_out; // @[mul.scala 95:35]
  wire  cell_20_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_20_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_20_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_20_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_20_io_B; // @[mul.scala 95:35]
  wire  cell_21_clock; // @[mul.scala 95:35]
  wire  cell_21_reset; // @[mul.scala 95:35]
  wire  cell_21_io_flush; // @[mul.scala 95:35]
  wire  cell_21_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_sum_in; // @[mul.scala 95:35]
  wire  cell_21_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_21_io_sum_out; // @[mul.scala 95:35]
  wire  cell_21_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_21_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_21_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_21_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_21_io_B; // @[mul.scala 95:35]
  wire  cell_22_clock; // @[mul.scala 95:35]
  wire  cell_22_reset; // @[mul.scala 95:35]
  wire  cell_22_io_flush; // @[mul.scala 95:35]
  wire  cell_22_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_sum_in; // @[mul.scala 95:35]
  wire  cell_22_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_22_io_sum_out; // @[mul.scala 95:35]
  wire  cell_22_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_22_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_22_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_22_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_22_io_B; // @[mul.scala 95:35]
  wire  cell_23_clock; // @[mul.scala 95:35]
  wire  cell_23_reset; // @[mul.scala 95:35]
  wire  cell_23_io_flush; // @[mul.scala 95:35]
  wire  cell_23_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_sum_in; // @[mul.scala 95:35]
  wire  cell_23_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_23_io_sum_out; // @[mul.scala 95:35]
  wire  cell_23_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_23_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_23_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_23_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_23_io_B; // @[mul.scala 95:35]
  wire  cell_24_clock; // @[mul.scala 95:35]
  wire  cell_24_reset; // @[mul.scala 95:35]
  wire  cell_24_io_flush; // @[mul.scala 95:35]
  wire  cell_24_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_sum_in; // @[mul.scala 95:35]
  wire  cell_24_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_24_io_sum_out; // @[mul.scala 95:35]
  wire  cell_24_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_24_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_24_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_24_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_24_io_B; // @[mul.scala 95:35]
  wire  cell_25_clock; // @[mul.scala 95:35]
  wire  cell_25_reset; // @[mul.scala 95:35]
  wire  cell_25_io_flush; // @[mul.scala 95:35]
  wire  cell_25_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_sum_in; // @[mul.scala 95:35]
  wire  cell_25_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_25_io_sum_out; // @[mul.scala 95:35]
  wire  cell_25_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_25_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_25_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_25_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_25_io_B; // @[mul.scala 95:35]
  wire  cell_26_clock; // @[mul.scala 95:35]
  wire  cell_26_reset; // @[mul.scala 95:35]
  wire  cell_26_io_flush; // @[mul.scala 95:35]
  wire  cell_26_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_sum_in; // @[mul.scala 95:35]
  wire  cell_26_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_26_io_sum_out; // @[mul.scala 95:35]
  wire  cell_26_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_26_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_26_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_26_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_26_io_B; // @[mul.scala 95:35]
  wire  cell_27_clock; // @[mul.scala 95:35]
  wire  cell_27_reset; // @[mul.scala 95:35]
  wire  cell_27_io_flush; // @[mul.scala 95:35]
  wire  cell_27_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_sum_in; // @[mul.scala 95:35]
  wire  cell_27_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_27_io_sum_out; // @[mul.scala 95:35]
  wire  cell_27_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_27_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_27_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_27_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_27_io_B; // @[mul.scala 95:35]
  wire  cell_28_clock; // @[mul.scala 95:35]
  wire  cell_28_reset; // @[mul.scala 95:35]
  wire  cell_28_io_flush; // @[mul.scala 95:35]
  wire  cell_28_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_sum_in; // @[mul.scala 95:35]
  wire  cell_28_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_28_io_sum_out; // @[mul.scala 95:35]
  wire  cell_28_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_28_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_28_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_28_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_28_io_B; // @[mul.scala 95:35]
  wire  cell_29_clock; // @[mul.scala 95:35]
  wire  cell_29_reset; // @[mul.scala 95:35]
  wire  cell_29_io_flush; // @[mul.scala 95:35]
  wire  cell_29_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_sum_in; // @[mul.scala 95:35]
  wire  cell_29_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_29_io_sum_out; // @[mul.scala 95:35]
  wire  cell_29_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_29_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_29_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_29_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_29_io_B; // @[mul.scala 95:35]
  wire  cell_30_clock; // @[mul.scala 95:35]
  wire  cell_30_reset; // @[mul.scala 95:35]
  wire  cell_30_io_flush; // @[mul.scala 95:35]
  wire  cell_30_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_sum_in; // @[mul.scala 95:35]
  wire  cell_30_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_30_io_sum_out; // @[mul.scala 95:35]
  wire  cell_30_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_30_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_30_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_30_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_30_io_B; // @[mul.scala 95:35]
  wire  cell_31_clock; // @[mul.scala 95:35]
  wire  cell_31_reset; // @[mul.scala 95:35]
  wire  cell_31_io_flush; // @[mul.scala 95:35]
  wire  cell_31_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_sum_in; // @[mul.scala 95:35]
  wire  cell_31_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_31_io_sum_out; // @[mul.scala 95:35]
  wire  cell_31_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_31_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_31_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_31_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_31_io_B; // @[mul.scala 95:35]
  wire  cell_32_clock; // @[mul.scala 95:35]
  wire  cell_32_reset; // @[mul.scala 95:35]
  wire  cell_32_io_flush; // @[mul.scala 95:35]
  wire  cell_32_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_sum_in; // @[mul.scala 95:35]
  wire  cell_32_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_32_io_sum_out; // @[mul.scala 95:35]
  wire  cell_32_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_32_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_32_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_32_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_32_io_B; // @[mul.scala 95:35]
  wire  cell_33_clock; // @[mul.scala 95:35]
  wire  cell_33_reset; // @[mul.scala 95:35]
  wire  cell_33_io_flush; // @[mul.scala 95:35]
  wire  cell_33_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_sum_in; // @[mul.scala 95:35]
  wire  cell_33_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_33_io_sum_out; // @[mul.scala 95:35]
  wire  cell_33_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_33_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_33_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_33_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_33_io_B; // @[mul.scala 95:35]
  wire  cell_34_clock; // @[mul.scala 95:35]
  wire  cell_34_reset; // @[mul.scala 95:35]
  wire  cell_34_io_flush; // @[mul.scala 95:35]
  wire  cell_34_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_sum_in; // @[mul.scala 95:35]
  wire  cell_34_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_34_io_sum_out; // @[mul.scala 95:35]
  wire  cell_34_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_34_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_34_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_34_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_34_io_B; // @[mul.scala 95:35]
  wire  cell_35_clock; // @[mul.scala 95:35]
  wire  cell_35_reset; // @[mul.scala 95:35]
  wire  cell_35_io_flush; // @[mul.scala 95:35]
  wire  cell_35_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_sum_in; // @[mul.scala 95:35]
  wire  cell_35_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_35_io_sum_out; // @[mul.scala 95:35]
  wire  cell_35_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_35_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_35_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_35_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_35_io_B; // @[mul.scala 95:35]
  wire  cell_36_clock; // @[mul.scala 95:35]
  wire  cell_36_reset; // @[mul.scala 95:35]
  wire  cell_36_io_flush; // @[mul.scala 95:35]
  wire  cell_36_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_sum_in; // @[mul.scala 95:35]
  wire  cell_36_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_36_io_sum_out; // @[mul.scala 95:35]
  wire  cell_36_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_36_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_36_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_36_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_36_io_B; // @[mul.scala 95:35]
  wire  cell_37_clock; // @[mul.scala 95:35]
  wire  cell_37_reset; // @[mul.scala 95:35]
  wire  cell_37_io_flush; // @[mul.scala 95:35]
  wire  cell_37_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_sum_in; // @[mul.scala 95:35]
  wire  cell_37_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_37_io_sum_out; // @[mul.scala 95:35]
  wire  cell_37_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_37_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_37_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_37_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_37_io_B; // @[mul.scala 95:35]
  wire  cell_38_clock; // @[mul.scala 95:35]
  wire  cell_38_reset; // @[mul.scala 95:35]
  wire  cell_38_io_flush; // @[mul.scala 95:35]
  wire  cell_38_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_sum_in; // @[mul.scala 95:35]
  wire  cell_38_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_38_io_sum_out; // @[mul.scala 95:35]
  wire  cell_38_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_38_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_38_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_38_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_38_io_B; // @[mul.scala 95:35]
  wire  cell_39_clock; // @[mul.scala 95:35]
  wire  cell_39_reset; // @[mul.scala 95:35]
  wire  cell_39_io_flush; // @[mul.scala 95:35]
  wire  cell_39_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_sum_in; // @[mul.scala 95:35]
  wire  cell_39_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_39_io_sum_out; // @[mul.scala 95:35]
  wire  cell_39_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_39_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_39_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_39_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_39_io_B; // @[mul.scala 95:35]
  wire  cell_40_clock; // @[mul.scala 95:35]
  wire  cell_40_reset; // @[mul.scala 95:35]
  wire  cell_40_io_flush; // @[mul.scala 95:35]
  wire  cell_40_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_sum_in; // @[mul.scala 95:35]
  wire  cell_40_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_40_io_sum_out; // @[mul.scala 95:35]
  wire  cell_40_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_40_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_40_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_40_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_40_io_B; // @[mul.scala 95:35]
  wire  cell_41_clock; // @[mul.scala 95:35]
  wire  cell_41_reset; // @[mul.scala 95:35]
  wire  cell_41_io_flush; // @[mul.scala 95:35]
  wire  cell_41_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_sum_in; // @[mul.scala 95:35]
  wire  cell_41_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_41_io_sum_out; // @[mul.scala 95:35]
  wire  cell_41_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_41_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_41_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_41_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_41_io_B; // @[mul.scala 95:35]
  wire  cell_42_clock; // @[mul.scala 95:35]
  wire  cell_42_reset; // @[mul.scala 95:35]
  wire  cell_42_io_flush; // @[mul.scala 95:35]
  wire  cell_42_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_sum_in; // @[mul.scala 95:35]
  wire  cell_42_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_42_io_sum_out; // @[mul.scala 95:35]
  wire  cell_42_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_42_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_42_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_42_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_42_io_B; // @[mul.scala 95:35]
  wire  cell_43_clock; // @[mul.scala 95:35]
  wire  cell_43_reset; // @[mul.scala 95:35]
  wire  cell_43_io_flush; // @[mul.scala 95:35]
  wire  cell_43_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_sum_in; // @[mul.scala 95:35]
  wire  cell_43_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_43_io_sum_out; // @[mul.scala 95:35]
  wire  cell_43_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_43_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_43_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_43_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_43_io_B; // @[mul.scala 95:35]
  wire  cell_44_clock; // @[mul.scala 95:35]
  wire  cell_44_reset; // @[mul.scala 95:35]
  wire  cell_44_io_flush; // @[mul.scala 95:35]
  wire  cell_44_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_sum_in; // @[mul.scala 95:35]
  wire  cell_44_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_44_io_sum_out; // @[mul.scala 95:35]
  wire  cell_44_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_44_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_44_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_44_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_44_io_B; // @[mul.scala 95:35]
  wire  cell_45_clock; // @[mul.scala 95:35]
  wire  cell_45_reset; // @[mul.scala 95:35]
  wire  cell_45_io_flush; // @[mul.scala 95:35]
  wire  cell_45_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_sum_in; // @[mul.scala 95:35]
  wire  cell_45_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_45_io_sum_out; // @[mul.scala 95:35]
  wire  cell_45_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_45_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_45_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_45_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_45_io_B; // @[mul.scala 95:35]
  wire  cell_46_clock; // @[mul.scala 95:35]
  wire  cell_46_reset; // @[mul.scala 95:35]
  wire  cell_46_io_flush; // @[mul.scala 95:35]
  wire  cell_46_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_sum_in; // @[mul.scala 95:35]
  wire  cell_46_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_46_io_sum_out; // @[mul.scala 95:35]
  wire  cell_46_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_46_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_46_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_46_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_46_io_B; // @[mul.scala 95:35]
  wire  cell_47_clock; // @[mul.scala 95:35]
  wire  cell_47_reset; // @[mul.scala 95:35]
  wire  cell_47_io_flush; // @[mul.scala 95:35]
  wire  cell_47_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_sum_in; // @[mul.scala 95:35]
  wire  cell_47_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_47_io_sum_out; // @[mul.scala 95:35]
  wire  cell_47_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_47_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_47_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_47_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_47_io_B; // @[mul.scala 95:35]
  wire  cell_48_clock; // @[mul.scala 95:35]
  wire  cell_48_reset; // @[mul.scala 95:35]
  wire  cell_48_io_flush; // @[mul.scala 95:35]
  wire  cell_48_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_sum_in; // @[mul.scala 95:35]
  wire  cell_48_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_48_io_sum_out; // @[mul.scala 95:35]
  wire  cell_48_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_48_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_48_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_48_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_48_io_B; // @[mul.scala 95:35]
  wire  cell_49_clock; // @[mul.scala 95:35]
  wire  cell_49_reset; // @[mul.scala 95:35]
  wire  cell_49_io_flush; // @[mul.scala 95:35]
  wire  cell_49_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_sum_in; // @[mul.scala 95:35]
  wire  cell_49_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_49_io_sum_out; // @[mul.scala 95:35]
  wire  cell_49_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_49_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_49_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_49_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_49_io_B; // @[mul.scala 95:35]
  wire  cell_50_clock; // @[mul.scala 95:35]
  wire  cell_50_reset; // @[mul.scala 95:35]
  wire  cell_50_io_flush; // @[mul.scala 95:35]
  wire  cell_50_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_sum_in; // @[mul.scala 95:35]
  wire  cell_50_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_50_io_sum_out; // @[mul.scala 95:35]
  wire  cell_50_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_50_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_50_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_50_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_50_io_B; // @[mul.scala 95:35]
  wire  cell_51_clock; // @[mul.scala 95:35]
  wire  cell_51_reset; // @[mul.scala 95:35]
  wire  cell_51_io_flush; // @[mul.scala 95:35]
  wire  cell_51_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_sum_in; // @[mul.scala 95:35]
  wire  cell_51_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_51_io_sum_out; // @[mul.scala 95:35]
  wire  cell_51_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_51_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_51_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_51_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_51_io_B; // @[mul.scala 95:35]
  wire  cell_52_clock; // @[mul.scala 95:35]
  wire  cell_52_reset; // @[mul.scala 95:35]
  wire  cell_52_io_flush; // @[mul.scala 95:35]
  wire  cell_52_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_sum_in; // @[mul.scala 95:35]
  wire  cell_52_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_52_io_sum_out; // @[mul.scala 95:35]
  wire  cell_52_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_52_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_52_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_52_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_52_io_B; // @[mul.scala 95:35]
  wire  cell_53_clock; // @[mul.scala 95:35]
  wire  cell_53_reset; // @[mul.scala 95:35]
  wire  cell_53_io_flush; // @[mul.scala 95:35]
  wire  cell_53_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_sum_in; // @[mul.scala 95:35]
  wire  cell_53_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_53_io_sum_out; // @[mul.scala 95:35]
  wire  cell_53_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_53_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_53_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_53_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_53_io_B; // @[mul.scala 95:35]
  wire  cell_54_clock; // @[mul.scala 95:35]
  wire  cell_54_reset; // @[mul.scala 95:35]
  wire  cell_54_io_flush; // @[mul.scala 95:35]
  wire  cell_54_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_sum_in; // @[mul.scala 95:35]
  wire  cell_54_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_54_io_sum_out; // @[mul.scala 95:35]
  wire  cell_54_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_54_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_54_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_54_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_54_io_B; // @[mul.scala 95:35]
  wire  cell_55_clock; // @[mul.scala 95:35]
  wire  cell_55_reset; // @[mul.scala 95:35]
  wire  cell_55_io_flush; // @[mul.scala 95:35]
  wire  cell_55_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_sum_in; // @[mul.scala 95:35]
  wire  cell_55_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_55_io_sum_out; // @[mul.scala 95:35]
  wire  cell_55_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_55_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_55_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_55_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_55_io_B; // @[mul.scala 95:35]
  wire  cell_56_clock; // @[mul.scala 95:35]
  wire  cell_56_reset; // @[mul.scala 95:35]
  wire  cell_56_io_flush; // @[mul.scala 95:35]
  wire  cell_56_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_sum_in; // @[mul.scala 95:35]
  wire  cell_56_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_56_io_sum_out; // @[mul.scala 95:35]
  wire  cell_56_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_56_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_56_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_56_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_56_io_B; // @[mul.scala 95:35]
  wire  cell_57_clock; // @[mul.scala 95:35]
  wire  cell_57_reset; // @[mul.scala 95:35]
  wire  cell_57_io_flush; // @[mul.scala 95:35]
  wire  cell_57_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_sum_in; // @[mul.scala 95:35]
  wire  cell_57_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_57_io_sum_out; // @[mul.scala 95:35]
  wire  cell_57_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_57_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_57_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_57_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_57_io_B; // @[mul.scala 95:35]
  wire  cell_58_clock; // @[mul.scala 95:35]
  wire  cell_58_reset; // @[mul.scala 95:35]
  wire  cell_58_io_flush; // @[mul.scala 95:35]
  wire  cell_58_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_sum_in; // @[mul.scala 95:35]
  wire  cell_58_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_58_io_sum_out; // @[mul.scala 95:35]
  wire  cell_58_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_58_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_58_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_58_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_58_io_B; // @[mul.scala 95:35]
  wire  cell_59_clock; // @[mul.scala 95:35]
  wire  cell_59_reset; // @[mul.scala 95:35]
  wire  cell_59_io_flush; // @[mul.scala 95:35]
  wire  cell_59_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_sum_in; // @[mul.scala 95:35]
  wire  cell_59_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_59_io_sum_out; // @[mul.scala 95:35]
  wire  cell_59_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_59_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_59_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_59_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_59_io_B; // @[mul.scala 95:35]
  wire  cell_60_clock; // @[mul.scala 95:35]
  wire  cell_60_reset; // @[mul.scala 95:35]
  wire  cell_60_io_flush; // @[mul.scala 95:35]
  wire  cell_60_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_sum_in; // @[mul.scala 95:35]
  wire  cell_60_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_60_io_sum_out; // @[mul.scala 95:35]
  wire  cell_60_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_60_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_60_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_60_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_60_io_B; // @[mul.scala 95:35]
  wire  cell_61_clock; // @[mul.scala 95:35]
  wire  cell_61_reset; // @[mul.scala 95:35]
  wire  cell_61_io_flush; // @[mul.scala 95:35]
  wire  cell_61_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_sum_in; // @[mul.scala 95:35]
  wire  cell_61_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_61_io_sum_out; // @[mul.scala 95:35]
  wire  cell_61_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_61_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_61_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_61_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_61_io_B; // @[mul.scala 95:35]
  wire  cell_62_clock; // @[mul.scala 95:35]
  wire  cell_62_reset; // @[mul.scala 95:35]
  wire  cell_62_io_flush; // @[mul.scala 95:35]
  wire  cell_62_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_sum_in; // @[mul.scala 95:35]
  wire  cell_62_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_62_io_sum_out; // @[mul.scala 95:35]
  wire  cell_62_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_62_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_62_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_62_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_62_io_B; // @[mul.scala 95:35]
  wire  cell_63_clock; // @[mul.scala 95:35]
  wire  cell_63_reset; // @[mul.scala 95:35]
  wire  cell_63_io_flush; // @[mul.scala 95:35]
  wire  cell_63_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_sum_in; // @[mul.scala 95:35]
  wire  cell_63_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_63_io_sum_out; // @[mul.scala 95:35]
  wire  cell_63_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_63_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_63_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_63_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_63_io_B; // @[mul.scala 95:35]
  wire  cell_64_clock; // @[mul.scala 95:35]
  wire  cell_64_reset; // @[mul.scala 95:35]
  wire  cell_64_io_flush; // @[mul.scala 95:35]
  wire  cell_64_io_valid; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_a_in; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_b_in; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_sum_in; // @[mul.scala 95:35]
  wire  cell_64_io_last; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_a_out; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_b_out; // @[mul.scala 95:35]
  wire [128:0] cell_64_io_sum_out; // @[mul.scala 95:35]
  wire  cell_64_io_ready; // @[mul.scala 95:35]
  wire [63:0] cell_64_io_a; // @[mul.scala 95:35]
  wire [63:0] cell_64_io_b; // @[mul.scala 95:35]
  wire [63:0] cell_64_io_A; // @[mul.scala 95:35]
  wire [63:0] cell_64_io_B; // @[mul.scala 95:35]
  reg [128:0] a; // @[mul.scala 77:20]
  reg [128:0] b; // @[mul.scala 78:20]
  reg  valid; // @[mul.scala 79:24]
  wire  _a_T_2 = io_mul_valid & io_mul_signed[1]; // @[mul.scala 82:26]
  wire [64:0] _a_T_16 = io_multiplicand[63] ? 65'h1ffffffffffffffff : 65'h0; // @[Bitwise.scala 77:12]
  wire [128:0] _a_T_17 = {_a_T_16,io_multiplicand}; // @[Cat.scala 33:92]
  wire [128:0] _a_T_19 = io_mul_valid ? {{65'd0}, io_multiplicand} : a; // @[mul.scala 84:12]
  wire [128:0] _a_T_20 = _a_T_2 ? _a_T_17 : _a_T_19; // @[mul.scala 83:12]
  wire [160:0] _a_T_21 = {{32'd0}, _a_T_20}; // @[mul.scala 82:12]
  wire [64:0] _b_T_16 = io_multiplier[63] ? 65'h1ffffffffffffffff : 65'h0; // @[Bitwise.scala 77:12]
  wire [128:0] _b_T_17 = {_b_T_16,io_multiplier}; // @[Cat.scala 33:92]
  wire [128:0] _b_T_19 = io_mul_valid ? {{65'd0}, io_multiplier} : b; // @[mul.scala 90:12]
  wire [128:0] _b_T_20 = _a_T_2 ? _b_T_17 : _b_T_19; // @[mul.scala 89:12]
  wire [160:0] _b_T_21 = {{32'd0}, _b_T_20}; // @[mul.scala 88:12]
  wire [127:0] _T_1 = cell_64_io_A * cell_64_io_B; // @[mul.scala 124:64]
  wire [128:0] _GEN_0 = {{1'd0}, _T_1}; // @[mul.scala 124:45]
  wire [160:0] _GEN_1 = reset ? 161'h0 : _a_T_21; // @[mul.scala 77:{20,20} 81:7]
  wire [160:0] _GEN_2 = reset ? 161'h0 : _b_T_21; // @[mul.scala 78:{20,20} 87:7]
  mul_cell cell_0 ( // @[mul.scala 95:35]
    .clock(cell_0_clock),
    .reset(cell_0_reset),
    .io_flush(cell_0_io_flush),
    .io_valid(cell_0_io_valid),
    .io_a_in(cell_0_io_a_in),
    .io_b_in(cell_0_io_b_in),
    .io_sum_in(cell_0_io_sum_in),
    .io_last(cell_0_io_last),
    .io_a_out(cell_0_io_a_out),
    .io_b_out(cell_0_io_b_out),
    .io_sum_out(cell_0_io_sum_out),
    .io_ready(cell_0_io_ready),
    .io_a(cell_0_io_a),
    .io_b(cell_0_io_b),
    .io_A(cell_0_io_A),
    .io_B(cell_0_io_B)
  );
  mul_cell cell_1 ( // @[mul.scala 95:35]
    .clock(cell_1_clock),
    .reset(cell_1_reset),
    .io_flush(cell_1_io_flush),
    .io_valid(cell_1_io_valid),
    .io_a_in(cell_1_io_a_in),
    .io_b_in(cell_1_io_b_in),
    .io_sum_in(cell_1_io_sum_in),
    .io_last(cell_1_io_last),
    .io_a_out(cell_1_io_a_out),
    .io_b_out(cell_1_io_b_out),
    .io_sum_out(cell_1_io_sum_out),
    .io_ready(cell_1_io_ready),
    .io_a(cell_1_io_a),
    .io_b(cell_1_io_b),
    .io_A(cell_1_io_A),
    .io_B(cell_1_io_B)
  );
  mul_cell cell_2 ( // @[mul.scala 95:35]
    .clock(cell_2_clock),
    .reset(cell_2_reset),
    .io_flush(cell_2_io_flush),
    .io_valid(cell_2_io_valid),
    .io_a_in(cell_2_io_a_in),
    .io_b_in(cell_2_io_b_in),
    .io_sum_in(cell_2_io_sum_in),
    .io_last(cell_2_io_last),
    .io_a_out(cell_2_io_a_out),
    .io_b_out(cell_2_io_b_out),
    .io_sum_out(cell_2_io_sum_out),
    .io_ready(cell_2_io_ready),
    .io_a(cell_2_io_a),
    .io_b(cell_2_io_b),
    .io_A(cell_2_io_A),
    .io_B(cell_2_io_B)
  );
  mul_cell cell_3 ( // @[mul.scala 95:35]
    .clock(cell_3_clock),
    .reset(cell_3_reset),
    .io_flush(cell_3_io_flush),
    .io_valid(cell_3_io_valid),
    .io_a_in(cell_3_io_a_in),
    .io_b_in(cell_3_io_b_in),
    .io_sum_in(cell_3_io_sum_in),
    .io_last(cell_3_io_last),
    .io_a_out(cell_3_io_a_out),
    .io_b_out(cell_3_io_b_out),
    .io_sum_out(cell_3_io_sum_out),
    .io_ready(cell_3_io_ready),
    .io_a(cell_3_io_a),
    .io_b(cell_3_io_b),
    .io_A(cell_3_io_A),
    .io_B(cell_3_io_B)
  );
  mul_cell cell_4 ( // @[mul.scala 95:35]
    .clock(cell_4_clock),
    .reset(cell_4_reset),
    .io_flush(cell_4_io_flush),
    .io_valid(cell_4_io_valid),
    .io_a_in(cell_4_io_a_in),
    .io_b_in(cell_4_io_b_in),
    .io_sum_in(cell_4_io_sum_in),
    .io_last(cell_4_io_last),
    .io_a_out(cell_4_io_a_out),
    .io_b_out(cell_4_io_b_out),
    .io_sum_out(cell_4_io_sum_out),
    .io_ready(cell_4_io_ready),
    .io_a(cell_4_io_a),
    .io_b(cell_4_io_b),
    .io_A(cell_4_io_A),
    .io_B(cell_4_io_B)
  );
  mul_cell cell_5 ( // @[mul.scala 95:35]
    .clock(cell_5_clock),
    .reset(cell_5_reset),
    .io_flush(cell_5_io_flush),
    .io_valid(cell_5_io_valid),
    .io_a_in(cell_5_io_a_in),
    .io_b_in(cell_5_io_b_in),
    .io_sum_in(cell_5_io_sum_in),
    .io_last(cell_5_io_last),
    .io_a_out(cell_5_io_a_out),
    .io_b_out(cell_5_io_b_out),
    .io_sum_out(cell_5_io_sum_out),
    .io_ready(cell_5_io_ready),
    .io_a(cell_5_io_a),
    .io_b(cell_5_io_b),
    .io_A(cell_5_io_A),
    .io_B(cell_5_io_B)
  );
  mul_cell cell_6 ( // @[mul.scala 95:35]
    .clock(cell_6_clock),
    .reset(cell_6_reset),
    .io_flush(cell_6_io_flush),
    .io_valid(cell_6_io_valid),
    .io_a_in(cell_6_io_a_in),
    .io_b_in(cell_6_io_b_in),
    .io_sum_in(cell_6_io_sum_in),
    .io_last(cell_6_io_last),
    .io_a_out(cell_6_io_a_out),
    .io_b_out(cell_6_io_b_out),
    .io_sum_out(cell_6_io_sum_out),
    .io_ready(cell_6_io_ready),
    .io_a(cell_6_io_a),
    .io_b(cell_6_io_b),
    .io_A(cell_6_io_A),
    .io_B(cell_6_io_B)
  );
  mul_cell cell_7 ( // @[mul.scala 95:35]
    .clock(cell_7_clock),
    .reset(cell_7_reset),
    .io_flush(cell_7_io_flush),
    .io_valid(cell_7_io_valid),
    .io_a_in(cell_7_io_a_in),
    .io_b_in(cell_7_io_b_in),
    .io_sum_in(cell_7_io_sum_in),
    .io_last(cell_7_io_last),
    .io_a_out(cell_7_io_a_out),
    .io_b_out(cell_7_io_b_out),
    .io_sum_out(cell_7_io_sum_out),
    .io_ready(cell_7_io_ready),
    .io_a(cell_7_io_a),
    .io_b(cell_7_io_b),
    .io_A(cell_7_io_A),
    .io_B(cell_7_io_B)
  );
  mul_cell cell_8 ( // @[mul.scala 95:35]
    .clock(cell_8_clock),
    .reset(cell_8_reset),
    .io_flush(cell_8_io_flush),
    .io_valid(cell_8_io_valid),
    .io_a_in(cell_8_io_a_in),
    .io_b_in(cell_8_io_b_in),
    .io_sum_in(cell_8_io_sum_in),
    .io_last(cell_8_io_last),
    .io_a_out(cell_8_io_a_out),
    .io_b_out(cell_8_io_b_out),
    .io_sum_out(cell_8_io_sum_out),
    .io_ready(cell_8_io_ready),
    .io_a(cell_8_io_a),
    .io_b(cell_8_io_b),
    .io_A(cell_8_io_A),
    .io_B(cell_8_io_B)
  );
  mul_cell cell_9 ( // @[mul.scala 95:35]
    .clock(cell_9_clock),
    .reset(cell_9_reset),
    .io_flush(cell_9_io_flush),
    .io_valid(cell_9_io_valid),
    .io_a_in(cell_9_io_a_in),
    .io_b_in(cell_9_io_b_in),
    .io_sum_in(cell_9_io_sum_in),
    .io_last(cell_9_io_last),
    .io_a_out(cell_9_io_a_out),
    .io_b_out(cell_9_io_b_out),
    .io_sum_out(cell_9_io_sum_out),
    .io_ready(cell_9_io_ready),
    .io_a(cell_9_io_a),
    .io_b(cell_9_io_b),
    .io_A(cell_9_io_A),
    .io_B(cell_9_io_B)
  );
  mul_cell cell_10 ( // @[mul.scala 95:35]
    .clock(cell_10_clock),
    .reset(cell_10_reset),
    .io_flush(cell_10_io_flush),
    .io_valid(cell_10_io_valid),
    .io_a_in(cell_10_io_a_in),
    .io_b_in(cell_10_io_b_in),
    .io_sum_in(cell_10_io_sum_in),
    .io_last(cell_10_io_last),
    .io_a_out(cell_10_io_a_out),
    .io_b_out(cell_10_io_b_out),
    .io_sum_out(cell_10_io_sum_out),
    .io_ready(cell_10_io_ready),
    .io_a(cell_10_io_a),
    .io_b(cell_10_io_b),
    .io_A(cell_10_io_A),
    .io_B(cell_10_io_B)
  );
  mul_cell cell_11 ( // @[mul.scala 95:35]
    .clock(cell_11_clock),
    .reset(cell_11_reset),
    .io_flush(cell_11_io_flush),
    .io_valid(cell_11_io_valid),
    .io_a_in(cell_11_io_a_in),
    .io_b_in(cell_11_io_b_in),
    .io_sum_in(cell_11_io_sum_in),
    .io_last(cell_11_io_last),
    .io_a_out(cell_11_io_a_out),
    .io_b_out(cell_11_io_b_out),
    .io_sum_out(cell_11_io_sum_out),
    .io_ready(cell_11_io_ready),
    .io_a(cell_11_io_a),
    .io_b(cell_11_io_b),
    .io_A(cell_11_io_A),
    .io_B(cell_11_io_B)
  );
  mul_cell cell_12 ( // @[mul.scala 95:35]
    .clock(cell_12_clock),
    .reset(cell_12_reset),
    .io_flush(cell_12_io_flush),
    .io_valid(cell_12_io_valid),
    .io_a_in(cell_12_io_a_in),
    .io_b_in(cell_12_io_b_in),
    .io_sum_in(cell_12_io_sum_in),
    .io_last(cell_12_io_last),
    .io_a_out(cell_12_io_a_out),
    .io_b_out(cell_12_io_b_out),
    .io_sum_out(cell_12_io_sum_out),
    .io_ready(cell_12_io_ready),
    .io_a(cell_12_io_a),
    .io_b(cell_12_io_b),
    .io_A(cell_12_io_A),
    .io_B(cell_12_io_B)
  );
  mul_cell cell_13 ( // @[mul.scala 95:35]
    .clock(cell_13_clock),
    .reset(cell_13_reset),
    .io_flush(cell_13_io_flush),
    .io_valid(cell_13_io_valid),
    .io_a_in(cell_13_io_a_in),
    .io_b_in(cell_13_io_b_in),
    .io_sum_in(cell_13_io_sum_in),
    .io_last(cell_13_io_last),
    .io_a_out(cell_13_io_a_out),
    .io_b_out(cell_13_io_b_out),
    .io_sum_out(cell_13_io_sum_out),
    .io_ready(cell_13_io_ready),
    .io_a(cell_13_io_a),
    .io_b(cell_13_io_b),
    .io_A(cell_13_io_A),
    .io_B(cell_13_io_B)
  );
  mul_cell cell_14 ( // @[mul.scala 95:35]
    .clock(cell_14_clock),
    .reset(cell_14_reset),
    .io_flush(cell_14_io_flush),
    .io_valid(cell_14_io_valid),
    .io_a_in(cell_14_io_a_in),
    .io_b_in(cell_14_io_b_in),
    .io_sum_in(cell_14_io_sum_in),
    .io_last(cell_14_io_last),
    .io_a_out(cell_14_io_a_out),
    .io_b_out(cell_14_io_b_out),
    .io_sum_out(cell_14_io_sum_out),
    .io_ready(cell_14_io_ready),
    .io_a(cell_14_io_a),
    .io_b(cell_14_io_b),
    .io_A(cell_14_io_A),
    .io_B(cell_14_io_B)
  );
  mul_cell cell_15 ( // @[mul.scala 95:35]
    .clock(cell_15_clock),
    .reset(cell_15_reset),
    .io_flush(cell_15_io_flush),
    .io_valid(cell_15_io_valid),
    .io_a_in(cell_15_io_a_in),
    .io_b_in(cell_15_io_b_in),
    .io_sum_in(cell_15_io_sum_in),
    .io_last(cell_15_io_last),
    .io_a_out(cell_15_io_a_out),
    .io_b_out(cell_15_io_b_out),
    .io_sum_out(cell_15_io_sum_out),
    .io_ready(cell_15_io_ready),
    .io_a(cell_15_io_a),
    .io_b(cell_15_io_b),
    .io_A(cell_15_io_A),
    .io_B(cell_15_io_B)
  );
  mul_cell cell_16 ( // @[mul.scala 95:35]
    .clock(cell_16_clock),
    .reset(cell_16_reset),
    .io_flush(cell_16_io_flush),
    .io_valid(cell_16_io_valid),
    .io_a_in(cell_16_io_a_in),
    .io_b_in(cell_16_io_b_in),
    .io_sum_in(cell_16_io_sum_in),
    .io_last(cell_16_io_last),
    .io_a_out(cell_16_io_a_out),
    .io_b_out(cell_16_io_b_out),
    .io_sum_out(cell_16_io_sum_out),
    .io_ready(cell_16_io_ready),
    .io_a(cell_16_io_a),
    .io_b(cell_16_io_b),
    .io_A(cell_16_io_A),
    .io_B(cell_16_io_B)
  );
  mul_cell cell_17 ( // @[mul.scala 95:35]
    .clock(cell_17_clock),
    .reset(cell_17_reset),
    .io_flush(cell_17_io_flush),
    .io_valid(cell_17_io_valid),
    .io_a_in(cell_17_io_a_in),
    .io_b_in(cell_17_io_b_in),
    .io_sum_in(cell_17_io_sum_in),
    .io_last(cell_17_io_last),
    .io_a_out(cell_17_io_a_out),
    .io_b_out(cell_17_io_b_out),
    .io_sum_out(cell_17_io_sum_out),
    .io_ready(cell_17_io_ready),
    .io_a(cell_17_io_a),
    .io_b(cell_17_io_b),
    .io_A(cell_17_io_A),
    .io_B(cell_17_io_B)
  );
  mul_cell cell_18 ( // @[mul.scala 95:35]
    .clock(cell_18_clock),
    .reset(cell_18_reset),
    .io_flush(cell_18_io_flush),
    .io_valid(cell_18_io_valid),
    .io_a_in(cell_18_io_a_in),
    .io_b_in(cell_18_io_b_in),
    .io_sum_in(cell_18_io_sum_in),
    .io_last(cell_18_io_last),
    .io_a_out(cell_18_io_a_out),
    .io_b_out(cell_18_io_b_out),
    .io_sum_out(cell_18_io_sum_out),
    .io_ready(cell_18_io_ready),
    .io_a(cell_18_io_a),
    .io_b(cell_18_io_b),
    .io_A(cell_18_io_A),
    .io_B(cell_18_io_B)
  );
  mul_cell cell_19 ( // @[mul.scala 95:35]
    .clock(cell_19_clock),
    .reset(cell_19_reset),
    .io_flush(cell_19_io_flush),
    .io_valid(cell_19_io_valid),
    .io_a_in(cell_19_io_a_in),
    .io_b_in(cell_19_io_b_in),
    .io_sum_in(cell_19_io_sum_in),
    .io_last(cell_19_io_last),
    .io_a_out(cell_19_io_a_out),
    .io_b_out(cell_19_io_b_out),
    .io_sum_out(cell_19_io_sum_out),
    .io_ready(cell_19_io_ready),
    .io_a(cell_19_io_a),
    .io_b(cell_19_io_b),
    .io_A(cell_19_io_A),
    .io_B(cell_19_io_B)
  );
  mul_cell cell_20 ( // @[mul.scala 95:35]
    .clock(cell_20_clock),
    .reset(cell_20_reset),
    .io_flush(cell_20_io_flush),
    .io_valid(cell_20_io_valid),
    .io_a_in(cell_20_io_a_in),
    .io_b_in(cell_20_io_b_in),
    .io_sum_in(cell_20_io_sum_in),
    .io_last(cell_20_io_last),
    .io_a_out(cell_20_io_a_out),
    .io_b_out(cell_20_io_b_out),
    .io_sum_out(cell_20_io_sum_out),
    .io_ready(cell_20_io_ready),
    .io_a(cell_20_io_a),
    .io_b(cell_20_io_b),
    .io_A(cell_20_io_A),
    .io_B(cell_20_io_B)
  );
  mul_cell cell_21 ( // @[mul.scala 95:35]
    .clock(cell_21_clock),
    .reset(cell_21_reset),
    .io_flush(cell_21_io_flush),
    .io_valid(cell_21_io_valid),
    .io_a_in(cell_21_io_a_in),
    .io_b_in(cell_21_io_b_in),
    .io_sum_in(cell_21_io_sum_in),
    .io_last(cell_21_io_last),
    .io_a_out(cell_21_io_a_out),
    .io_b_out(cell_21_io_b_out),
    .io_sum_out(cell_21_io_sum_out),
    .io_ready(cell_21_io_ready),
    .io_a(cell_21_io_a),
    .io_b(cell_21_io_b),
    .io_A(cell_21_io_A),
    .io_B(cell_21_io_B)
  );
  mul_cell cell_22 ( // @[mul.scala 95:35]
    .clock(cell_22_clock),
    .reset(cell_22_reset),
    .io_flush(cell_22_io_flush),
    .io_valid(cell_22_io_valid),
    .io_a_in(cell_22_io_a_in),
    .io_b_in(cell_22_io_b_in),
    .io_sum_in(cell_22_io_sum_in),
    .io_last(cell_22_io_last),
    .io_a_out(cell_22_io_a_out),
    .io_b_out(cell_22_io_b_out),
    .io_sum_out(cell_22_io_sum_out),
    .io_ready(cell_22_io_ready),
    .io_a(cell_22_io_a),
    .io_b(cell_22_io_b),
    .io_A(cell_22_io_A),
    .io_B(cell_22_io_B)
  );
  mul_cell cell_23 ( // @[mul.scala 95:35]
    .clock(cell_23_clock),
    .reset(cell_23_reset),
    .io_flush(cell_23_io_flush),
    .io_valid(cell_23_io_valid),
    .io_a_in(cell_23_io_a_in),
    .io_b_in(cell_23_io_b_in),
    .io_sum_in(cell_23_io_sum_in),
    .io_last(cell_23_io_last),
    .io_a_out(cell_23_io_a_out),
    .io_b_out(cell_23_io_b_out),
    .io_sum_out(cell_23_io_sum_out),
    .io_ready(cell_23_io_ready),
    .io_a(cell_23_io_a),
    .io_b(cell_23_io_b),
    .io_A(cell_23_io_A),
    .io_B(cell_23_io_B)
  );
  mul_cell cell_24 ( // @[mul.scala 95:35]
    .clock(cell_24_clock),
    .reset(cell_24_reset),
    .io_flush(cell_24_io_flush),
    .io_valid(cell_24_io_valid),
    .io_a_in(cell_24_io_a_in),
    .io_b_in(cell_24_io_b_in),
    .io_sum_in(cell_24_io_sum_in),
    .io_last(cell_24_io_last),
    .io_a_out(cell_24_io_a_out),
    .io_b_out(cell_24_io_b_out),
    .io_sum_out(cell_24_io_sum_out),
    .io_ready(cell_24_io_ready),
    .io_a(cell_24_io_a),
    .io_b(cell_24_io_b),
    .io_A(cell_24_io_A),
    .io_B(cell_24_io_B)
  );
  mul_cell cell_25 ( // @[mul.scala 95:35]
    .clock(cell_25_clock),
    .reset(cell_25_reset),
    .io_flush(cell_25_io_flush),
    .io_valid(cell_25_io_valid),
    .io_a_in(cell_25_io_a_in),
    .io_b_in(cell_25_io_b_in),
    .io_sum_in(cell_25_io_sum_in),
    .io_last(cell_25_io_last),
    .io_a_out(cell_25_io_a_out),
    .io_b_out(cell_25_io_b_out),
    .io_sum_out(cell_25_io_sum_out),
    .io_ready(cell_25_io_ready),
    .io_a(cell_25_io_a),
    .io_b(cell_25_io_b),
    .io_A(cell_25_io_A),
    .io_B(cell_25_io_B)
  );
  mul_cell cell_26 ( // @[mul.scala 95:35]
    .clock(cell_26_clock),
    .reset(cell_26_reset),
    .io_flush(cell_26_io_flush),
    .io_valid(cell_26_io_valid),
    .io_a_in(cell_26_io_a_in),
    .io_b_in(cell_26_io_b_in),
    .io_sum_in(cell_26_io_sum_in),
    .io_last(cell_26_io_last),
    .io_a_out(cell_26_io_a_out),
    .io_b_out(cell_26_io_b_out),
    .io_sum_out(cell_26_io_sum_out),
    .io_ready(cell_26_io_ready),
    .io_a(cell_26_io_a),
    .io_b(cell_26_io_b),
    .io_A(cell_26_io_A),
    .io_B(cell_26_io_B)
  );
  mul_cell cell_27 ( // @[mul.scala 95:35]
    .clock(cell_27_clock),
    .reset(cell_27_reset),
    .io_flush(cell_27_io_flush),
    .io_valid(cell_27_io_valid),
    .io_a_in(cell_27_io_a_in),
    .io_b_in(cell_27_io_b_in),
    .io_sum_in(cell_27_io_sum_in),
    .io_last(cell_27_io_last),
    .io_a_out(cell_27_io_a_out),
    .io_b_out(cell_27_io_b_out),
    .io_sum_out(cell_27_io_sum_out),
    .io_ready(cell_27_io_ready),
    .io_a(cell_27_io_a),
    .io_b(cell_27_io_b),
    .io_A(cell_27_io_A),
    .io_B(cell_27_io_B)
  );
  mul_cell cell_28 ( // @[mul.scala 95:35]
    .clock(cell_28_clock),
    .reset(cell_28_reset),
    .io_flush(cell_28_io_flush),
    .io_valid(cell_28_io_valid),
    .io_a_in(cell_28_io_a_in),
    .io_b_in(cell_28_io_b_in),
    .io_sum_in(cell_28_io_sum_in),
    .io_last(cell_28_io_last),
    .io_a_out(cell_28_io_a_out),
    .io_b_out(cell_28_io_b_out),
    .io_sum_out(cell_28_io_sum_out),
    .io_ready(cell_28_io_ready),
    .io_a(cell_28_io_a),
    .io_b(cell_28_io_b),
    .io_A(cell_28_io_A),
    .io_B(cell_28_io_B)
  );
  mul_cell cell_29 ( // @[mul.scala 95:35]
    .clock(cell_29_clock),
    .reset(cell_29_reset),
    .io_flush(cell_29_io_flush),
    .io_valid(cell_29_io_valid),
    .io_a_in(cell_29_io_a_in),
    .io_b_in(cell_29_io_b_in),
    .io_sum_in(cell_29_io_sum_in),
    .io_last(cell_29_io_last),
    .io_a_out(cell_29_io_a_out),
    .io_b_out(cell_29_io_b_out),
    .io_sum_out(cell_29_io_sum_out),
    .io_ready(cell_29_io_ready),
    .io_a(cell_29_io_a),
    .io_b(cell_29_io_b),
    .io_A(cell_29_io_A),
    .io_B(cell_29_io_B)
  );
  mul_cell cell_30 ( // @[mul.scala 95:35]
    .clock(cell_30_clock),
    .reset(cell_30_reset),
    .io_flush(cell_30_io_flush),
    .io_valid(cell_30_io_valid),
    .io_a_in(cell_30_io_a_in),
    .io_b_in(cell_30_io_b_in),
    .io_sum_in(cell_30_io_sum_in),
    .io_last(cell_30_io_last),
    .io_a_out(cell_30_io_a_out),
    .io_b_out(cell_30_io_b_out),
    .io_sum_out(cell_30_io_sum_out),
    .io_ready(cell_30_io_ready),
    .io_a(cell_30_io_a),
    .io_b(cell_30_io_b),
    .io_A(cell_30_io_A),
    .io_B(cell_30_io_B)
  );
  mul_cell cell_31 ( // @[mul.scala 95:35]
    .clock(cell_31_clock),
    .reset(cell_31_reset),
    .io_flush(cell_31_io_flush),
    .io_valid(cell_31_io_valid),
    .io_a_in(cell_31_io_a_in),
    .io_b_in(cell_31_io_b_in),
    .io_sum_in(cell_31_io_sum_in),
    .io_last(cell_31_io_last),
    .io_a_out(cell_31_io_a_out),
    .io_b_out(cell_31_io_b_out),
    .io_sum_out(cell_31_io_sum_out),
    .io_ready(cell_31_io_ready),
    .io_a(cell_31_io_a),
    .io_b(cell_31_io_b),
    .io_A(cell_31_io_A),
    .io_B(cell_31_io_B)
  );
  mul_cell cell_32 ( // @[mul.scala 95:35]
    .clock(cell_32_clock),
    .reset(cell_32_reset),
    .io_flush(cell_32_io_flush),
    .io_valid(cell_32_io_valid),
    .io_a_in(cell_32_io_a_in),
    .io_b_in(cell_32_io_b_in),
    .io_sum_in(cell_32_io_sum_in),
    .io_last(cell_32_io_last),
    .io_a_out(cell_32_io_a_out),
    .io_b_out(cell_32_io_b_out),
    .io_sum_out(cell_32_io_sum_out),
    .io_ready(cell_32_io_ready),
    .io_a(cell_32_io_a),
    .io_b(cell_32_io_b),
    .io_A(cell_32_io_A),
    .io_B(cell_32_io_B)
  );
  mul_cell cell_33 ( // @[mul.scala 95:35]
    .clock(cell_33_clock),
    .reset(cell_33_reset),
    .io_flush(cell_33_io_flush),
    .io_valid(cell_33_io_valid),
    .io_a_in(cell_33_io_a_in),
    .io_b_in(cell_33_io_b_in),
    .io_sum_in(cell_33_io_sum_in),
    .io_last(cell_33_io_last),
    .io_a_out(cell_33_io_a_out),
    .io_b_out(cell_33_io_b_out),
    .io_sum_out(cell_33_io_sum_out),
    .io_ready(cell_33_io_ready),
    .io_a(cell_33_io_a),
    .io_b(cell_33_io_b),
    .io_A(cell_33_io_A),
    .io_B(cell_33_io_B)
  );
  mul_cell cell_34 ( // @[mul.scala 95:35]
    .clock(cell_34_clock),
    .reset(cell_34_reset),
    .io_flush(cell_34_io_flush),
    .io_valid(cell_34_io_valid),
    .io_a_in(cell_34_io_a_in),
    .io_b_in(cell_34_io_b_in),
    .io_sum_in(cell_34_io_sum_in),
    .io_last(cell_34_io_last),
    .io_a_out(cell_34_io_a_out),
    .io_b_out(cell_34_io_b_out),
    .io_sum_out(cell_34_io_sum_out),
    .io_ready(cell_34_io_ready),
    .io_a(cell_34_io_a),
    .io_b(cell_34_io_b),
    .io_A(cell_34_io_A),
    .io_B(cell_34_io_B)
  );
  mul_cell cell_35 ( // @[mul.scala 95:35]
    .clock(cell_35_clock),
    .reset(cell_35_reset),
    .io_flush(cell_35_io_flush),
    .io_valid(cell_35_io_valid),
    .io_a_in(cell_35_io_a_in),
    .io_b_in(cell_35_io_b_in),
    .io_sum_in(cell_35_io_sum_in),
    .io_last(cell_35_io_last),
    .io_a_out(cell_35_io_a_out),
    .io_b_out(cell_35_io_b_out),
    .io_sum_out(cell_35_io_sum_out),
    .io_ready(cell_35_io_ready),
    .io_a(cell_35_io_a),
    .io_b(cell_35_io_b),
    .io_A(cell_35_io_A),
    .io_B(cell_35_io_B)
  );
  mul_cell cell_36 ( // @[mul.scala 95:35]
    .clock(cell_36_clock),
    .reset(cell_36_reset),
    .io_flush(cell_36_io_flush),
    .io_valid(cell_36_io_valid),
    .io_a_in(cell_36_io_a_in),
    .io_b_in(cell_36_io_b_in),
    .io_sum_in(cell_36_io_sum_in),
    .io_last(cell_36_io_last),
    .io_a_out(cell_36_io_a_out),
    .io_b_out(cell_36_io_b_out),
    .io_sum_out(cell_36_io_sum_out),
    .io_ready(cell_36_io_ready),
    .io_a(cell_36_io_a),
    .io_b(cell_36_io_b),
    .io_A(cell_36_io_A),
    .io_B(cell_36_io_B)
  );
  mul_cell cell_37 ( // @[mul.scala 95:35]
    .clock(cell_37_clock),
    .reset(cell_37_reset),
    .io_flush(cell_37_io_flush),
    .io_valid(cell_37_io_valid),
    .io_a_in(cell_37_io_a_in),
    .io_b_in(cell_37_io_b_in),
    .io_sum_in(cell_37_io_sum_in),
    .io_last(cell_37_io_last),
    .io_a_out(cell_37_io_a_out),
    .io_b_out(cell_37_io_b_out),
    .io_sum_out(cell_37_io_sum_out),
    .io_ready(cell_37_io_ready),
    .io_a(cell_37_io_a),
    .io_b(cell_37_io_b),
    .io_A(cell_37_io_A),
    .io_B(cell_37_io_B)
  );
  mul_cell cell_38 ( // @[mul.scala 95:35]
    .clock(cell_38_clock),
    .reset(cell_38_reset),
    .io_flush(cell_38_io_flush),
    .io_valid(cell_38_io_valid),
    .io_a_in(cell_38_io_a_in),
    .io_b_in(cell_38_io_b_in),
    .io_sum_in(cell_38_io_sum_in),
    .io_last(cell_38_io_last),
    .io_a_out(cell_38_io_a_out),
    .io_b_out(cell_38_io_b_out),
    .io_sum_out(cell_38_io_sum_out),
    .io_ready(cell_38_io_ready),
    .io_a(cell_38_io_a),
    .io_b(cell_38_io_b),
    .io_A(cell_38_io_A),
    .io_B(cell_38_io_B)
  );
  mul_cell cell_39 ( // @[mul.scala 95:35]
    .clock(cell_39_clock),
    .reset(cell_39_reset),
    .io_flush(cell_39_io_flush),
    .io_valid(cell_39_io_valid),
    .io_a_in(cell_39_io_a_in),
    .io_b_in(cell_39_io_b_in),
    .io_sum_in(cell_39_io_sum_in),
    .io_last(cell_39_io_last),
    .io_a_out(cell_39_io_a_out),
    .io_b_out(cell_39_io_b_out),
    .io_sum_out(cell_39_io_sum_out),
    .io_ready(cell_39_io_ready),
    .io_a(cell_39_io_a),
    .io_b(cell_39_io_b),
    .io_A(cell_39_io_A),
    .io_B(cell_39_io_B)
  );
  mul_cell cell_40 ( // @[mul.scala 95:35]
    .clock(cell_40_clock),
    .reset(cell_40_reset),
    .io_flush(cell_40_io_flush),
    .io_valid(cell_40_io_valid),
    .io_a_in(cell_40_io_a_in),
    .io_b_in(cell_40_io_b_in),
    .io_sum_in(cell_40_io_sum_in),
    .io_last(cell_40_io_last),
    .io_a_out(cell_40_io_a_out),
    .io_b_out(cell_40_io_b_out),
    .io_sum_out(cell_40_io_sum_out),
    .io_ready(cell_40_io_ready),
    .io_a(cell_40_io_a),
    .io_b(cell_40_io_b),
    .io_A(cell_40_io_A),
    .io_B(cell_40_io_B)
  );
  mul_cell cell_41 ( // @[mul.scala 95:35]
    .clock(cell_41_clock),
    .reset(cell_41_reset),
    .io_flush(cell_41_io_flush),
    .io_valid(cell_41_io_valid),
    .io_a_in(cell_41_io_a_in),
    .io_b_in(cell_41_io_b_in),
    .io_sum_in(cell_41_io_sum_in),
    .io_last(cell_41_io_last),
    .io_a_out(cell_41_io_a_out),
    .io_b_out(cell_41_io_b_out),
    .io_sum_out(cell_41_io_sum_out),
    .io_ready(cell_41_io_ready),
    .io_a(cell_41_io_a),
    .io_b(cell_41_io_b),
    .io_A(cell_41_io_A),
    .io_B(cell_41_io_B)
  );
  mul_cell cell_42 ( // @[mul.scala 95:35]
    .clock(cell_42_clock),
    .reset(cell_42_reset),
    .io_flush(cell_42_io_flush),
    .io_valid(cell_42_io_valid),
    .io_a_in(cell_42_io_a_in),
    .io_b_in(cell_42_io_b_in),
    .io_sum_in(cell_42_io_sum_in),
    .io_last(cell_42_io_last),
    .io_a_out(cell_42_io_a_out),
    .io_b_out(cell_42_io_b_out),
    .io_sum_out(cell_42_io_sum_out),
    .io_ready(cell_42_io_ready),
    .io_a(cell_42_io_a),
    .io_b(cell_42_io_b),
    .io_A(cell_42_io_A),
    .io_B(cell_42_io_B)
  );
  mul_cell cell_43 ( // @[mul.scala 95:35]
    .clock(cell_43_clock),
    .reset(cell_43_reset),
    .io_flush(cell_43_io_flush),
    .io_valid(cell_43_io_valid),
    .io_a_in(cell_43_io_a_in),
    .io_b_in(cell_43_io_b_in),
    .io_sum_in(cell_43_io_sum_in),
    .io_last(cell_43_io_last),
    .io_a_out(cell_43_io_a_out),
    .io_b_out(cell_43_io_b_out),
    .io_sum_out(cell_43_io_sum_out),
    .io_ready(cell_43_io_ready),
    .io_a(cell_43_io_a),
    .io_b(cell_43_io_b),
    .io_A(cell_43_io_A),
    .io_B(cell_43_io_B)
  );
  mul_cell cell_44 ( // @[mul.scala 95:35]
    .clock(cell_44_clock),
    .reset(cell_44_reset),
    .io_flush(cell_44_io_flush),
    .io_valid(cell_44_io_valid),
    .io_a_in(cell_44_io_a_in),
    .io_b_in(cell_44_io_b_in),
    .io_sum_in(cell_44_io_sum_in),
    .io_last(cell_44_io_last),
    .io_a_out(cell_44_io_a_out),
    .io_b_out(cell_44_io_b_out),
    .io_sum_out(cell_44_io_sum_out),
    .io_ready(cell_44_io_ready),
    .io_a(cell_44_io_a),
    .io_b(cell_44_io_b),
    .io_A(cell_44_io_A),
    .io_B(cell_44_io_B)
  );
  mul_cell cell_45 ( // @[mul.scala 95:35]
    .clock(cell_45_clock),
    .reset(cell_45_reset),
    .io_flush(cell_45_io_flush),
    .io_valid(cell_45_io_valid),
    .io_a_in(cell_45_io_a_in),
    .io_b_in(cell_45_io_b_in),
    .io_sum_in(cell_45_io_sum_in),
    .io_last(cell_45_io_last),
    .io_a_out(cell_45_io_a_out),
    .io_b_out(cell_45_io_b_out),
    .io_sum_out(cell_45_io_sum_out),
    .io_ready(cell_45_io_ready),
    .io_a(cell_45_io_a),
    .io_b(cell_45_io_b),
    .io_A(cell_45_io_A),
    .io_B(cell_45_io_B)
  );
  mul_cell cell_46 ( // @[mul.scala 95:35]
    .clock(cell_46_clock),
    .reset(cell_46_reset),
    .io_flush(cell_46_io_flush),
    .io_valid(cell_46_io_valid),
    .io_a_in(cell_46_io_a_in),
    .io_b_in(cell_46_io_b_in),
    .io_sum_in(cell_46_io_sum_in),
    .io_last(cell_46_io_last),
    .io_a_out(cell_46_io_a_out),
    .io_b_out(cell_46_io_b_out),
    .io_sum_out(cell_46_io_sum_out),
    .io_ready(cell_46_io_ready),
    .io_a(cell_46_io_a),
    .io_b(cell_46_io_b),
    .io_A(cell_46_io_A),
    .io_B(cell_46_io_B)
  );
  mul_cell cell_47 ( // @[mul.scala 95:35]
    .clock(cell_47_clock),
    .reset(cell_47_reset),
    .io_flush(cell_47_io_flush),
    .io_valid(cell_47_io_valid),
    .io_a_in(cell_47_io_a_in),
    .io_b_in(cell_47_io_b_in),
    .io_sum_in(cell_47_io_sum_in),
    .io_last(cell_47_io_last),
    .io_a_out(cell_47_io_a_out),
    .io_b_out(cell_47_io_b_out),
    .io_sum_out(cell_47_io_sum_out),
    .io_ready(cell_47_io_ready),
    .io_a(cell_47_io_a),
    .io_b(cell_47_io_b),
    .io_A(cell_47_io_A),
    .io_B(cell_47_io_B)
  );
  mul_cell cell_48 ( // @[mul.scala 95:35]
    .clock(cell_48_clock),
    .reset(cell_48_reset),
    .io_flush(cell_48_io_flush),
    .io_valid(cell_48_io_valid),
    .io_a_in(cell_48_io_a_in),
    .io_b_in(cell_48_io_b_in),
    .io_sum_in(cell_48_io_sum_in),
    .io_last(cell_48_io_last),
    .io_a_out(cell_48_io_a_out),
    .io_b_out(cell_48_io_b_out),
    .io_sum_out(cell_48_io_sum_out),
    .io_ready(cell_48_io_ready),
    .io_a(cell_48_io_a),
    .io_b(cell_48_io_b),
    .io_A(cell_48_io_A),
    .io_B(cell_48_io_B)
  );
  mul_cell cell_49 ( // @[mul.scala 95:35]
    .clock(cell_49_clock),
    .reset(cell_49_reset),
    .io_flush(cell_49_io_flush),
    .io_valid(cell_49_io_valid),
    .io_a_in(cell_49_io_a_in),
    .io_b_in(cell_49_io_b_in),
    .io_sum_in(cell_49_io_sum_in),
    .io_last(cell_49_io_last),
    .io_a_out(cell_49_io_a_out),
    .io_b_out(cell_49_io_b_out),
    .io_sum_out(cell_49_io_sum_out),
    .io_ready(cell_49_io_ready),
    .io_a(cell_49_io_a),
    .io_b(cell_49_io_b),
    .io_A(cell_49_io_A),
    .io_B(cell_49_io_B)
  );
  mul_cell cell_50 ( // @[mul.scala 95:35]
    .clock(cell_50_clock),
    .reset(cell_50_reset),
    .io_flush(cell_50_io_flush),
    .io_valid(cell_50_io_valid),
    .io_a_in(cell_50_io_a_in),
    .io_b_in(cell_50_io_b_in),
    .io_sum_in(cell_50_io_sum_in),
    .io_last(cell_50_io_last),
    .io_a_out(cell_50_io_a_out),
    .io_b_out(cell_50_io_b_out),
    .io_sum_out(cell_50_io_sum_out),
    .io_ready(cell_50_io_ready),
    .io_a(cell_50_io_a),
    .io_b(cell_50_io_b),
    .io_A(cell_50_io_A),
    .io_B(cell_50_io_B)
  );
  mul_cell cell_51 ( // @[mul.scala 95:35]
    .clock(cell_51_clock),
    .reset(cell_51_reset),
    .io_flush(cell_51_io_flush),
    .io_valid(cell_51_io_valid),
    .io_a_in(cell_51_io_a_in),
    .io_b_in(cell_51_io_b_in),
    .io_sum_in(cell_51_io_sum_in),
    .io_last(cell_51_io_last),
    .io_a_out(cell_51_io_a_out),
    .io_b_out(cell_51_io_b_out),
    .io_sum_out(cell_51_io_sum_out),
    .io_ready(cell_51_io_ready),
    .io_a(cell_51_io_a),
    .io_b(cell_51_io_b),
    .io_A(cell_51_io_A),
    .io_B(cell_51_io_B)
  );
  mul_cell cell_52 ( // @[mul.scala 95:35]
    .clock(cell_52_clock),
    .reset(cell_52_reset),
    .io_flush(cell_52_io_flush),
    .io_valid(cell_52_io_valid),
    .io_a_in(cell_52_io_a_in),
    .io_b_in(cell_52_io_b_in),
    .io_sum_in(cell_52_io_sum_in),
    .io_last(cell_52_io_last),
    .io_a_out(cell_52_io_a_out),
    .io_b_out(cell_52_io_b_out),
    .io_sum_out(cell_52_io_sum_out),
    .io_ready(cell_52_io_ready),
    .io_a(cell_52_io_a),
    .io_b(cell_52_io_b),
    .io_A(cell_52_io_A),
    .io_B(cell_52_io_B)
  );
  mul_cell cell_53 ( // @[mul.scala 95:35]
    .clock(cell_53_clock),
    .reset(cell_53_reset),
    .io_flush(cell_53_io_flush),
    .io_valid(cell_53_io_valid),
    .io_a_in(cell_53_io_a_in),
    .io_b_in(cell_53_io_b_in),
    .io_sum_in(cell_53_io_sum_in),
    .io_last(cell_53_io_last),
    .io_a_out(cell_53_io_a_out),
    .io_b_out(cell_53_io_b_out),
    .io_sum_out(cell_53_io_sum_out),
    .io_ready(cell_53_io_ready),
    .io_a(cell_53_io_a),
    .io_b(cell_53_io_b),
    .io_A(cell_53_io_A),
    .io_B(cell_53_io_B)
  );
  mul_cell cell_54 ( // @[mul.scala 95:35]
    .clock(cell_54_clock),
    .reset(cell_54_reset),
    .io_flush(cell_54_io_flush),
    .io_valid(cell_54_io_valid),
    .io_a_in(cell_54_io_a_in),
    .io_b_in(cell_54_io_b_in),
    .io_sum_in(cell_54_io_sum_in),
    .io_last(cell_54_io_last),
    .io_a_out(cell_54_io_a_out),
    .io_b_out(cell_54_io_b_out),
    .io_sum_out(cell_54_io_sum_out),
    .io_ready(cell_54_io_ready),
    .io_a(cell_54_io_a),
    .io_b(cell_54_io_b),
    .io_A(cell_54_io_A),
    .io_B(cell_54_io_B)
  );
  mul_cell cell_55 ( // @[mul.scala 95:35]
    .clock(cell_55_clock),
    .reset(cell_55_reset),
    .io_flush(cell_55_io_flush),
    .io_valid(cell_55_io_valid),
    .io_a_in(cell_55_io_a_in),
    .io_b_in(cell_55_io_b_in),
    .io_sum_in(cell_55_io_sum_in),
    .io_last(cell_55_io_last),
    .io_a_out(cell_55_io_a_out),
    .io_b_out(cell_55_io_b_out),
    .io_sum_out(cell_55_io_sum_out),
    .io_ready(cell_55_io_ready),
    .io_a(cell_55_io_a),
    .io_b(cell_55_io_b),
    .io_A(cell_55_io_A),
    .io_B(cell_55_io_B)
  );
  mul_cell cell_56 ( // @[mul.scala 95:35]
    .clock(cell_56_clock),
    .reset(cell_56_reset),
    .io_flush(cell_56_io_flush),
    .io_valid(cell_56_io_valid),
    .io_a_in(cell_56_io_a_in),
    .io_b_in(cell_56_io_b_in),
    .io_sum_in(cell_56_io_sum_in),
    .io_last(cell_56_io_last),
    .io_a_out(cell_56_io_a_out),
    .io_b_out(cell_56_io_b_out),
    .io_sum_out(cell_56_io_sum_out),
    .io_ready(cell_56_io_ready),
    .io_a(cell_56_io_a),
    .io_b(cell_56_io_b),
    .io_A(cell_56_io_A),
    .io_B(cell_56_io_B)
  );
  mul_cell cell_57 ( // @[mul.scala 95:35]
    .clock(cell_57_clock),
    .reset(cell_57_reset),
    .io_flush(cell_57_io_flush),
    .io_valid(cell_57_io_valid),
    .io_a_in(cell_57_io_a_in),
    .io_b_in(cell_57_io_b_in),
    .io_sum_in(cell_57_io_sum_in),
    .io_last(cell_57_io_last),
    .io_a_out(cell_57_io_a_out),
    .io_b_out(cell_57_io_b_out),
    .io_sum_out(cell_57_io_sum_out),
    .io_ready(cell_57_io_ready),
    .io_a(cell_57_io_a),
    .io_b(cell_57_io_b),
    .io_A(cell_57_io_A),
    .io_B(cell_57_io_B)
  );
  mul_cell cell_58 ( // @[mul.scala 95:35]
    .clock(cell_58_clock),
    .reset(cell_58_reset),
    .io_flush(cell_58_io_flush),
    .io_valid(cell_58_io_valid),
    .io_a_in(cell_58_io_a_in),
    .io_b_in(cell_58_io_b_in),
    .io_sum_in(cell_58_io_sum_in),
    .io_last(cell_58_io_last),
    .io_a_out(cell_58_io_a_out),
    .io_b_out(cell_58_io_b_out),
    .io_sum_out(cell_58_io_sum_out),
    .io_ready(cell_58_io_ready),
    .io_a(cell_58_io_a),
    .io_b(cell_58_io_b),
    .io_A(cell_58_io_A),
    .io_B(cell_58_io_B)
  );
  mul_cell cell_59 ( // @[mul.scala 95:35]
    .clock(cell_59_clock),
    .reset(cell_59_reset),
    .io_flush(cell_59_io_flush),
    .io_valid(cell_59_io_valid),
    .io_a_in(cell_59_io_a_in),
    .io_b_in(cell_59_io_b_in),
    .io_sum_in(cell_59_io_sum_in),
    .io_last(cell_59_io_last),
    .io_a_out(cell_59_io_a_out),
    .io_b_out(cell_59_io_b_out),
    .io_sum_out(cell_59_io_sum_out),
    .io_ready(cell_59_io_ready),
    .io_a(cell_59_io_a),
    .io_b(cell_59_io_b),
    .io_A(cell_59_io_A),
    .io_B(cell_59_io_B)
  );
  mul_cell cell_60 ( // @[mul.scala 95:35]
    .clock(cell_60_clock),
    .reset(cell_60_reset),
    .io_flush(cell_60_io_flush),
    .io_valid(cell_60_io_valid),
    .io_a_in(cell_60_io_a_in),
    .io_b_in(cell_60_io_b_in),
    .io_sum_in(cell_60_io_sum_in),
    .io_last(cell_60_io_last),
    .io_a_out(cell_60_io_a_out),
    .io_b_out(cell_60_io_b_out),
    .io_sum_out(cell_60_io_sum_out),
    .io_ready(cell_60_io_ready),
    .io_a(cell_60_io_a),
    .io_b(cell_60_io_b),
    .io_A(cell_60_io_A),
    .io_B(cell_60_io_B)
  );
  mul_cell cell_61 ( // @[mul.scala 95:35]
    .clock(cell_61_clock),
    .reset(cell_61_reset),
    .io_flush(cell_61_io_flush),
    .io_valid(cell_61_io_valid),
    .io_a_in(cell_61_io_a_in),
    .io_b_in(cell_61_io_b_in),
    .io_sum_in(cell_61_io_sum_in),
    .io_last(cell_61_io_last),
    .io_a_out(cell_61_io_a_out),
    .io_b_out(cell_61_io_b_out),
    .io_sum_out(cell_61_io_sum_out),
    .io_ready(cell_61_io_ready),
    .io_a(cell_61_io_a),
    .io_b(cell_61_io_b),
    .io_A(cell_61_io_A),
    .io_B(cell_61_io_B)
  );
  mul_cell cell_62 ( // @[mul.scala 95:35]
    .clock(cell_62_clock),
    .reset(cell_62_reset),
    .io_flush(cell_62_io_flush),
    .io_valid(cell_62_io_valid),
    .io_a_in(cell_62_io_a_in),
    .io_b_in(cell_62_io_b_in),
    .io_sum_in(cell_62_io_sum_in),
    .io_last(cell_62_io_last),
    .io_a_out(cell_62_io_a_out),
    .io_b_out(cell_62_io_b_out),
    .io_sum_out(cell_62_io_sum_out),
    .io_ready(cell_62_io_ready),
    .io_a(cell_62_io_a),
    .io_b(cell_62_io_b),
    .io_A(cell_62_io_A),
    .io_B(cell_62_io_B)
  );
  mul_cell cell_63 ( // @[mul.scala 95:35]
    .clock(cell_63_clock),
    .reset(cell_63_reset),
    .io_flush(cell_63_io_flush),
    .io_valid(cell_63_io_valid),
    .io_a_in(cell_63_io_a_in),
    .io_b_in(cell_63_io_b_in),
    .io_sum_in(cell_63_io_sum_in),
    .io_last(cell_63_io_last),
    .io_a_out(cell_63_io_a_out),
    .io_b_out(cell_63_io_b_out),
    .io_sum_out(cell_63_io_sum_out),
    .io_ready(cell_63_io_ready),
    .io_a(cell_63_io_a),
    .io_b(cell_63_io_b),
    .io_A(cell_63_io_A),
    .io_B(cell_63_io_B)
  );
  mul_cell cell_64 ( // @[mul.scala 95:35]
    .clock(cell_64_clock),
    .reset(cell_64_reset),
    .io_flush(cell_64_io_flush),
    .io_valid(cell_64_io_valid),
    .io_a_in(cell_64_io_a_in),
    .io_b_in(cell_64_io_b_in),
    .io_sum_in(cell_64_io_sum_in),
    .io_last(cell_64_io_last),
    .io_a_out(cell_64_io_a_out),
    .io_b_out(cell_64_io_b_out),
    .io_sum_out(cell_64_io_sum_out),
    .io_ready(cell_64_io_ready),
    .io_a(cell_64_io_a),
    .io_b(cell_64_io_b),
    .io_A(cell_64_io_A),
    .io_B(cell_64_io_B)
  );
  assign io_out_valid = cell_64_io_ready; // @[mul.scala 118:18]
  assign io_result_lo = cell_64_io_sum_out[63:0]; // @[mul.scala 120:41]
  assign cell_0_clock = clock;
  assign cell_0_reset = reset;
  assign cell_0_io_flush = 1'h0; // @[mul.scala 97:23]
  assign cell_0_io_valid = valid; // @[mul.scala 98:23]
  assign cell_0_io_a_in = a; // @[mul.scala 99:23]
  assign cell_0_io_b_in = b; // @[mul.scala 100:23]
  assign cell_0_io_sum_in = 129'h0; // @[mul.scala 101:23]
  assign cell_0_io_last = 1'h0; // @[mul.scala 102:23]
  assign cell_0_io_a = io_multiplicand; // @[mul.scala 103:23]
  assign cell_0_io_b = io_multiplier; // @[mul.scala 104:23]
  assign cell_1_clock = clock;
  assign cell_1_reset = reset;
  assign cell_1_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_1_io_valid = cell_0_io_ready; // @[mul.scala 108:25]
  assign cell_1_io_a_in = cell_0_io_a_out; // @[mul.scala 109:25]
  assign cell_1_io_b_in = cell_0_io_b_out; // @[mul.scala 110:25]
  assign cell_1_io_sum_in = cell_0_io_sum_out; // @[mul.scala 111:25]
  assign cell_1_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_1_io_a = cell_0_io_A; // @[mul.scala 113:25]
  assign cell_1_io_b = cell_0_io_B; // @[mul.scala 114:25]
  assign cell_2_clock = clock;
  assign cell_2_reset = reset;
  assign cell_2_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_2_io_valid = cell_1_io_ready; // @[mul.scala 108:25]
  assign cell_2_io_a_in = cell_1_io_a_out; // @[mul.scala 109:25]
  assign cell_2_io_b_in = cell_1_io_b_out; // @[mul.scala 110:25]
  assign cell_2_io_sum_in = cell_1_io_sum_out; // @[mul.scala 111:25]
  assign cell_2_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_2_io_a = cell_1_io_A; // @[mul.scala 113:25]
  assign cell_2_io_b = cell_1_io_B; // @[mul.scala 114:25]
  assign cell_3_clock = clock;
  assign cell_3_reset = reset;
  assign cell_3_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_3_io_valid = cell_2_io_ready; // @[mul.scala 108:25]
  assign cell_3_io_a_in = cell_2_io_a_out; // @[mul.scala 109:25]
  assign cell_3_io_b_in = cell_2_io_b_out; // @[mul.scala 110:25]
  assign cell_3_io_sum_in = cell_2_io_sum_out; // @[mul.scala 111:25]
  assign cell_3_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_3_io_a = cell_2_io_A; // @[mul.scala 113:25]
  assign cell_3_io_b = cell_2_io_B; // @[mul.scala 114:25]
  assign cell_4_clock = clock;
  assign cell_4_reset = reset;
  assign cell_4_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_4_io_valid = cell_3_io_ready; // @[mul.scala 108:25]
  assign cell_4_io_a_in = cell_3_io_a_out; // @[mul.scala 109:25]
  assign cell_4_io_b_in = cell_3_io_b_out; // @[mul.scala 110:25]
  assign cell_4_io_sum_in = cell_3_io_sum_out; // @[mul.scala 111:25]
  assign cell_4_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_4_io_a = cell_3_io_A; // @[mul.scala 113:25]
  assign cell_4_io_b = cell_3_io_B; // @[mul.scala 114:25]
  assign cell_5_clock = clock;
  assign cell_5_reset = reset;
  assign cell_5_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_5_io_valid = cell_4_io_ready; // @[mul.scala 108:25]
  assign cell_5_io_a_in = cell_4_io_a_out; // @[mul.scala 109:25]
  assign cell_5_io_b_in = cell_4_io_b_out; // @[mul.scala 110:25]
  assign cell_5_io_sum_in = cell_4_io_sum_out; // @[mul.scala 111:25]
  assign cell_5_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_5_io_a = cell_4_io_A; // @[mul.scala 113:25]
  assign cell_5_io_b = cell_4_io_B; // @[mul.scala 114:25]
  assign cell_6_clock = clock;
  assign cell_6_reset = reset;
  assign cell_6_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_6_io_valid = cell_5_io_ready; // @[mul.scala 108:25]
  assign cell_6_io_a_in = cell_5_io_a_out; // @[mul.scala 109:25]
  assign cell_6_io_b_in = cell_5_io_b_out; // @[mul.scala 110:25]
  assign cell_6_io_sum_in = cell_5_io_sum_out; // @[mul.scala 111:25]
  assign cell_6_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_6_io_a = cell_5_io_A; // @[mul.scala 113:25]
  assign cell_6_io_b = cell_5_io_B; // @[mul.scala 114:25]
  assign cell_7_clock = clock;
  assign cell_7_reset = reset;
  assign cell_7_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_7_io_valid = cell_6_io_ready; // @[mul.scala 108:25]
  assign cell_7_io_a_in = cell_6_io_a_out; // @[mul.scala 109:25]
  assign cell_7_io_b_in = cell_6_io_b_out; // @[mul.scala 110:25]
  assign cell_7_io_sum_in = cell_6_io_sum_out; // @[mul.scala 111:25]
  assign cell_7_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_7_io_a = cell_6_io_A; // @[mul.scala 113:25]
  assign cell_7_io_b = cell_6_io_B; // @[mul.scala 114:25]
  assign cell_8_clock = clock;
  assign cell_8_reset = reset;
  assign cell_8_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_8_io_valid = cell_7_io_ready; // @[mul.scala 108:25]
  assign cell_8_io_a_in = cell_7_io_a_out; // @[mul.scala 109:25]
  assign cell_8_io_b_in = cell_7_io_b_out; // @[mul.scala 110:25]
  assign cell_8_io_sum_in = cell_7_io_sum_out; // @[mul.scala 111:25]
  assign cell_8_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_8_io_a = cell_7_io_A; // @[mul.scala 113:25]
  assign cell_8_io_b = cell_7_io_B; // @[mul.scala 114:25]
  assign cell_9_clock = clock;
  assign cell_9_reset = reset;
  assign cell_9_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_9_io_valid = cell_8_io_ready; // @[mul.scala 108:25]
  assign cell_9_io_a_in = cell_8_io_a_out; // @[mul.scala 109:25]
  assign cell_9_io_b_in = cell_8_io_b_out; // @[mul.scala 110:25]
  assign cell_9_io_sum_in = cell_8_io_sum_out; // @[mul.scala 111:25]
  assign cell_9_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_9_io_a = cell_8_io_A; // @[mul.scala 113:25]
  assign cell_9_io_b = cell_8_io_B; // @[mul.scala 114:25]
  assign cell_10_clock = clock;
  assign cell_10_reset = reset;
  assign cell_10_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_10_io_valid = cell_9_io_ready; // @[mul.scala 108:25]
  assign cell_10_io_a_in = cell_9_io_a_out; // @[mul.scala 109:25]
  assign cell_10_io_b_in = cell_9_io_b_out; // @[mul.scala 110:25]
  assign cell_10_io_sum_in = cell_9_io_sum_out; // @[mul.scala 111:25]
  assign cell_10_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_10_io_a = cell_9_io_A; // @[mul.scala 113:25]
  assign cell_10_io_b = cell_9_io_B; // @[mul.scala 114:25]
  assign cell_11_clock = clock;
  assign cell_11_reset = reset;
  assign cell_11_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_11_io_valid = cell_10_io_ready; // @[mul.scala 108:25]
  assign cell_11_io_a_in = cell_10_io_a_out; // @[mul.scala 109:25]
  assign cell_11_io_b_in = cell_10_io_b_out; // @[mul.scala 110:25]
  assign cell_11_io_sum_in = cell_10_io_sum_out; // @[mul.scala 111:25]
  assign cell_11_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_11_io_a = cell_10_io_A; // @[mul.scala 113:25]
  assign cell_11_io_b = cell_10_io_B; // @[mul.scala 114:25]
  assign cell_12_clock = clock;
  assign cell_12_reset = reset;
  assign cell_12_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_12_io_valid = cell_11_io_ready; // @[mul.scala 108:25]
  assign cell_12_io_a_in = cell_11_io_a_out; // @[mul.scala 109:25]
  assign cell_12_io_b_in = cell_11_io_b_out; // @[mul.scala 110:25]
  assign cell_12_io_sum_in = cell_11_io_sum_out; // @[mul.scala 111:25]
  assign cell_12_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_12_io_a = cell_11_io_A; // @[mul.scala 113:25]
  assign cell_12_io_b = cell_11_io_B; // @[mul.scala 114:25]
  assign cell_13_clock = clock;
  assign cell_13_reset = reset;
  assign cell_13_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_13_io_valid = cell_12_io_ready; // @[mul.scala 108:25]
  assign cell_13_io_a_in = cell_12_io_a_out; // @[mul.scala 109:25]
  assign cell_13_io_b_in = cell_12_io_b_out; // @[mul.scala 110:25]
  assign cell_13_io_sum_in = cell_12_io_sum_out; // @[mul.scala 111:25]
  assign cell_13_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_13_io_a = cell_12_io_A; // @[mul.scala 113:25]
  assign cell_13_io_b = cell_12_io_B; // @[mul.scala 114:25]
  assign cell_14_clock = clock;
  assign cell_14_reset = reset;
  assign cell_14_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_14_io_valid = cell_13_io_ready; // @[mul.scala 108:25]
  assign cell_14_io_a_in = cell_13_io_a_out; // @[mul.scala 109:25]
  assign cell_14_io_b_in = cell_13_io_b_out; // @[mul.scala 110:25]
  assign cell_14_io_sum_in = cell_13_io_sum_out; // @[mul.scala 111:25]
  assign cell_14_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_14_io_a = cell_13_io_A; // @[mul.scala 113:25]
  assign cell_14_io_b = cell_13_io_B; // @[mul.scala 114:25]
  assign cell_15_clock = clock;
  assign cell_15_reset = reset;
  assign cell_15_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_15_io_valid = cell_14_io_ready; // @[mul.scala 108:25]
  assign cell_15_io_a_in = cell_14_io_a_out; // @[mul.scala 109:25]
  assign cell_15_io_b_in = cell_14_io_b_out; // @[mul.scala 110:25]
  assign cell_15_io_sum_in = cell_14_io_sum_out; // @[mul.scala 111:25]
  assign cell_15_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_15_io_a = cell_14_io_A; // @[mul.scala 113:25]
  assign cell_15_io_b = cell_14_io_B; // @[mul.scala 114:25]
  assign cell_16_clock = clock;
  assign cell_16_reset = reset;
  assign cell_16_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_16_io_valid = cell_15_io_ready; // @[mul.scala 108:25]
  assign cell_16_io_a_in = cell_15_io_a_out; // @[mul.scala 109:25]
  assign cell_16_io_b_in = cell_15_io_b_out; // @[mul.scala 110:25]
  assign cell_16_io_sum_in = cell_15_io_sum_out; // @[mul.scala 111:25]
  assign cell_16_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_16_io_a = cell_15_io_A; // @[mul.scala 113:25]
  assign cell_16_io_b = cell_15_io_B; // @[mul.scala 114:25]
  assign cell_17_clock = clock;
  assign cell_17_reset = reset;
  assign cell_17_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_17_io_valid = cell_16_io_ready; // @[mul.scala 108:25]
  assign cell_17_io_a_in = cell_16_io_a_out; // @[mul.scala 109:25]
  assign cell_17_io_b_in = cell_16_io_b_out; // @[mul.scala 110:25]
  assign cell_17_io_sum_in = cell_16_io_sum_out; // @[mul.scala 111:25]
  assign cell_17_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_17_io_a = cell_16_io_A; // @[mul.scala 113:25]
  assign cell_17_io_b = cell_16_io_B; // @[mul.scala 114:25]
  assign cell_18_clock = clock;
  assign cell_18_reset = reset;
  assign cell_18_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_18_io_valid = cell_17_io_ready; // @[mul.scala 108:25]
  assign cell_18_io_a_in = cell_17_io_a_out; // @[mul.scala 109:25]
  assign cell_18_io_b_in = cell_17_io_b_out; // @[mul.scala 110:25]
  assign cell_18_io_sum_in = cell_17_io_sum_out; // @[mul.scala 111:25]
  assign cell_18_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_18_io_a = cell_17_io_A; // @[mul.scala 113:25]
  assign cell_18_io_b = cell_17_io_B; // @[mul.scala 114:25]
  assign cell_19_clock = clock;
  assign cell_19_reset = reset;
  assign cell_19_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_19_io_valid = cell_18_io_ready; // @[mul.scala 108:25]
  assign cell_19_io_a_in = cell_18_io_a_out; // @[mul.scala 109:25]
  assign cell_19_io_b_in = cell_18_io_b_out; // @[mul.scala 110:25]
  assign cell_19_io_sum_in = cell_18_io_sum_out; // @[mul.scala 111:25]
  assign cell_19_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_19_io_a = cell_18_io_A; // @[mul.scala 113:25]
  assign cell_19_io_b = cell_18_io_B; // @[mul.scala 114:25]
  assign cell_20_clock = clock;
  assign cell_20_reset = reset;
  assign cell_20_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_20_io_valid = cell_19_io_ready; // @[mul.scala 108:25]
  assign cell_20_io_a_in = cell_19_io_a_out; // @[mul.scala 109:25]
  assign cell_20_io_b_in = cell_19_io_b_out; // @[mul.scala 110:25]
  assign cell_20_io_sum_in = cell_19_io_sum_out; // @[mul.scala 111:25]
  assign cell_20_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_20_io_a = cell_19_io_A; // @[mul.scala 113:25]
  assign cell_20_io_b = cell_19_io_B; // @[mul.scala 114:25]
  assign cell_21_clock = clock;
  assign cell_21_reset = reset;
  assign cell_21_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_21_io_valid = cell_20_io_ready; // @[mul.scala 108:25]
  assign cell_21_io_a_in = cell_20_io_a_out; // @[mul.scala 109:25]
  assign cell_21_io_b_in = cell_20_io_b_out; // @[mul.scala 110:25]
  assign cell_21_io_sum_in = cell_20_io_sum_out; // @[mul.scala 111:25]
  assign cell_21_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_21_io_a = cell_20_io_A; // @[mul.scala 113:25]
  assign cell_21_io_b = cell_20_io_B; // @[mul.scala 114:25]
  assign cell_22_clock = clock;
  assign cell_22_reset = reset;
  assign cell_22_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_22_io_valid = cell_21_io_ready; // @[mul.scala 108:25]
  assign cell_22_io_a_in = cell_21_io_a_out; // @[mul.scala 109:25]
  assign cell_22_io_b_in = cell_21_io_b_out; // @[mul.scala 110:25]
  assign cell_22_io_sum_in = cell_21_io_sum_out; // @[mul.scala 111:25]
  assign cell_22_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_22_io_a = cell_21_io_A; // @[mul.scala 113:25]
  assign cell_22_io_b = cell_21_io_B; // @[mul.scala 114:25]
  assign cell_23_clock = clock;
  assign cell_23_reset = reset;
  assign cell_23_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_23_io_valid = cell_22_io_ready; // @[mul.scala 108:25]
  assign cell_23_io_a_in = cell_22_io_a_out; // @[mul.scala 109:25]
  assign cell_23_io_b_in = cell_22_io_b_out; // @[mul.scala 110:25]
  assign cell_23_io_sum_in = cell_22_io_sum_out; // @[mul.scala 111:25]
  assign cell_23_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_23_io_a = cell_22_io_A; // @[mul.scala 113:25]
  assign cell_23_io_b = cell_22_io_B; // @[mul.scala 114:25]
  assign cell_24_clock = clock;
  assign cell_24_reset = reset;
  assign cell_24_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_24_io_valid = cell_23_io_ready; // @[mul.scala 108:25]
  assign cell_24_io_a_in = cell_23_io_a_out; // @[mul.scala 109:25]
  assign cell_24_io_b_in = cell_23_io_b_out; // @[mul.scala 110:25]
  assign cell_24_io_sum_in = cell_23_io_sum_out; // @[mul.scala 111:25]
  assign cell_24_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_24_io_a = cell_23_io_A; // @[mul.scala 113:25]
  assign cell_24_io_b = cell_23_io_B; // @[mul.scala 114:25]
  assign cell_25_clock = clock;
  assign cell_25_reset = reset;
  assign cell_25_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_25_io_valid = cell_24_io_ready; // @[mul.scala 108:25]
  assign cell_25_io_a_in = cell_24_io_a_out; // @[mul.scala 109:25]
  assign cell_25_io_b_in = cell_24_io_b_out; // @[mul.scala 110:25]
  assign cell_25_io_sum_in = cell_24_io_sum_out; // @[mul.scala 111:25]
  assign cell_25_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_25_io_a = cell_24_io_A; // @[mul.scala 113:25]
  assign cell_25_io_b = cell_24_io_B; // @[mul.scala 114:25]
  assign cell_26_clock = clock;
  assign cell_26_reset = reset;
  assign cell_26_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_26_io_valid = cell_25_io_ready; // @[mul.scala 108:25]
  assign cell_26_io_a_in = cell_25_io_a_out; // @[mul.scala 109:25]
  assign cell_26_io_b_in = cell_25_io_b_out; // @[mul.scala 110:25]
  assign cell_26_io_sum_in = cell_25_io_sum_out; // @[mul.scala 111:25]
  assign cell_26_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_26_io_a = cell_25_io_A; // @[mul.scala 113:25]
  assign cell_26_io_b = cell_25_io_B; // @[mul.scala 114:25]
  assign cell_27_clock = clock;
  assign cell_27_reset = reset;
  assign cell_27_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_27_io_valid = cell_26_io_ready; // @[mul.scala 108:25]
  assign cell_27_io_a_in = cell_26_io_a_out; // @[mul.scala 109:25]
  assign cell_27_io_b_in = cell_26_io_b_out; // @[mul.scala 110:25]
  assign cell_27_io_sum_in = cell_26_io_sum_out; // @[mul.scala 111:25]
  assign cell_27_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_27_io_a = cell_26_io_A; // @[mul.scala 113:25]
  assign cell_27_io_b = cell_26_io_B; // @[mul.scala 114:25]
  assign cell_28_clock = clock;
  assign cell_28_reset = reset;
  assign cell_28_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_28_io_valid = cell_27_io_ready; // @[mul.scala 108:25]
  assign cell_28_io_a_in = cell_27_io_a_out; // @[mul.scala 109:25]
  assign cell_28_io_b_in = cell_27_io_b_out; // @[mul.scala 110:25]
  assign cell_28_io_sum_in = cell_27_io_sum_out; // @[mul.scala 111:25]
  assign cell_28_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_28_io_a = cell_27_io_A; // @[mul.scala 113:25]
  assign cell_28_io_b = cell_27_io_B; // @[mul.scala 114:25]
  assign cell_29_clock = clock;
  assign cell_29_reset = reset;
  assign cell_29_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_29_io_valid = cell_28_io_ready; // @[mul.scala 108:25]
  assign cell_29_io_a_in = cell_28_io_a_out; // @[mul.scala 109:25]
  assign cell_29_io_b_in = cell_28_io_b_out; // @[mul.scala 110:25]
  assign cell_29_io_sum_in = cell_28_io_sum_out; // @[mul.scala 111:25]
  assign cell_29_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_29_io_a = cell_28_io_A; // @[mul.scala 113:25]
  assign cell_29_io_b = cell_28_io_B; // @[mul.scala 114:25]
  assign cell_30_clock = clock;
  assign cell_30_reset = reset;
  assign cell_30_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_30_io_valid = cell_29_io_ready; // @[mul.scala 108:25]
  assign cell_30_io_a_in = cell_29_io_a_out; // @[mul.scala 109:25]
  assign cell_30_io_b_in = cell_29_io_b_out; // @[mul.scala 110:25]
  assign cell_30_io_sum_in = cell_29_io_sum_out; // @[mul.scala 111:25]
  assign cell_30_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_30_io_a = cell_29_io_A; // @[mul.scala 113:25]
  assign cell_30_io_b = cell_29_io_B; // @[mul.scala 114:25]
  assign cell_31_clock = clock;
  assign cell_31_reset = reset;
  assign cell_31_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_31_io_valid = cell_30_io_ready; // @[mul.scala 108:25]
  assign cell_31_io_a_in = cell_30_io_a_out; // @[mul.scala 109:25]
  assign cell_31_io_b_in = cell_30_io_b_out; // @[mul.scala 110:25]
  assign cell_31_io_sum_in = cell_30_io_sum_out; // @[mul.scala 111:25]
  assign cell_31_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_31_io_a = cell_30_io_A; // @[mul.scala 113:25]
  assign cell_31_io_b = cell_30_io_B; // @[mul.scala 114:25]
  assign cell_32_clock = clock;
  assign cell_32_reset = reset;
  assign cell_32_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_32_io_valid = cell_31_io_ready; // @[mul.scala 108:25]
  assign cell_32_io_a_in = cell_31_io_a_out; // @[mul.scala 109:25]
  assign cell_32_io_b_in = cell_31_io_b_out; // @[mul.scala 110:25]
  assign cell_32_io_sum_in = cell_31_io_sum_out; // @[mul.scala 111:25]
  assign cell_32_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_32_io_a = cell_31_io_A; // @[mul.scala 113:25]
  assign cell_32_io_b = cell_31_io_B; // @[mul.scala 114:25]
  assign cell_33_clock = clock;
  assign cell_33_reset = reset;
  assign cell_33_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_33_io_valid = cell_32_io_ready; // @[mul.scala 108:25]
  assign cell_33_io_a_in = cell_32_io_a_out; // @[mul.scala 109:25]
  assign cell_33_io_b_in = cell_32_io_b_out; // @[mul.scala 110:25]
  assign cell_33_io_sum_in = cell_32_io_sum_out; // @[mul.scala 111:25]
  assign cell_33_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_33_io_a = cell_32_io_A; // @[mul.scala 113:25]
  assign cell_33_io_b = cell_32_io_B; // @[mul.scala 114:25]
  assign cell_34_clock = clock;
  assign cell_34_reset = reset;
  assign cell_34_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_34_io_valid = cell_33_io_ready; // @[mul.scala 108:25]
  assign cell_34_io_a_in = cell_33_io_a_out; // @[mul.scala 109:25]
  assign cell_34_io_b_in = cell_33_io_b_out; // @[mul.scala 110:25]
  assign cell_34_io_sum_in = cell_33_io_sum_out; // @[mul.scala 111:25]
  assign cell_34_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_34_io_a = cell_33_io_A; // @[mul.scala 113:25]
  assign cell_34_io_b = cell_33_io_B; // @[mul.scala 114:25]
  assign cell_35_clock = clock;
  assign cell_35_reset = reset;
  assign cell_35_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_35_io_valid = cell_34_io_ready; // @[mul.scala 108:25]
  assign cell_35_io_a_in = cell_34_io_a_out; // @[mul.scala 109:25]
  assign cell_35_io_b_in = cell_34_io_b_out; // @[mul.scala 110:25]
  assign cell_35_io_sum_in = cell_34_io_sum_out; // @[mul.scala 111:25]
  assign cell_35_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_35_io_a = cell_34_io_A; // @[mul.scala 113:25]
  assign cell_35_io_b = cell_34_io_B; // @[mul.scala 114:25]
  assign cell_36_clock = clock;
  assign cell_36_reset = reset;
  assign cell_36_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_36_io_valid = cell_35_io_ready; // @[mul.scala 108:25]
  assign cell_36_io_a_in = cell_35_io_a_out; // @[mul.scala 109:25]
  assign cell_36_io_b_in = cell_35_io_b_out; // @[mul.scala 110:25]
  assign cell_36_io_sum_in = cell_35_io_sum_out; // @[mul.scala 111:25]
  assign cell_36_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_36_io_a = cell_35_io_A; // @[mul.scala 113:25]
  assign cell_36_io_b = cell_35_io_B; // @[mul.scala 114:25]
  assign cell_37_clock = clock;
  assign cell_37_reset = reset;
  assign cell_37_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_37_io_valid = cell_36_io_ready; // @[mul.scala 108:25]
  assign cell_37_io_a_in = cell_36_io_a_out; // @[mul.scala 109:25]
  assign cell_37_io_b_in = cell_36_io_b_out; // @[mul.scala 110:25]
  assign cell_37_io_sum_in = cell_36_io_sum_out; // @[mul.scala 111:25]
  assign cell_37_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_37_io_a = cell_36_io_A; // @[mul.scala 113:25]
  assign cell_37_io_b = cell_36_io_B; // @[mul.scala 114:25]
  assign cell_38_clock = clock;
  assign cell_38_reset = reset;
  assign cell_38_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_38_io_valid = cell_37_io_ready; // @[mul.scala 108:25]
  assign cell_38_io_a_in = cell_37_io_a_out; // @[mul.scala 109:25]
  assign cell_38_io_b_in = cell_37_io_b_out; // @[mul.scala 110:25]
  assign cell_38_io_sum_in = cell_37_io_sum_out; // @[mul.scala 111:25]
  assign cell_38_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_38_io_a = cell_37_io_A; // @[mul.scala 113:25]
  assign cell_38_io_b = cell_37_io_B; // @[mul.scala 114:25]
  assign cell_39_clock = clock;
  assign cell_39_reset = reset;
  assign cell_39_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_39_io_valid = cell_38_io_ready; // @[mul.scala 108:25]
  assign cell_39_io_a_in = cell_38_io_a_out; // @[mul.scala 109:25]
  assign cell_39_io_b_in = cell_38_io_b_out; // @[mul.scala 110:25]
  assign cell_39_io_sum_in = cell_38_io_sum_out; // @[mul.scala 111:25]
  assign cell_39_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_39_io_a = cell_38_io_A; // @[mul.scala 113:25]
  assign cell_39_io_b = cell_38_io_B; // @[mul.scala 114:25]
  assign cell_40_clock = clock;
  assign cell_40_reset = reset;
  assign cell_40_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_40_io_valid = cell_39_io_ready; // @[mul.scala 108:25]
  assign cell_40_io_a_in = cell_39_io_a_out; // @[mul.scala 109:25]
  assign cell_40_io_b_in = cell_39_io_b_out; // @[mul.scala 110:25]
  assign cell_40_io_sum_in = cell_39_io_sum_out; // @[mul.scala 111:25]
  assign cell_40_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_40_io_a = cell_39_io_A; // @[mul.scala 113:25]
  assign cell_40_io_b = cell_39_io_B; // @[mul.scala 114:25]
  assign cell_41_clock = clock;
  assign cell_41_reset = reset;
  assign cell_41_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_41_io_valid = cell_40_io_ready; // @[mul.scala 108:25]
  assign cell_41_io_a_in = cell_40_io_a_out; // @[mul.scala 109:25]
  assign cell_41_io_b_in = cell_40_io_b_out; // @[mul.scala 110:25]
  assign cell_41_io_sum_in = cell_40_io_sum_out; // @[mul.scala 111:25]
  assign cell_41_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_41_io_a = cell_40_io_A; // @[mul.scala 113:25]
  assign cell_41_io_b = cell_40_io_B; // @[mul.scala 114:25]
  assign cell_42_clock = clock;
  assign cell_42_reset = reset;
  assign cell_42_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_42_io_valid = cell_41_io_ready; // @[mul.scala 108:25]
  assign cell_42_io_a_in = cell_41_io_a_out; // @[mul.scala 109:25]
  assign cell_42_io_b_in = cell_41_io_b_out; // @[mul.scala 110:25]
  assign cell_42_io_sum_in = cell_41_io_sum_out; // @[mul.scala 111:25]
  assign cell_42_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_42_io_a = cell_41_io_A; // @[mul.scala 113:25]
  assign cell_42_io_b = cell_41_io_B; // @[mul.scala 114:25]
  assign cell_43_clock = clock;
  assign cell_43_reset = reset;
  assign cell_43_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_43_io_valid = cell_42_io_ready; // @[mul.scala 108:25]
  assign cell_43_io_a_in = cell_42_io_a_out; // @[mul.scala 109:25]
  assign cell_43_io_b_in = cell_42_io_b_out; // @[mul.scala 110:25]
  assign cell_43_io_sum_in = cell_42_io_sum_out; // @[mul.scala 111:25]
  assign cell_43_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_43_io_a = cell_42_io_A; // @[mul.scala 113:25]
  assign cell_43_io_b = cell_42_io_B; // @[mul.scala 114:25]
  assign cell_44_clock = clock;
  assign cell_44_reset = reset;
  assign cell_44_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_44_io_valid = cell_43_io_ready; // @[mul.scala 108:25]
  assign cell_44_io_a_in = cell_43_io_a_out; // @[mul.scala 109:25]
  assign cell_44_io_b_in = cell_43_io_b_out; // @[mul.scala 110:25]
  assign cell_44_io_sum_in = cell_43_io_sum_out; // @[mul.scala 111:25]
  assign cell_44_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_44_io_a = cell_43_io_A; // @[mul.scala 113:25]
  assign cell_44_io_b = cell_43_io_B; // @[mul.scala 114:25]
  assign cell_45_clock = clock;
  assign cell_45_reset = reset;
  assign cell_45_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_45_io_valid = cell_44_io_ready; // @[mul.scala 108:25]
  assign cell_45_io_a_in = cell_44_io_a_out; // @[mul.scala 109:25]
  assign cell_45_io_b_in = cell_44_io_b_out; // @[mul.scala 110:25]
  assign cell_45_io_sum_in = cell_44_io_sum_out; // @[mul.scala 111:25]
  assign cell_45_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_45_io_a = cell_44_io_A; // @[mul.scala 113:25]
  assign cell_45_io_b = cell_44_io_B; // @[mul.scala 114:25]
  assign cell_46_clock = clock;
  assign cell_46_reset = reset;
  assign cell_46_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_46_io_valid = cell_45_io_ready; // @[mul.scala 108:25]
  assign cell_46_io_a_in = cell_45_io_a_out; // @[mul.scala 109:25]
  assign cell_46_io_b_in = cell_45_io_b_out; // @[mul.scala 110:25]
  assign cell_46_io_sum_in = cell_45_io_sum_out; // @[mul.scala 111:25]
  assign cell_46_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_46_io_a = cell_45_io_A; // @[mul.scala 113:25]
  assign cell_46_io_b = cell_45_io_B; // @[mul.scala 114:25]
  assign cell_47_clock = clock;
  assign cell_47_reset = reset;
  assign cell_47_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_47_io_valid = cell_46_io_ready; // @[mul.scala 108:25]
  assign cell_47_io_a_in = cell_46_io_a_out; // @[mul.scala 109:25]
  assign cell_47_io_b_in = cell_46_io_b_out; // @[mul.scala 110:25]
  assign cell_47_io_sum_in = cell_46_io_sum_out; // @[mul.scala 111:25]
  assign cell_47_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_47_io_a = cell_46_io_A; // @[mul.scala 113:25]
  assign cell_47_io_b = cell_46_io_B; // @[mul.scala 114:25]
  assign cell_48_clock = clock;
  assign cell_48_reset = reset;
  assign cell_48_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_48_io_valid = cell_47_io_ready; // @[mul.scala 108:25]
  assign cell_48_io_a_in = cell_47_io_a_out; // @[mul.scala 109:25]
  assign cell_48_io_b_in = cell_47_io_b_out; // @[mul.scala 110:25]
  assign cell_48_io_sum_in = cell_47_io_sum_out; // @[mul.scala 111:25]
  assign cell_48_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_48_io_a = cell_47_io_A; // @[mul.scala 113:25]
  assign cell_48_io_b = cell_47_io_B; // @[mul.scala 114:25]
  assign cell_49_clock = clock;
  assign cell_49_reset = reset;
  assign cell_49_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_49_io_valid = cell_48_io_ready; // @[mul.scala 108:25]
  assign cell_49_io_a_in = cell_48_io_a_out; // @[mul.scala 109:25]
  assign cell_49_io_b_in = cell_48_io_b_out; // @[mul.scala 110:25]
  assign cell_49_io_sum_in = cell_48_io_sum_out; // @[mul.scala 111:25]
  assign cell_49_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_49_io_a = cell_48_io_A; // @[mul.scala 113:25]
  assign cell_49_io_b = cell_48_io_B; // @[mul.scala 114:25]
  assign cell_50_clock = clock;
  assign cell_50_reset = reset;
  assign cell_50_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_50_io_valid = cell_49_io_ready; // @[mul.scala 108:25]
  assign cell_50_io_a_in = cell_49_io_a_out; // @[mul.scala 109:25]
  assign cell_50_io_b_in = cell_49_io_b_out; // @[mul.scala 110:25]
  assign cell_50_io_sum_in = cell_49_io_sum_out; // @[mul.scala 111:25]
  assign cell_50_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_50_io_a = cell_49_io_A; // @[mul.scala 113:25]
  assign cell_50_io_b = cell_49_io_B; // @[mul.scala 114:25]
  assign cell_51_clock = clock;
  assign cell_51_reset = reset;
  assign cell_51_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_51_io_valid = cell_50_io_ready; // @[mul.scala 108:25]
  assign cell_51_io_a_in = cell_50_io_a_out; // @[mul.scala 109:25]
  assign cell_51_io_b_in = cell_50_io_b_out; // @[mul.scala 110:25]
  assign cell_51_io_sum_in = cell_50_io_sum_out; // @[mul.scala 111:25]
  assign cell_51_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_51_io_a = cell_50_io_A; // @[mul.scala 113:25]
  assign cell_51_io_b = cell_50_io_B; // @[mul.scala 114:25]
  assign cell_52_clock = clock;
  assign cell_52_reset = reset;
  assign cell_52_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_52_io_valid = cell_51_io_ready; // @[mul.scala 108:25]
  assign cell_52_io_a_in = cell_51_io_a_out; // @[mul.scala 109:25]
  assign cell_52_io_b_in = cell_51_io_b_out; // @[mul.scala 110:25]
  assign cell_52_io_sum_in = cell_51_io_sum_out; // @[mul.scala 111:25]
  assign cell_52_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_52_io_a = cell_51_io_A; // @[mul.scala 113:25]
  assign cell_52_io_b = cell_51_io_B; // @[mul.scala 114:25]
  assign cell_53_clock = clock;
  assign cell_53_reset = reset;
  assign cell_53_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_53_io_valid = cell_52_io_ready; // @[mul.scala 108:25]
  assign cell_53_io_a_in = cell_52_io_a_out; // @[mul.scala 109:25]
  assign cell_53_io_b_in = cell_52_io_b_out; // @[mul.scala 110:25]
  assign cell_53_io_sum_in = cell_52_io_sum_out; // @[mul.scala 111:25]
  assign cell_53_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_53_io_a = cell_52_io_A; // @[mul.scala 113:25]
  assign cell_53_io_b = cell_52_io_B; // @[mul.scala 114:25]
  assign cell_54_clock = clock;
  assign cell_54_reset = reset;
  assign cell_54_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_54_io_valid = cell_53_io_ready; // @[mul.scala 108:25]
  assign cell_54_io_a_in = cell_53_io_a_out; // @[mul.scala 109:25]
  assign cell_54_io_b_in = cell_53_io_b_out; // @[mul.scala 110:25]
  assign cell_54_io_sum_in = cell_53_io_sum_out; // @[mul.scala 111:25]
  assign cell_54_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_54_io_a = cell_53_io_A; // @[mul.scala 113:25]
  assign cell_54_io_b = cell_53_io_B; // @[mul.scala 114:25]
  assign cell_55_clock = clock;
  assign cell_55_reset = reset;
  assign cell_55_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_55_io_valid = cell_54_io_ready; // @[mul.scala 108:25]
  assign cell_55_io_a_in = cell_54_io_a_out; // @[mul.scala 109:25]
  assign cell_55_io_b_in = cell_54_io_b_out; // @[mul.scala 110:25]
  assign cell_55_io_sum_in = cell_54_io_sum_out; // @[mul.scala 111:25]
  assign cell_55_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_55_io_a = cell_54_io_A; // @[mul.scala 113:25]
  assign cell_55_io_b = cell_54_io_B; // @[mul.scala 114:25]
  assign cell_56_clock = clock;
  assign cell_56_reset = reset;
  assign cell_56_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_56_io_valid = cell_55_io_ready; // @[mul.scala 108:25]
  assign cell_56_io_a_in = cell_55_io_a_out; // @[mul.scala 109:25]
  assign cell_56_io_b_in = cell_55_io_b_out; // @[mul.scala 110:25]
  assign cell_56_io_sum_in = cell_55_io_sum_out; // @[mul.scala 111:25]
  assign cell_56_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_56_io_a = cell_55_io_A; // @[mul.scala 113:25]
  assign cell_56_io_b = cell_55_io_B; // @[mul.scala 114:25]
  assign cell_57_clock = clock;
  assign cell_57_reset = reset;
  assign cell_57_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_57_io_valid = cell_56_io_ready; // @[mul.scala 108:25]
  assign cell_57_io_a_in = cell_56_io_a_out; // @[mul.scala 109:25]
  assign cell_57_io_b_in = cell_56_io_b_out; // @[mul.scala 110:25]
  assign cell_57_io_sum_in = cell_56_io_sum_out; // @[mul.scala 111:25]
  assign cell_57_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_57_io_a = cell_56_io_A; // @[mul.scala 113:25]
  assign cell_57_io_b = cell_56_io_B; // @[mul.scala 114:25]
  assign cell_58_clock = clock;
  assign cell_58_reset = reset;
  assign cell_58_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_58_io_valid = cell_57_io_ready; // @[mul.scala 108:25]
  assign cell_58_io_a_in = cell_57_io_a_out; // @[mul.scala 109:25]
  assign cell_58_io_b_in = cell_57_io_b_out; // @[mul.scala 110:25]
  assign cell_58_io_sum_in = cell_57_io_sum_out; // @[mul.scala 111:25]
  assign cell_58_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_58_io_a = cell_57_io_A; // @[mul.scala 113:25]
  assign cell_58_io_b = cell_57_io_B; // @[mul.scala 114:25]
  assign cell_59_clock = clock;
  assign cell_59_reset = reset;
  assign cell_59_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_59_io_valid = cell_58_io_ready; // @[mul.scala 108:25]
  assign cell_59_io_a_in = cell_58_io_a_out; // @[mul.scala 109:25]
  assign cell_59_io_b_in = cell_58_io_b_out; // @[mul.scala 110:25]
  assign cell_59_io_sum_in = cell_58_io_sum_out; // @[mul.scala 111:25]
  assign cell_59_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_59_io_a = cell_58_io_A; // @[mul.scala 113:25]
  assign cell_59_io_b = cell_58_io_B; // @[mul.scala 114:25]
  assign cell_60_clock = clock;
  assign cell_60_reset = reset;
  assign cell_60_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_60_io_valid = cell_59_io_ready; // @[mul.scala 108:25]
  assign cell_60_io_a_in = cell_59_io_a_out; // @[mul.scala 109:25]
  assign cell_60_io_b_in = cell_59_io_b_out; // @[mul.scala 110:25]
  assign cell_60_io_sum_in = cell_59_io_sum_out; // @[mul.scala 111:25]
  assign cell_60_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_60_io_a = cell_59_io_A; // @[mul.scala 113:25]
  assign cell_60_io_b = cell_59_io_B; // @[mul.scala 114:25]
  assign cell_61_clock = clock;
  assign cell_61_reset = reset;
  assign cell_61_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_61_io_valid = cell_60_io_ready; // @[mul.scala 108:25]
  assign cell_61_io_a_in = cell_60_io_a_out; // @[mul.scala 109:25]
  assign cell_61_io_b_in = cell_60_io_b_out; // @[mul.scala 110:25]
  assign cell_61_io_sum_in = cell_60_io_sum_out; // @[mul.scala 111:25]
  assign cell_61_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_61_io_a = cell_60_io_A; // @[mul.scala 113:25]
  assign cell_61_io_b = cell_60_io_B; // @[mul.scala 114:25]
  assign cell_62_clock = clock;
  assign cell_62_reset = reset;
  assign cell_62_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_62_io_valid = cell_61_io_ready; // @[mul.scala 108:25]
  assign cell_62_io_a_in = cell_61_io_a_out; // @[mul.scala 109:25]
  assign cell_62_io_b_in = cell_61_io_b_out; // @[mul.scala 110:25]
  assign cell_62_io_sum_in = cell_61_io_sum_out; // @[mul.scala 111:25]
  assign cell_62_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_62_io_a = cell_61_io_A; // @[mul.scala 113:25]
  assign cell_62_io_b = cell_61_io_B; // @[mul.scala 114:25]
  assign cell_63_clock = clock;
  assign cell_63_reset = reset;
  assign cell_63_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_63_io_valid = cell_62_io_ready; // @[mul.scala 108:25]
  assign cell_63_io_a_in = cell_62_io_a_out; // @[mul.scala 109:25]
  assign cell_63_io_b_in = cell_62_io_b_out; // @[mul.scala 110:25]
  assign cell_63_io_sum_in = cell_62_io_sum_out; // @[mul.scala 111:25]
  assign cell_63_io_last = 1'h0; // @[mul.scala 112:25]
  assign cell_63_io_a = cell_62_io_A; // @[mul.scala 113:25]
  assign cell_63_io_b = cell_62_io_B; // @[mul.scala 114:25]
  assign cell_64_clock = clock;
  assign cell_64_reset = reset;
  assign cell_64_io_flush = 1'h0; // @[mul.scala 107:25]
  assign cell_64_io_valid = cell_63_io_ready; // @[mul.scala 108:25]
  assign cell_64_io_a_in = cell_63_io_a_out; // @[mul.scala 109:25]
  assign cell_64_io_b_in = cell_63_io_b_out; // @[mul.scala 110:25]
  assign cell_64_io_sum_in = cell_63_io_sum_out; // @[mul.scala 111:25]
  assign cell_64_io_last = 1'h1; // @[mul.scala 112:25]
  assign cell_64_io_a = cell_63_io_A; // @[mul.scala 113:25]
  assign cell_64_io_b = cell_63_io_B; // @[mul.scala 114:25]
  always @(posedge clock) begin
    a <= _GEN_1[128:0]; // @[mul.scala 77:{20,20} 81:7]
    b <= _GEN_2[128:0]; // @[mul.scala 78:{20,20} 87:7]
    if (reset) begin // @[mul.scala 79:24]
      valid <= 1'h0; // @[mul.scala 79:24]
    end else begin
      valid <= io_mul_valid; // @[mul.scala 93:10]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_out_valid & ~reset & ~(cell_64_io_sum_out == _GEN_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at mul.scala:124 chisel3.assert( cell(64).io.sum_out === (cell(64).io.A * cell(64).io.B))\n"
            ); // @[mul.scala 124:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_out_valid & ~reset & ~(cell_64_io_sum_out == _GEN_0)) begin
          $fatal; // @[mul.scala 124:23]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  a = _RAND_0[128:0];
  _RAND_1 = {5{`RANDOM}};
  b = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module div(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _dividend_abs_T_3 = ~io_dividend; // @[div.scala 20:27]
  wire [63:0] _dividend_abs_T_5 = _dividend_abs_T_3 + 64'h1; // @[div.scala 20:48]
  wire [63:0] dividend_abs = io_div_signed & io_dividend[63] ? _dividend_abs_T_5 : io_dividend; // @[div.scala 19:25]
  wire [63:0] _divisor_abs_T_3 = ~io_divisor; // @[div.scala 22:26]
  wire [63:0] _divisor_abs_T_5 = _divisor_abs_T_3 + 64'h1; // @[div.scala 22:46]
  wire [63:0] divisor_abs = io_div_signed & io_divisor[63] ? _divisor_abs_T_5 : io_divisor; // @[div.scala 21:24]
  reg [63:0] quotient; // @[div.scala 24:25]
  reg [63:0] remainder; // @[div.scala 25:26]
  reg [127:0] dividend; // @[div.scala 26:25]
  reg [64:0] divisor; // @[div.scala 27:24]
  reg [6:0] shift_count; // @[div.scala 29:28]
  reg  is_dividing; // @[div.scala 31:28]
  reg  is_dividing_signed; // @[div.scala 33:35]
  reg  quotient_sign; // @[div.scala 39:30]
  reg  remainder_sign; // @[div.scala 40:31]
  reg  out_valid; // @[div.scala 41:26]
  wire [64:0] sub = dividend[127:63] - divisor; // @[div.scala 43:36]
  wire  _io_div_ready_T = ~is_dividing; // @[div.scala 45:19]
  wire  _T_1 = io_div_valid & _io_div_ready_T; // @[div.scala 51:27]
  wire [127:0] _dividend_T = {64'h0,dividend_abs}; // @[Cat.scala 33:92]
  wire [64:0] _divisor_T = {1'h0,divisor_abs}; // @[Cat.scala 33:92]
  wire [63:0] _quotient_T = ~quotient; // @[div.scala 70:41]
  wire [63:0] _quotient_T_2 = _quotient_T + 64'h1; // @[div.scala 70:59]
  wire [63:0] _quotient_T_3 = quotient_sign ? _quotient_T_2 : quotient; // @[div.scala 70:24]
  wire [63:0] _remainder_T_1 = ~remainder; // @[div.scala 71:43]
  wire [63:0] _remainder_T_3 = _remainder_T_1 + 64'h1; // @[div.scala 71:62]
  wire [63:0] _remainder_T_4 = remainder_sign ? _remainder_T_3 : remainder; // @[div.scala 71:25]
  wire [63:0] _GEN_0 = is_dividing_signed ? _quotient_T_3 : quotient; // @[div.scala 69:32 70:18 24:25]
  wire [63:0] _GEN_1 = is_dividing_signed ? _remainder_T_4 : dividend[63:0]; // @[div.scala 67:17 69:32 71:19]
  wire [128:0] _dividend_T_1 = {dividend, 1'h0}; // @[div.scala 77:28]
  wire [64:0] _quotient_T_4 = {quotient, 1'h0}; // @[div.scala 78:28]
  wire [64:0] _quotient_T_6 = _quotient_T_4 | 65'h1; // @[div.scala 80:37]
  wire [127:0] _dividend_T_3 = {sub,dividend[62:0]}; // @[Cat.scala 33:92]
  wire [128:0] _dividend_T_4 = {_dividend_T_3, 1'h0}; // @[div.scala 81:47]
  wire [128:0] _GEN_2 = sub[64] ? _dividend_T_1 : _dividend_T_4; // @[div.scala 76:33 77:16 81:16]
  wire [64:0] _GEN_3 = sub[64] ? _quotient_T_4 : _quotient_T_6; // @[div.scala 76:33 78:16 80:16]
  wire  _GEN_4 = shift_count == 7'h0 ? 1'h0 : is_dividing; // @[div.scala 64:30 65:19 31:28]
  wire [64:0] _GEN_6 = shift_count == 7'h0 ? {{1'd0}, _GEN_0} : _GEN_3; // @[div.scala 64:30]
  wire  _GEN_7 = shift_count == 7'h0 | out_valid; // @[div.scala 64:30 74:17 41:26]
  wire [128:0] _GEN_8 = shift_count == 7'h0 ? {{1'd0}, dividend} : _GEN_2; // @[div.scala 26:25 64:30]
  wire [6:0] _shift_count_T_1 = shift_count - 7'h1; // @[div.scala 84:32]
  wire  _GEN_9 = is_dividing ? _GEN_4 : is_dividing; // @[div.scala 63:27 31:28]
  wire [64:0] _GEN_11 = is_dividing ? _GEN_6 : {{1'd0}, quotient}; // @[div.scala 24:25 63:27]
  wire  _GEN_12 = is_dividing & _GEN_7; // @[div.scala 63:27 88:15]
  wire [128:0] _GEN_13 = is_dividing ? _GEN_8 : {{1'd0}, dividend}; // @[div.scala 26:25 63:27]
  wire  _GEN_15 = io_div_valid & _io_div_ready_T | _GEN_9; // @[div.scala 51:44 52:17]
  wire [128:0] _GEN_18 = io_div_valid & _io_div_ready_T ? {{1'd0}, _dividend_T} : _GEN_13; // @[div.scala 51:44 55:14]
  wire [64:0] _GEN_20 = io_div_valid & _io_div_ready_T ? 65'h0 : _GEN_11; // @[div.scala 51:44 57:14]
  wire [64:0] _GEN_37 = reset ? 65'h0 : _GEN_20; // @[div.scala 24:{25,25}]
  wire [128:0] _GEN_38 = reset ? 129'h0 : _GEN_18; // @[div.scala 26:{25,25}]
  assign io_out_valid = out_valid; // @[div.scala 91:16]
  assign io_quotient = quotient; // @[div.scala 92:15]
  assign io_remainder = remainder; // @[div.scala 93:16]
  always @(posedge clock) begin
    quotient <= _GEN_37[63:0]; // @[div.scala 24:{25,25}]
    if (reset) begin // @[div.scala 25:26]
      remainder <= 64'h0; // @[div.scala 25:26]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      remainder <= 64'h0; // @[div.scala 58:15]
    end else if (is_dividing) begin // @[div.scala 63:27]
      if (shift_count == 7'h0) begin // @[div.scala 64:30]
        remainder <= _GEN_1;
      end
    end
    dividend <= _GEN_38[127:0]; // @[div.scala 26:{25,25}]
    if (reset) begin // @[div.scala 27:24]
      divisor <= 65'h0; // @[div.scala 27:24]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      divisor <= _divisor_T; // @[div.scala 56:13]
    end
    if (reset) begin // @[div.scala 29:28]
      shift_count <= 7'h40; // @[div.scala 29:28]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      shift_count <= 7'h40; // @[div.scala 59:17]
    end else if (is_dividing) begin // @[div.scala 63:27]
      shift_count <= _shift_count_T_1; // @[div.scala 84:17]
    end
    if (reset) begin // @[div.scala 31:28]
      is_dividing <= 1'h0; // @[div.scala 31:28]
    end else begin
      is_dividing <= _GEN_15;
    end
    if (reset) begin // @[div.scala 33:35]
      is_dividing_signed <= 1'h0; // @[div.scala 33:35]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      is_dividing_signed <= io_div_signed; // @[div.scala 54:24]
    end
    if (reset) begin // @[div.scala 39:30]
      quotient_sign <= 1'h0; // @[div.scala 39:30]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      quotient_sign <= io_dividend[63] ^ io_divisor[63]; // @[div.scala 60:19]
    end
    if (reset) begin // @[div.scala 40:31]
      remainder_sign <= 1'h0; // @[div.scala 40:31]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      remainder_sign <= io_dividend[63]; // @[div.scala 61:20]
    end
    if (reset) begin // @[div.scala 41:26]
      out_valid <= 1'h0; // @[div.scala 41:26]
    end else if (io_div_valid & _io_div_ready_T) begin // @[div.scala 51:44]
      out_valid <= 1'h0; // @[div.scala 62:15]
    end else begin
      out_valid <= _GEN_12;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_1 & is_dividing & ~reset) begin
          $fwrite(32'h80000002,"%d %x %x %x %x %x\n",shift_count,dividend,divisor,quotient,remainder,sub[64]); // @[div.scala 86:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  quotient = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  remainder = _RAND_1[63:0];
  _RAND_2 = {4{`RANDOM}};
  dividend = _RAND_2[127:0];
  _RAND_3 = {3{`RANDOM}};
  divisor = _RAND_3[64:0];
  _RAND_4 = {1{`RANDOM}};
  shift_count = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  is_dividing = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  is_dividing_signed = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quotient_sign = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  remainder_sign = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_valid = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [18:0] io_op,
  output [63:0] io_result,
  input         io_validin,
  output        io_validout
);
  wire  mul_pipe_clock; // @[ALU.scala 38:19]
  wire  mul_pipe_reset; // @[ALU.scala 38:19]
  wire  mul_pipe_io_mul_valid; // @[ALU.scala 38:19]
  wire [1:0] mul_pipe_io_mul_signed; // @[ALU.scala 38:19]
  wire [63:0] mul_pipe_io_multiplicand; // @[ALU.scala 38:19]
  wire [63:0] mul_pipe_io_multiplier; // @[ALU.scala 38:19]
  wire  mul_pipe_io_out_valid; // @[ALU.scala 38:19]
  wire [63:0] mul_pipe_io_result_lo; // @[ALU.scala 38:19]
  wire  div_clock; // @[ALU.scala 46:19]
  wire  div_reset; // @[ALU.scala 46:19]
  wire [63:0] div_io_dividend; // @[ALU.scala 46:19]
  wire [63:0] div_io_divisor; // @[ALU.scala 46:19]
  wire  div_io_div_valid; // @[ALU.scala 46:19]
  wire  div_io_div_signed; // @[ALU.scala 46:19]
  wire  div_io_out_valid; // @[ALU.scala 46:19]
  wire [63:0] div_io_quotient; // @[ALU.scala 46:19]
  wire [63:0] div_io_remainder; // @[ALU.scala 46:19]
  wire  _adder_b_T_6 = io_op[1] | io_op[8] | io_op[9] | io_op[11]; // @[ALU.scala 27:44]
  wire [63:0] _adder_b_T_7 = ~io_src2; // @[ALU.scala 27:55]
  wire [63:0] adder_b = io_op[1] | io_op[8] | io_op[9] | io_op[11] ? _adder_b_T_7 : io_src2; // @[ALU.scala 27:17]
  wire [64:0] _sum_T = io_src1 + adder_b; // @[ALU.scala 29:17]
  wire [64:0] _GEN_0 = {{64'd0}, _adder_b_T_6}; // @[ALU.scala 29:26]
  wire [65:0] _sum_T_1 = _sum_T + _GEN_0; // @[ALU.scala 29:26]
  wire [64:0] sum = _sum_T_1[64:0]; // @[ALU.scala 22:17 29:8]
  wire  adder_cout = sum[64]; // @[ALU.scala 30:20]
  wire [63:0] adder_result = sum[63:0]; // @[ALU.scala 31:22]
  wire  _slt_result_T_11 = io_src1[63] & ~io_src2[63] | ~(io_src1[63] ^ io_src2[63]) & adder_result[63]; // @[ALU.scala 33:61]
  wire [63:0] slt_result = {63'h0,_slt_result_T_11}; // @[Cat.scala 33:92]
  wire  _sltu_result_T_1 = ~adder_cout; // @[ALU.scala 34:35]
  wire [63:0] sltu_result = {63'h0,_sltu_result_T_1}; // @[Cat.scala 33:92]
  wire  _eql_result_T_1 = adder_result == 64'h0; // @[ALU.scala 35:46]
  wire [63:0] eql_result = {63'h0,_eql_result_T_1}; // @[Cat.scala 33:92]
  wire  _T_4 = io_op[12] | io_op[13] | io_op[14]; // @[ALU.scala 39:42]
  wire  _T_8 = io_op[13] | io_op[14]; // @[ALU.scala 41:35]
  wire  _T_13 = io_op[15] | io_op[16]; // @[ALU.scala 47:32]
  wire [63:0] _io_result_T_4 = io_src1 & io_src2; // @[ALU.scala 60:36]
  wire [63:0] _io_result_T_6 = io_src1 | io_src2; // @[ALU.scala 61:36]
  wire [63:0] _io_result_T_8 = io_src1 ^ io_src2; // @[ALU.scala 62:36]
  wire [126:0] _GEN_1 = {{63'd0}, io_src1}; // @[ALU.scala 63:37]
  wire [126:0] _io_result_T_11 = _GEN_1 << io_src2[5:0]; // @[ALU.scala 63:37]
  wire [63:0] _io_result_T_15 = io_src1 >> io_src2[5:0]; // @[ALU.scala 64:36]
  wire [63:0] _io_result_T_20 = $signed(io_src1) >>> io_src2[5:0]; // @[ALU.scala 65:62]
  wire [63:0] _io_result_T_25 = adder_result & 64'hfffffffffffffffe; // @[ALU.scala 68:42]
  wire [63:0] _io_result_T_38 = io_op[17] | io_op[18] ? div_io_remainder : 64'h0; // @[ALU.scala 72:19]
  wire [63:0] _io_result_T_39 = _T_13 ? div_io_quotient : _io_result_T_38; // @[ALU.scala 71:19]
  wire [63:0] _io_result_T_40 = _T_4 ? mul_pipe_io_result_lo : _io_result_T_39; // @[ALU.scala 70:19]
  wire [63:0] _io_result_T_41 = io_op[11] ? eql_result : _io_result_T_40; // @[ALU.scala 69:19]
  wire [63:0] _io_result_T_42 = io_op[10] ? _io_result_T_25 : _io_result_T_41; // @[ALU.scala 68:19]
  wire [63:0] _io_result_T_43 = io_op[9] ? sltu_result : _io_result_T_42; // @[ALU.scala 67:19]
  wire [63:0] _io_result_T_44 = io_op[8] ? slt_result : _io_result_T_43; // @[ALU.scala 66:19]
  wire [63:0] _io_result_T_45 = io_op[7] ? _io_result_T_20 : _io_result_T_44; // @[ALU.scala 65:19]
  wire [63:0] _io_result_T_46 = io_op[6] ? _io_result_T_15 : _io_result_T_45; // @[ALU.scala 64:19]
  wire [63:0] _io_result_T_47 = io_op[5] ? _io_result_T_11[63:0] : _io_result_T_46; // @[ALU.scala 63:19]
  wire [63:0] _io_result_T_48 = io_op[4] ? _io_result_T_8 : _io_result_T_47; // @[ALU.scala 62:19]
  wire [63:0] _io_result_T_49 = io_op[3] ? _io_result_T_6 : _io_result_T_48; // @[ALU.scala 61:19]
  wire [63:0] _io_result_T_50 = io_op[2] ? _io_result_T_4 : _io_result_T_49; // @[ALU.scala 60:19]
  mul_pipe mul_pipe ( // @[ALU.scala 38:19]
    .clock(mul_pipe_clock),
    .reset(mul_pipe_reset),
    .io_mul_valid(mul_pipe_io_mul_valid),
    .io_mul_signed(mul_pipe_io_mul_signed),
    .io_multiplicand(mul_pipe_io_multiplicand),
    .io_multiplier(mul_pipe_io_multiplier),
    .io_out_valid(mul_pipe_io_out_valid),
    .io_result_lo(mul_pipe_io_result_lo)
  );
  div div ( // @[ALU.scala 46:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_dividend(div_io_dividend),
    .io_divisor(div_io_divisor),
    .io_div_valid(div_io_div_valid),
    .io_div_signed(div_io_div_signed),
    .io_out_valid(div_io_out_valid),
    .io_quotient(div_io_quotient),
    .io_remainder(div_io_remainder)
  );
  assign io_result = io_op[0] | io_op[1] ? adder_result : _io_result_T_50; // @[ALU.scala 59:19]
  assign io_validout = ~(_T_4 | io_op[15] | io_op[16] | io_op[17] | io_op[18]) | mul_pipe_io_out_valid |
    div_io_out_valid; // @[ALU.scala 57:108]
  assign mul_pipe_clock = clock;
  assign mul_pipe_reset = reset;
  assign mul_pipe_io_mul_valid = (io_op[12] | io_op[13] | io_op[14]) & io_validin; // @[ALU.scala 39:53]
  assign mul_pipe_io_mul_signed = {_T_8,io_op[13]}; // @[Cat.scala 33:92]
  assign mul_pipe_io_multiplicand = io_src1; // @[ALU.scala 42:21]
  assign mul_pipe_io_multiplier = io_src2; // @[ALU.scala 43:19]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_dividend = io_src1; // @[ALU.scala 50:17]
  assign div_io_divisor = io_src2; // @[ALU.scala 51:16]
  assign div_io_div_valid = (io_op[15] | io_op[16] | io_op[17] | io_op[18]) & io_validin; // @[ALU.scala 47:63]
  assign div_io_div_signed = io_op[15] | io_op[17]; // @[ALU.scala 49:30]
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [31:0] io_in_bits_inst,
  input  [4:0]  io_in_bits_rs1,
  input  [4:0]  io_in_bits_rs2,
  input  [4:0]  io_in_bits_rd,
  input  [63:0] io_in_bits_imm,
  input  [79:0] io_in_bits_op,
  input  [5:0]  io_in_bits_typ,
  input         io_in_bits_isJump,
  input  [4:0]  io_in_bits_clearidx,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_pc,
  output [63:0] io_out_bits_pc_dnpc,
  output [4:0]  io_out_bits_gpr_idx_w,
  output        io_out_bits_gpr_en_w,
  output [63:0] io_out_bits_gpr_val_w,
  output        io_out_bits_csr_en_w,
  output [11:0] io_out_bits_csr_idx_w,
  output [63:0] io_out_bits_csr_val_w,
  output [63:0] io_out_bits_csr_no,
  output [63:0] io_out_bits_csr_epc,
  output        io_out_bits_isJump,
  output [4:0]  io_out_bits_clearidx,
  output [4:0]  io_gpr_idx_r1,
  output [4:0]  io_gpr_idx_r2,
  output        io_gpr_en_r1,
  output        io_gpr_en_r2,
  input  [63:0] io_gpr_val_r1,
  input  [63:0] io_gpr_val_r2,
  output [11:0] io_csr_idx_r,
  output        io_csr_en_r,
  input  [63:0] io_csr_val_r,
  input         io_lm_ar_ready,
  output        io_lm_ar_valid,
  output [31:0] io_lm_ar_bits_addr,
  output        io_lm_r_ready,
  input         io_lm_r_valid,
  input  [63:0] io_lm_r_bits_data,
  input         io_lm_aw_ready,
  output        io_lm_aw_valid,
  output [31:0] io_lm_aw_bits_addr,
  input         io_lm_w_ready,
  output        io_lm_w_valid,
  output [63:0] io_lm_w_bits_data,
  output [7:0]  io_lm_w_bits_strb,
  input         io_lm_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  lsu_clock; // @[EXU.scala 39:25]
  wire  lsu_reset; // @[EXU.scala 39:25]
  wire  lsu_io_ls_in_valid; // @[EXU.scala 39:25]
  wire [31:0] lsu_io_ls_in_bits_raddr; // @[EXU.scala 39:25]
  wire [31:0] lsu_io_ls_in_bits_waddr; // @[EXU.scala 39:25]
  wire [63:0] lsu_io_ls_in_bits_wdata; // @[EXU.scala 39:25]
  wire [7:0] lsu_io_ls_in_bits_wmask; // @[EXU.scala 39:25]
  wire  lsu_io_ls_out_ready; // @[EXU.scala 39:25]
  wire  lsu_io_ls_out_valid; // @[EXU.scala 39:25]
  wire [63:0] lsu_io_ls_out_bits_rdata; // @[EXU.scala 39:25]
  wire  lsu_io_en_r; // @[EXU.scala 39:25]
  wire  lsu_io_en_w; // @[EXU.scala 39:25]
  wire  lsu_io_lm_ar_ready; // @[EXU.scala 39:25]
  wire  lsu_io_lm_ar_valid; // @[EXU.scala 39:25]
  wire [31:0] lsu_io_lm_ar_bits_addr; // @[EXU.scala 39:25]
  wire  lsu_io_lm_r_ready; // @[EXU.scala 39:25]
  wire  lsu_io_lm_r_valid; // @[EXU.scala 39:25]
  wire [63:0] lsu_io_lm_r_bits_data; // @[EXU.scala 39:25]
  wire  lsu_io_lm_aw_ready; // @[EXU.scala 39:25]
  wire  lsu_io_lm_aw_valid; // @[EXU.scala 39:25]
  wire [31:0] lsu_io_lm_aw_bits_addr; // @[EXU.scala 39:25]
  wire  lsu_io_lm_w_ready; // @[EXU.scala 39:25]
  wire  lsu_io_lm_w_valid; // @[EXU.scala 39:25]
  wire [63:0] lsu_io_lm_w_bits_data; // @[EXU.scala 39:25]
  wire [7:0] lsu_io_lm_w_bits_strb; // @[EXU.scala 39:25]
  wire  lsu_io_lm_b_ready; // @[EXU.scala 39:25]
  wire  lsu_io_lm_b_valid; // @[EXU.scala 39:25]
  wire  alu_clock; // @[EXU.scala 64:23]
  wire  alu_reset; // @[EXU.scala 64:23]
  wire [63:0] alu_io_src1; // @[EXU.scala 64:23]
  wire [63:0] alu_io_src2; // @[EXU.scala 64:23]
  wire [18:0] alu_io_op; // @[EXU.scala 64:23]
  wire [63:0] alu_io_result; // @[EXU.scala 64:23]
  wire  alu_io_validin; // @[EXU.scala 64:23]
  wire  alu_io_validout; // @[EXU.scala 64:23]
  wire  ebreak1_en_break; // @[EXU.scala 108:27]
  wire  ebreak1_clk; // @[EXU.scala 108:27]
  wire  _EXE_reg_pc_T = io_in_ready & io_in_valid; // @[Decoupled.scala 52:35]
  reg [31:0] EXE_reg_pc; // @[Reg.scala 35:20]
  reg [31:0] EXE_reg_inst; // @[Reg.scala 35:20]
  reg [4:0] EXE_reg_rs1; // @[Reg.scala 35:20]
  reg [4:0] EXE_reg_rs2; // @[Reg.scala 35:20]
  reg [4:0] EXE_reg_rd; // @[Reg.scala 35:20]
  reg [63:0] EXE_reg_imm; // @[Reg.scala 35:20]
  reg [79:0] EXE_reg_op; // @[Reg.scala 35:20]
  reg [5:0] EXE_reg_typ; // @[Reg.scala 35:20]
  reg  EXE_reg_isJump; // @[Reg.scala 35:20]
  reg [4:0] EXE_reg_clearidx; // @[Reg.scala 35:20]
  wire  op_r = EXE_reg_op[38] | EXE_reg_op[39] | EXE_reg_op[40] | EXE_reg_op[41] | EXE_reg_op[46] | EXE_reg_op[47] |
    EXE_reg_op[48]; // @[EXU.scala 45:110]
  wire  op_w = EXE_reg_op[42] | EXE_reg_op[43] | EXE_reg_op[44] | EXE_reg_op[45]; // @[EXU.scala 46:62]
  wire  _op_mul_T_2 = EXE_reg_op[50] | EXE_reg_op[51]; // @[EXU.scala 47:31]
  wire  op_mul = EXE_reg_op[50] | EXE_reg_op[51] | EXE_reg_op[52] | EXE_reg_op[53] | EXE_reg_op[54]; // @[EXU.scala 47:76]
  wire  _op_div_T_2 = EXE_reg_op[55] | EXE_reg_op[56]; // @[EXU.scala 48:31]
  wire  op_div = EXE_reg_op[55] | EXE_reg_op[56] | EXE_reg_op[57] | EXE_reg_op[58]; // @[EXU.scala 48:61]
  wire  _src1_T_4 = EXE_reg_typ[0] | EXE_reg_typ[2] | EXE_reg_typ[4]; // @[EXU.scala 53:49]
  wire [63:0] _src1_T_10 = EXE_reg_typ[1] | EXE_reg_typ[3] ? EXE_reg_imm : 64'h0; // @[EXU.scala 54:16]
  wire [63:0] src1 = EXE_reg_typ[0] | EXE_reg_typ[2] | EXE_reg_typ[4] | EXE_reg_typ[5] ? io_gpr_val_r1 : _src1_T_10; // @[EXU.scala 53:18]
  wire  _src2_T_2 = EXE_reg_typ[2] | EXE_reg_typ[4]; // @[EXU.scala 57:34]
  wire [63:0] _src2_T_6 = EXE_reg_typ[0] ? EXE_reg_imm : 64'h0; // @[EXU.scala 58:16]
  wire [63:0] src2 = EXE_reg_typ[2] | EXE_reg_typ[4] | EXE_reg_typ[5] ? io_gpr_val_r2 : _src2_T_6; // @[EXU.scala 57:18]
  wire [63:0] dest = _src2_T_2 ? EXE_reg_imm : {{59'd0}, EXE_reg_rd}; // @[EXU.scala 61:18]
  reg  lsu_finish; // @[EXU.scala 66:31]
  reg  alu_finish; // @[EXU.scala 67:31]
  reg [1:0] state; // @[EXU.scala 71:28]
  wire  _lsu_finish_T = state != 2'h1; // @[EXU.scala 73:33]
  wire  _lsu_finish_T_1 = lsu_io_ls_out_ready & lsu_io_ls_out_valid; // @[Decoupled.scala 52:35]
  wire  _lsu_finish_T_7 = _lsu_finish_T_1 | ~op_r & ~op_w | lsu_finish; // @[EXU.scala 74:26]
  wire  _alu_finish_T_6 = alu_io_validout | ~op_mul & ~op_div | alu_finish; // @[EXU.scala 76:26]
  wire [1:0] _state_T_1 = _EXE_reg_pc_T ? 2'h1 : 2'h0; // @[EXU.scala 80:26]
  wire  _state_T_6 = io_out_ready & io_out_valid; // @[Decoupled.scala 52:35]
  wire  _lsu_io_ls_in_valid_T = state == 2'h1; // @[EXU.scala 95:36]
  wire [63:0] _lsu_io_ls_in_bits_raddr_T_13 = op_r ? alu_io_result : 64'h0; // @[EXU.scala 96:37]
  wire [63:0] _lsu_io_ls_in_bits_waddr_T_7 = op_w ? alu_io_result : 64'h0; // @[EXU.scala 97:37]
  wire [7:0] _lsu_io_ls_in_bits_wmask_T_13 = EXE_reg_op[45] ? 8'hff : 8'h0; // @[EXU.scala 102:35]
  wire [7:0] _lsu_io_ls_in_bits_wmask_T_14 = EXE_reg_op[44] ? 8'hf : _lsu_io_ls_in_bits_wmask_T_13; // @[EXU.scala 101:35]
  wire [7:0] _lsu_io_ls_in_bits_wmask_T_15 = EXE_reg_op[43] ? 8'h3 : _lsu_io_ls_in_bits_wmask_T_14; // @[EXU.scala 100:35]
  wire  _io_csr_en_r_T_2 = EXE_reg_op[63] | EXE_reg_op[64]; // @[EXU.scala 120:40]
  wire [63:0] _io_csr_idx_r_T_3 = _io_csr_en_r_T_2 ? src2 : 64'h0; // @[EXU.scala 121:26]
  reg  alu_wait; // @[EXU.scala 129:29]
  wire [63:0] _alu_io_src1_T_15 = {32'h0,src1[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _alu_io_src1_T_21 = src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _alu_io_src1_T_23 = {_alu_io_src1_T_21,src1[31:0]}; // @[Cat.scala 33:92]
  wire  _alu_io_src1_T_26 = EXE_reg_op[36] | EXE_reg_op[37]; // @[EXU.scala 135:43]
  wire [63:0] _alu_io_src1_T_27 = EXE_reg_op[36] | EXE_reg_op[37] ? {{32'd0}, EXE_reg_pc} : src1; // @[EXU.scala 135:28]
  wire [63:0] _alu_io_src1_T_28 = EXE_reg_op[17] | EXE_reg_op[19] ? _alu_io_src1_T_23 : _alu_io_src1_T_27; // @[EXU.scala 134:28]
  wire [63:0] _alu_io_src2_T_7 = {59'h0,src2[4:0]}; // @[Cat.scala 33:92]
  wire [63:0] _alu_io_src2_T_28 = {32'h0,src2[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _alu_io_src2_T_30 = EXE_reg_op[64] ? io_csr_val_r : src2; // @[EXU.scala 142:28]
  wire [63:0] _alu_io_src2_T_31 = EXE_reg_op[56] | EXE_reg_op[58] | EXE_reg_op[60] | EXE_reg_op[62] ? _alu_io_src2_T_28
     : _alu_io_src2_T_30; // @[EXU.scala 141:28]
  wire [63:0] _alu_io_src2_T_32 = op_w ? dest : _alu_io_src2_T_31; // @[EXU.scala 140:28]
  wire [63:0] _alu_io_src2_T_33 = _alu_io_src1_T_26 ? 64'h4 : _alu_io_src2_T_32; // @[EXU.scala 139:28]
  wire [63:0] _alu_io_src2_T_34 = EXE_reg_op[25] ? {{32'd0}, EXE_reg_pc} : _alu_io_src2_T_33; // @[EXU.scala 138:28]
  wire [18:0] _alu_io_op_T_108 = EXE_reg_op[61] | EXE_reg_op[62] ? 19'h40000 : 19'h0; // @[EXU.scala 161:28]
  wire [18:0] _alu_io_op_T_109 = EXE_reg_op[59] | EXE_reg_op[60] ? 19'h20000 : _alu_io_op_T_108; // @[EXU.scala 160:28]
  wire [18:0] _alu_io_op_T_110 = EXE_reg_op[57] | EXE_reg_op[58] ? 19'h10000 : _alu_io_op_T_109; // @[EXU.scala 159:28]
  wire [18:0] _alu_io_op_T_111 = _op_div_T_2 ? 19'h8000 : _alu_io_op_T_110; // @[EXU.scala 158:28]
  wire [18:0] _alu_io_op_T_112 = EXE_reg_op[54] ? 19'h4000 : _alu_io_op_T_111; // @[EXU.scala 157:28]
  wire [18:0] _alu_io_op_T_113 = EXE_reg_op[52] ? 19'h2000 : _alu_io_op_T_112; // @[EXU.scala 156:28]
  wire [18:0] _alu_io_op_T_114 = _op_mul_T_2 | EXE_reg_op[53] ? 19'h1000 : _alu_io_op_T_113; // @[EXU.scala 155:28]
  wire [18:0] _alu_io_op_T_115 = EXE_reg_op[30] | EXE_reg_op[31] ? 19'h800 : _alu_io_op_T_114; // @[EXU.scala 154:28]
  wire [18:0] _alu_io_op_T_116 = EXE_reg_op[27] | EXE_reg_op[29] | EXE_reg_op[33] | EXE_reg_op[35] ? 19'h200 :
    _alu_io_op_T_115; // @[EXU.scala 153:28]
  wire [18:0] _alu_io_op_T_117 = EXE_reg_op[26] | EXE_reg_op[28] | EXE_reg_op[32] | EXE_reg_op[34] ? 19'h100 :
    _alu_io_op_T_116; // @[EXU.scala 152:28]
  wire [18:0] _alu_io_op_T_118 = EXE_reg_op[16] | EXE_reg_op[17] | EXE_reg_op[18] | EXE_reg_op[19] ? 19'h80 :
    _alu_io_op_T_117; // @[EXU.scala 151:28]
  wire [18:0] _alu_io_op_T_119 = EXE_reg_op[20] | EXE_reg_op[21] | EXE_reg_op[22] | EXE_reg_op[23] ? 19'h40 :
    _alu_io_op_T_118; // @[EXU.scala 150:28]
  wire [18:0] _alu_io_op_T_120 = EXE_reg_op[12] | EXE_reg_op[13] | EXE_reg_op[14] | EXE_reg_op[15] ? 19'h20 :
    _alu_io_op_T_119; // @[EXU.scala 149:28]
  wire [18:0] _alu_io_op_T_121 = EXE_reg_op[10] | EXE_reg_op[11] ? 19'h10 : _alu_io_op_T_120; // @[EXU.scala 148:28]
  wire [18:0] _alu_io_op_T_122 = EXE_reg_op[8] | EXE_reg_op[9] | EXE_reg_op[64] ? 19'h8 : _alu_io_op_T_121; // @[EXU.scala 147:28]
  wire [18:0] _alu_io_op_T_123 = EXE_reg_op[6] | EXE_reg_op[7] ? 19'h4 : _alu_io_op_T_122; // @[EXU.scala 146:28]
  wire [18:0] _alu_io_op_T_124 = EXE_reg_op[4] | EXE_reg_op[5] ? 19'h2 : _alu_io_op_T_123; // @[EXU.scala 145:28]
  wire [63:0] next_pc_src1 = EXE_reg_op[37] ? src1 : {{32'd0}, EXE_reg_pc}; // @[EXU.scala 168:26]
  wire  _next_pc_src2_T_5 = ~alu_io_result[0]; // @[EXU.scala 170:43]
  wire [63:0] _next_pc_src2_T_23 = EXE_reg_op[37] ? src2 : 64'h4; // @[EXU.scala 176:26]
  wire [63:0] _next_pc_src2_T_24 = EXE_reg_op[36] ? src1 : _next_pc_src2_T_23; // @[EXU.scala 175:26]
  wire [63:0] _next_pc_src2_T_25 = EXE_reg_op[35] & alu_io_result[0] ? dest : _next_pc_src2_T_24; // @[EXU.scala 174:26]
  wire [63:0] _next_pc_src2_T_26 = EXE_reg_op[34] & alu_io_result[0] ? dest : _next_pc_src2_T_25; // @[EXU.scala 173:26]
  wire [63:0] _next_pc_src2_T_27 = EXE_reg_op[33] & _next_pc_src2_T_5 ? dest : _next_pc_src2_T_26; // @[EXU.scala 172:26]
  wire [63:0] _next_pc_src2_T_28 = EXE_reg_op[32] & _next_pc_src2_T_5 ? dest : _next_pc_src2_T_27; // @[EXU.scala 171:26]
  wire [63:0] _next_pc_src2_T_29 = EXE_reg_op[31] & ~alu_io_result[0] ? dest : _next_pc_src2_T_28; // @[EXU.scala 170:26]
  wire [63:0] next_pc_src2 = EXE_reg_op[30] & alu_io_result[0] ? dest : _next_pc_src2_T_29; // @[EXU.scala 169:26]
  wire [63:0] next_pc_sum = next_pc_src1 + next_pc_src2; // @[EXU.scala 178:34]
  wire [1:0] _io_out_bits_csr_no_T_2 = EXE_reg_op[66] ? 2'h2 : 2'h0; // @[EXU.scala 187:32]
  wire [1:0] _io_out_bits_csr_no_T_3 = EXE_reg_op[65] ? 2'h1 : _io_out_bits_csr_no_T_2; // @[EXU.scala 186:32]
  wire [31:0] _io_out_bits_gpr_val_w_T_25 = alu_io_result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_gpr_val_w_T_27 = {_io_out_bits_gpr_val_w_T_25,alu_io_result[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_gpr_val_w_T_35 = {32'h0,alu_io_result[63:32]}; // @[Cat.scala 33:92]
  wire [55:0] _io_out_bits_gpr_val_w_T_42 = lsu_io_ls_out_bits_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_gpr_val_w_T_44 = {_io_out_bits_gpr_val_w_T_42,lsu_io_ls_out_bits_rdata[7:0]}; // @[Cat.scala 33:92]
  wire [47:0] _io_out_bits_gpr_val_w_T_48 = lsu_io_ls_out_bits_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_gpr_val_w_T_50 = {_io_out_bits_gpr_val_w_T_48,lsu_io_ls_out_bits_rdata[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _io_out_bits_gpr_val_w_T_54 = lsu_io_ls_out_bits_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_bits_gpr_val_w_T_56 = {_io_out_bits_gpr_val_w_T_54,lsu_io_ls_out_bits_rdata[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_gpr_val_w_T_61 = {56'h0,lsu_io_ls_out_bits_rdata[7:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_gpr_val_w_T_65 = {48'h0,lsu_io_ls_out_bits_rdata[15:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_gpr_val_w_T_69 = {32'h0,lsu_io_ls_out_bits_rdata[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _io_out_bits_gpr_val_w_T_70 = EXE_reg_op[48] ? _io_out_bits_gpr_val_w_T_69 : alu_io_result; // @[EXU.scala 199:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_71 = EXE_reg_op[47] ? _io_out_bits_gpr_val_w_T_65 : _io_out_bits_gpr_val_w_T_70; // @[EXU.scala 198:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_72 = EXE_reg_op[46] ? _io_out_bits_gpr_val_w_T_61 : _io_out_bits_gpr_val_w_T_71; // @[EXU.scala 197:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_73 = EXE_reg_op[41] ? lsu_io_ls_out_bits_rdata : _io_out_bits_gpr_val_w_T_72; // @[EXU.scala 196:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_74 = EXE_reg_op[40] ? _io_out_bits_gpr_val_w_T_56 : _io_out_bits_gpr_val_w_T_73; // @[EXU.scala 195:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_75 = EXE_reg_op[39] ? _io_out_bits_gpr_val_w_T_50 : _io_out_bits_gpr_val_w_T_74; // @[EXU.scala 194:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_76 = EXE_reg_op[38] ? _io_out_bits_gpr_val_w_T_44 : _io_out_bits_gpr_val_w_T_75; // @[EXU.scala 193:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_77 = _io_csr_en_r_T_2 ? io_csr_val_r : _io_out_bits_gpr_val_w_T_76; // @[EXU.scala 192:26]
  wire [63:0] _io_out_bits_gpr_val_w_T_78 = EXE_reg_op[52] | EXE_reg_op[53] | EXE_reg_op[54] ?
    _io_out_bits_gpr_val_w_T_35 : _io_out_bits_gpr_val_w_T_77; // @[EXU.scala 191:26]
  wire [63:0] _io_out_bits_csr_val_w_T_2 = EXE_reg_op[64] ? alu_io_result : 64'h0; // @[EXU.scala 203:26]
  wire [63:0] _io_out_bits_pc_dnpc_T_5 = next_pc_sum & 64'hfffffffffffffffe; // @[EXU.scala 206:60]
  wire [63:0] _io_out_bits_pc_dnpc_T_6 = EXE_reg_op[37] ? _io_out_bits_pc_dnpc_T_5 : next_pc_sum; // @[EXU.scala 206:33]
  LSU lsu ( // @[EXU.scala 39:25]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_ls_in_valid(lsu_io_ls_in_valid),
    .io_ls_in_bits_raddr(lsu_io_ls_in_bits_raddr),
    .io_ls_in_bits_waddr(lsu_io_ls_in_bits_waddr),
    .io_ls_in_bits_wdata(lsu_io_ls_in_bits_wdata),
    .io_ls_in_bits_wmask(lsu_io_ls_in_bits_wmask),
    .io_ls_out_ready(lsu_io_ls_out_ready),
    .io_ls_out_valid(lsu_io_ls_out_valid),
    .io_ls_out_bits_rdata(lsu_io_ls_out_bits_rdata),
    .io_en_r(lsu_io_en_r),
    .io_en_w(lsu_io_en_w),
    .io_lm_ar_ready(lsu_io_lm_ar_ready),
    .io_lm_ar_valid(lsu_io_lm_ar_valid),
    .io_lm_ar_bits_addr(lsu_io_lm_ar_bits_addr),
    .io_lm_r_ready(lsu_io_lm_r_ready),
    .io_lm_r_valid(lsu_io_lm_r_valid),
    .io_lm_r_bits_data(lsu_io_lm_r_bits_data),
    .io_lm_aw_ready(lsu_io_lm_aw_ready),
    .io_lm_aw_valid(lsu_io_lm_aw_valid),
    .io_lm_aw_bits_addr(lsu_io_lm_aw_bits_addr),
    .io_lm_w_ready(lsu_io_lm_w_ready),
    .io_lm_w_valid(lsu_io_lm_w_valid),
    .io_lm_w_bits_data(lsu_io_lm_w_bits_data),
    .io_lm_w_bits_strb(lsu_io_lm_w_bits_strb),
    .io_lm_b_ready(lsu_io_lm_b_ready),
    .io_lm_b_valid(lsu_io_lm_b_valid)
  );
  ALU alu ( // @[EXU.scala 64:23]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_src1(alu_io_src1),
    .io_src2(alu_io_src2),
    .io_op(alu_io_op),
    .io_result(alu_io_result),
    .io_validin(alu_io_validin),
    .io_validout(alu_io_validout)
  );
  ebreak ebreak1 ( // @[EXU.scala 108:27]
    .en_break(ebreak1_en_break),
    .clk(ebreak1_clk)
  );
  assign io_in_ready = state == 2'h0; // @[EXU.scala 88:29]
  assign io_out_valid = state == 2'h2; // @[EXU.scala 89:30]
  assign io_out_bits_pc = EXE_reg_pc; // @[EXU.scala 209:23]
  assign io_out_bits_pc_dnpc = EXE_reg_op[65] | EXE_reg_op[66] ? io_csr_val_r : _io_out_bits_pc_dnpc_T_6; // @[EXU.scala 205:33]
  assign io_out_bits_gpr_idx_w = dest[4:0]; // @[EXU.scala 182:30]
  assign io_out_bits_gpr_en_w = EXE_reg_typ[0] | EXE_reg_typ[1] | EXE_reg_typ[3] | EXE_reg_typ[5]; // @[EXU.scala 181:80]
  assign io_out_bits_gpr_val_w = EXE_reg_op[1] | EXE_reg_op[3] | EXE_reg_op[5] | EXE_reg_op[13] | EXE_reg_op[15] |
    EXE_reg_op[17] | EXE_reg_op[21] | EXE_reg_op[23] | EXE_reg_op[51] | EXE_reg_op[56] | EXE_reg_op[60] | EXE_reg_op[62]
     ? _io_out_bits_gpr_val_w_T_27 : _io_out_bits_gpr_val_w_T_78; // @[EXU.scala 190:35]
  assign io_out_bits_csr_en_w = EXE_reg_op[63] | EXE_reg_op[64]; // @[EXU.scala 184:50]
  assign io_out_bits_csr_idx_w = _io_csr_idx_r_T_3[11:0]; // @[EXU.scala 185:30]
  assign io_out_bits_csr_val_w = EXE_reg_op[63] ? src1 : _io_out_bits_csr_val_w_T_2; // @[EXU.scala 202:35]
  assign io_out_bits_csr_no = {{62'd0}, _io_out_bits_csr_no_T_3}; // @[EXU.scala 186:27]
  assign io_out_bits_csr_epc = {{32'd0}, EXE_reg_pc}; // @[EXU.scala 189:28]
  assign io_out_bits_isJump = EXE_reg_isJump; // @[EXU.scala 35:27]
  assign io_out_bits_clearidx = EXE_reg_clearidx; // @[EXU.scala 37:29]
  assign io_gpr_idx_r1 = EXE_reg_rs1; // @[EXU.scala 116:22]
  assign io_gpr_idx_r2 = EXE_reg_rs2; // @[EXU.scala 117:22]
  assign io_gpr_en_r1 = _src1_T_4 | EXE_reg_typ[5]; // @[EXU.scala 114:72]
  assign io_gpr_en_r2 = _src2_T_2 | EXE_reg_typ[5]; // @[EXU.scala 115:57]
  assign io_csr_idx_r = _io_csr_idx_r_T_3[11:0]; // @[EXU.scala 121:21]
  assign io_csr_en_r = EXE_reg_op[63] | EXE_reg_op[64]; // @[EXU.scala 120:40]
  assign io_lm_ar_valid = lsu_io_lm_ar_valid; // @[EXU.scala 105:14]
  assign io_lm_ar_bits_addr = lsu_io_lm_ar_bits_addr; // @[EXU.scala 105:14]
  assign io_lm_r_ready = lsu_io_lm_r_ready; // @[EXU.scala 105:14]
  assign io_lm_aw_valid = lsu_io_lm_aw_valid; // @[EXU.scala 105:14]
  assign io_lm_aw_bits_addr = lsu_io_lm_aw_bits_addr; // @[EXU.scala 105:14]
  assign io_lm_w_valid = lsu_io_lm_w_valid; // @[EXU.scala 105:14]
  assign io_lm_w_bits_data = lsu_io_lm_w_bits_data; // @[EXU.scala 105:14]
  assign io_lm_w_bits_strb = lsu_io_lm_w_bits_strb; // @[EXU.scala 105:14]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_ls_in_valid = state == 2'h1 & (op_w | op_r) & ~lsu_finish; // @[EXU.scala 95:62]
  assign lsu_io_ls_in_bits_raddr = _lsu_io_ls_in_bits_raddr_T_13[31:0]; // @[EXU.scala 96:32]
  assign lsu_io_ls_in_bits_waddr = _lsu_io_ls_in_bits_waddr_T_7[31:0]; // @[EXU.scala 97:32]
  assign lsu_io_ls_in_bits_wdata = op_w ? io_gpr_val_r2 : 64'h0; // @[EXU.scala 98:37]
  assign lsu_io_ls_in_bits_wmask = EXE_reg_op[42] ? 8'h1 : _lsu_io_ls_in_bits_wmask_T_15; // @[EXU.scala 99:37]
  assign lsu_io_ls_out_ready = 1'h1; // @[EXU.scala 94:28]
  assign lsu_io_en_r = EXE_reg_op[38] | EXE_reg_op[39] | EXE_reg_op[40] | EXE_reg_op[41] | EXE_reg_op[46] | EXE_reg_op[
    47] | EXE_reg_op[48]; // @[EXU.scala 45:110]
  assign lsu_io_en_w = EXE_reg_op[42] | EXE_reg_op[43] | EXE_reg_op[44] | EXE_reg_op[45]; // @[EXU.scala 46:62]
  assign lsu_io_lm_ar_ready = io_lm_ar_ready; // @[EXU.scala 105:14]
  assign lsu_io_lm_r_valid = io_lm_r_valid; // @[EXU.scala 105:14]
  assign lsu_io_lm_r_bits_data = io_lm_r_bits_data; // @[EXU.scala 105:14]
  assign lsu_io_lm_aw_ready = io_lm_aw_ready; // @[EXU.scala 105:14]
  assign lsu_io_lm_w_ready = io_lm_w_ready; // @[EXU.scala 105:14]
  assign lsu_io_lm_b_valid = io_lm_b_valid; // @[EXU.scala 105:14]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_src1 = EXE_reg_op[13] | EXE_reg_op[21] | EXE_reg_op[23] | EXE_reg_op[56] | EXE_reg_op[58] | EXE_reg_op[
    60] | EXE_reg_op[62] ? _alu_io_src1_T_15 : _alu_io_src1_T_28; // @[EXU.scala 133:28]
  assign alu_io_src2 = EXE_reg_op[13] | EXE_reg_op[17] | EXE_reg_op[21] ? _alu_io_src2_T_7 : _alu_io_src2_T_34; // @[EXU.scala 137:28]
  assign alu_io_op = EXE_reg_op[0] | EXE_reg_op[1] | EXE_reg_op[2] | EXE_reg_op[3] | EXE_reg_op[24] | EXE_reg_op[25] |
    EXE_reg_op[36] | EXE_reg_op[37] | EXE_reg_op[38] | EXE_reg_op[39] | EXE_reg_op[40] | EXE_reg_op[41] | EXE_reg_op[42]
     | EXE_reg_op[43] | EXE_reg_op[44] | EXE_reg_op[45] | EXE_reg_op[46] | EXE_reg_op[47] | EXE_reg_op[48] ? 19'h1 :
    _alu_io_op_T_124; // @[EXU.scala 144:28]
  assign alu_io_validin = _lsu_io_ls_in_valid_T & (op_mul | op_div) & ~alu_finish & ~alu_wait; // @[EXU.scala 131:79]
  assign ebreak1_en_break = EXE_reg_op[49] & _EXE_reg_pc_T; // @[EXU.scala 109:44]
  assign ebreak1_clk = clock; // @[EXU.scala 110:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_pc <= 32'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_pc <= io_in_bits_pc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_inst <= 32'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_inst <= io_in_bits_inst; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_rs1 <= 5'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_rs1 <= io_in_bits_rs1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_rs2 <= 5'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_rs2 <= io_in_bits_rs2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_rd <= 5'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_rd <= io_in_bits_rd; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_imm <= 64'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_imm <= io_in_bits_imm; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_op <= 80'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_op <= io_in_bits_op; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_typ <= 6'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_typ <= io_in_bits_typ; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_isJump <= 1'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_isJump <= io_in_bits_isJump; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      EXE_reg_clearidx <= 5'h0; // @[Reg.scala 35:20]
    end else if (_EXE_reg_pc_T) begin // @[Reg.scala 36:18]
      EXE_reg_clearidx <= io_in_bits_clearidx; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[EXU.scala 66:31]
      lsu_finish <= 1'h0; // @[EXU.scala 66:31]
    end else if (state != 2'h1) begin // @[EXU.scala 73:26]
      lsu_finish <= 1'h0;
    end else begin
      lsu_finish <= _lsu_finish_T_7;
    end
    if (reset) begin // @[EXU.scala 67:31]
      alu_finish <= 1'h0; // @[EXU.scala 67:31]
    end else if (_lsu_finish_T) begin // @[EXU.scala 75:26]
      alu_finish <= 1'h0;
    end else begin
      alu_finish <= _alu_finish_T_6;
    end
    if (reset) begin // @[EXU.scala 71:28]
      state <= 2'h0; // @[EXU.scala 71:28]
    end else if (2'h2 == state) begin // @[Mux.scala 81:58]
      if (_state_T_6) begin // @[EXU.scala 82:31]
        state <= 2'h0;
      end else begin
        state <= 2'h2;
      end
    end else if (2'h1 == state) begin // @[Mux.scala 81:58]
      if (lsu_finish & alu_finish) begin // @[EXU.scala 81:26]
        state <= 2'h2;
      end else begin
        state <= 2'h1;
      end
    end else if (2'h0 == state) begin // @[Mux.scala 81:58]
      state <= _state_T_1;
    end else begin
      state <= 2'h0;
    end
    if (reset) begin // @[EXU.scala 129:29]
      alu_wait <= 1'h0; // @[EXU.scala 129:29]
    end else begin
      alu_wait <= _lsu_io_ls_in_valid_T; // @[EXU.scala 130:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  EXE_reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  EXE_reg_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  EXE_reg_rs1 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  EXE_reg_rs2 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  EXE_reg_rd = _RAND_4[4:0];
  _RAND_5 = {2{`RANDOM}};
  EXE_reg_imm = _RAND_5[63:0];
  _RAND_6 = {3{`RANDOM}};
  EXE_reg_op = _RAND_6[79:0];
  _RAND_7 = {1{`RANDOM}};
  EXE_reg_typ = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  EXE_reg_isJump = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  EXE_reg_clearidx = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  lsu_finish = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  alu_finish = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  alu_wait = _RAND_13[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_pc,
  input  [63:0] io_in_bits_pc_dnpc,
  input  [4:0]  io_in_bits_gpr_idx_w,
  input         io_in_bits_gpr_en_w,
  input  [63:0] io_in_bits_gpr_val_w,
  input         io_in_bits_csr_en_w,
  input  [11:0] io_in_bits_csr_idx_w,
  input  [63:0] io_in_bits_csr_val_w,
  input  [63:0] io_in_bits_csr_no,
  input  [63:0] io_in_bits_csr_epc,
  input         io_in_bits_isJump,
  input  [4:0]  io_in_bits_clearidx,
  output [4:0]  io_gpr_idx_w,
  output        io_gpr_en_w,
  output [63:0] io_gpr_val_w,
  output        io_csr_en_w,
  output [11:0] io_csr_idx_w,
  output [63:0] io_csr_val_w,
  output [63:0] io_csr_no,
  output [63:0] io_csr_epc,
  output [63:0] io_pc_dnpc,
  output        io_valid,
  output        io_isJump,
  output [4:0]  io_sb_clearidx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  _WB_reg_pc_T = io_in_ready & io_in_valid; // @[Decoupled.scala 52:35]
  reg [31:0] WB_reg_pc; // @[Reg.scala 19:16]
  reg [31:0] WB_reg_pc_dnpc; // @[Reg.scala 35:20]
  wire [63:0] _GEN_2 = _WB_reg_pc_T ? io_in_bits_pc_dnpc : {{32'd0}, WB_reg_pc_dnpc}; // @[Reg.scala 36:18 35:20 36:22]
  reg  WB_reg_gpr_en_w; // @[Reg.scala 19:16]
  reg [4:0] WB_reg_gpr_idx_w; // @[Reg.scala 19:16]
  reg [63:0] WB_reg_gpr_val_w; // @[Reg.scala 19:16]
  reg  WB_reg_csr_en_w; // @[Reg.scala 19:16]
  reg [11:0] WB_reg_csr_idx_w; // @[Reg.scala 19:16]
  reg [63:0] WB_reg_csr_val_w; // @[Reg.scala 19:16]
  reg [63:0] WB_reg_csr_no; // @[Reg.scala 19:16]
  reg [63:0] WB_reg_csr_epc; // @[Reg.scala 19:16]
  reg  WB_reg_isJump; // @[Reg.scala 35:20]
  reg [4:0] WB_reg_clearidx; // @[Reg.scala 35:20]
  reg  state; // @[WBU.scala 32:24]
  wire [63:0] _GEN_14 = reset ? 64'h80000000 : _GEN_2; // @[Reg.scala 35:{20,20}]
  assign io_in_ready = ~state; // @[WBU.scala 39:25]
  assign io_gpr_idx_w = WB_reg_gpr_idx_w; // @[WBU.scala 42:17]
  assign io_gpr_en_w = WB_reg_gpr_en_w & state; // @[WBU.scala 41:34]
  assign io_gpr_val_w = WB_reg_gpr_val_w; // @[WBU.scala 43:17]
  assign io_csr_en_w = WB_reg_csr_en_w & state; // @[WBU.scala 45:34]
  assign io_csr_idx_w = WB_reg_csr_idx_w; // @[WBU.scala 46:17]
  assign io_csr_val_w = WB_reg_csr_val_w; // @[WBU.scala 47:17]
  assign io_csr_no = state ? WB_reg_csr_no : 64'h0; // @[WBU.scala 48:19]
  assign io_csr_epc = WB_reg_csr_epc; // @[WBU.scala 49:15]
  assign io_pc_dnpc = {{32'd0}, WB_reg_pc_dnpc}; // @[WBU.scala 51:15]
  assign io_valid = state; // @[WBU.scala 52:22]
  assign io_isJump = WB_reg_isJump & state; // @[WBU.scala 37:30]
  assign io_sb_clearidx = state ? WB_reg_clearidx : 5'h0; // @[WBU.scala 54:24]
  always @(posedge clock) begin
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_pc <= io_in_bits_pc; // @[Reg.scala 20:22]
    end
    WB_reg_pc_dnpc <= _GEN_14[31:0]; // @[Reg.scala 35:{20,20}]
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_gpr_en_w <= io_in_bits_gpr_en_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_gpr_idx_w <= io_in_bits_gpr_idx_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_gpr_val_w <= io_in_bits_gpr_val_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_csr_en_w <= io_in_bits_csr_en_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_csr_idx_w <= io_in_bits_csr_idx_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_csr_val_w <= io_in_bits_csr_val_w; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_csr_no <= io_in_bits_csr_no; // @[Reg.scala 20:22]
    end
    if (_WB_reg_pc_T) begin // @[Reg.scala 20:18]
      WB_reg_csr_epc <= io_in_bits_csr_epc; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      WB_reg_isJump <= 1'h0; // @[Reg.scala 35:20]
    end else if (_WB_reg_pc_T) begin // @[Reg.scala 36:18]
      WB_reg_isJump <= io_in_bits_isJump; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      WB_reg_clearidx <= 5'h0; // @[Reg.scala 35:20]
    end else if (_WB_reg_pc_T) begin // @[Reg.scala 36:18]
      WB_reg_clearidx <= io_in_bits_clearidx; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[WBU.scala 32:24]
      state <= 1'h0; // @[WBU.scala 32:24]
    end else if (state) begin // @[Mux.scala 81:58]
      state <= 1'h0;
    end else begin
      state <= _WB_reg_pc_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  WB_reg_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  WB_reg_pc_dnpc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  WB_reg_gpr_en_w = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  WB_reg_gpr_idx_w = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  WB_reg_gpr_val_w = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  WB_reg_csr_en_w = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  WB_reg_csr_idx_w = _RAND_6[11:0];
  _RAND_7 = {2{`RANDOM}};
  WB_reg_csr_val_w = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  WB_reg_csr_no = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  WB_reg_csr_epc = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  WB_reg_isJump = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  WB_reg_clearidx = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GPR(
  input         clock,
  input         reset,
  input  [4:0]  io_r_idx_r1,
  input  [4:0]  io_r_idx_r2,
  input         io_r_en_r1,
  input         io_r_en_r2,
  output [63:0] io_r_val_r1,
  output [63:0] io_r_val_r2,
  input  [4:0]  io_w_idx_w,
  input         io_w_en_w,
  input  [63:0] io_w_val_w
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] p_rf_0; // @[GPR.scala 31:17]
  wire [63:0] p_rf_1; // @[GPR.scala 31:17]
  wire [63:0] p_rf_2; // @[GPR.scala 31:17]
  wire [63:0] p_rf_3; // @[GPR.scala 31:17]
  wire [63:0] p_rf_4; // @[GPR.scala 31:17]
  wire [63:0] p_rf_5; // @[GPR.scala 31:17]
  wire [63:0] p_rf_6; // @[GPR.scala 31:17]
  wire [63:0] p_rf_7; // @[GPR.scala 31:17]
  wire [63:0] p_rf_8; // @[GPR.scala 31:17]
  wire [63:0] p_rf_9; // @[GPR.scala 31:17]
  wire [63:0] p_rf_10; // @[GPR.scala 31:17]
  wire [63:0] p_rf_11; // @[GPR.scala 31:17]
  wire [63:0] p_rf_12; // @[GPR.scala 31:17]
  wire [63:0] p_rf_13; // @[GPR.scala 31:17]
  wire [63:0] p_rf_14; // @[GPR.scala 31:17]
  wire [63:0] p_rf_15; // @[GPR.scala 31:17]
  wire [63:0] p_rf_16; // @[GPR.scala 31:17]
  wire [63:0] p_rf_17; // @[GPR.scala 31:17]
  wire [63:0] p_rf_18; // @[GPR.scala 31:17]
  wire [63:0] p_rf_19; // @[GPR.scala 31:17]
  wire [63:0] p_rf_20; // @[GPR.scala 31:17]
  wire [63:0] p_rf_21; // @[GPR.scala 31:17]
  wire [63:0] p_rf_22; // @[GPR.scala 31:17]
  wire [63:0] p_rf_23; // @[GPR.scala 31:17]
  wire [63:0] p_rf_24; // @[GPR.scala 31:17]
  wire [63:0] p_rf_25; // @[GPR.scala 31:17]
  wire [63:0] p_rf_26; // @[GPR.scala 31:17]
  wire [63:0] p_rf_27; // @[GPR.scala 31:17]
  wire [63:0] p_rf_28; // @[GPR.scala 31:17]
  wire [63:0] p_rf_29; // @[GPR.scala 31:17]
  wire [63:0] p_rf_30; // @[GPR.scala 31:17]
  wire [63:0] p_rf_31; // @[GPR.scala 31:17]
  reg [63:0] gpr_1; // @[GPR.scala 25:20]
  reg [63:0] gpr_2; // @[GPR.scala 25:20]
  reg [63:0] gpr_3; // @[GPR.scala 25:20]
  reg [63:0] gpr_4; // @[GPR.scala 25:20]
  reg [63:0] gpr_5; // @[GPR.scala 25:20]
  reg [63:0] gpr_6; // @[GPR.scala 25:20]
  reg [63:0] gpr_7; // @[GPR.scala 25:20]
  reg [63:0] gpr_8; // @[GPR.scala 25:20]
  reg [63:0] gpr_9; // @[GPR.scala 25:20]
  reg [63:0] gpr_10; // @[GPR.scala 25:20]
  reg [63:0] gpr_11; // @[GPR.scala 25:20]
  reg [63:0] gpr_12; // @[GPR.scala 25:20]
  reg [63:0] gpr_13; // @[GPR.scala 25:20]
  reg [63:0] gpr_14; // @[GPR.scala 25:20]
  reg [63:0] gpr_15; // @[GPR.scala 25:20]
  reg [63:0] gpr_16; // @[GPR.scala 25:20]
  reg [63:0] gpr_17; // @[GPR.scala 25:20]
  reg [63:0] gpr_18; // @[GPR.scala 25:20]
  reg [63:0] gpr_19; // @[GPR.scala 25:20]
  reg [63:0] gpr_20; // @[GPR.scala 25:20]
  reg [63:0] gpr_21; // @[GPR.scala 25:20]
  reg [63:0] gpr_22; // @[GPR.scala 25:20]
  reg [63:0] gpr_23; // @[GPR.scala 25:20]
  reg [63:0] gpr_24; // @[GPR.scala 25:20]
  reg [63:0] gpr_25; // @[GPR.scala 25:20]
  reg [63:0] gpr_26; // @[GPR.scala 25:20]
  reg [63:0] gpr_27; // @[GPR.scala 25:20]
  reg [63:0] gpr_28; // @[GPR.scala 25:20]
  reg [63:0] gpr_29; // @[GPR.scala 25:20]
  reg [63:0] gpr_30; // @[GPR.scala 25:20]
  reg [63:0] gpr_31; // @[GPR.scala 25:20]
  wire [63:0] _GEN_1 = 5'h1 == io_r_idx_r1 ? gpr_1 : 64'h0; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_2 = 5'h2 == io_r_idx_r1 ? gpr_2 : _GEN_1; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_3 = 5'h3 == io_r_idx_r1 ? gpr_3 : _GEN_2; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_4 = 5'h4 == io_r_idx_r1 ? gpr_4 : _GEN_3; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_5 = 5'h5 == io_r_idx_r1 ? gpr_5 : _GEN_4; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_6 = 5'h6 == io_r_idx_r1 ? gpr_6 : _GEN_5; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_7 = 5'h7 == io_r_idx_r1 ? gpr_7 : _GEN_6; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_8 = 5'h8 == io_r_idx_r1 ? gpr_8 : _GEN_7; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_9 = 5'h9 == io_r_idx_r1 ? gpr_9 : _GEN_8; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_10 = 5'ha == io_r_idx_r1 ? gpr_10 : _GEN_9; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_11 = 5'hb == io_r_idx_r1 ? gpr_11 : _GEN_10; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_12 = 5'hc == io_r_idx_r1 ? gpr_12 : _GEN_11; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_13 = 5'hd == io_r_idx_r1 ? gpr_13 : _GEN_12; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_14 = 5'he == io_r_idx_r1 ? gpr_14 : _GEN_13; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_15 = 5'hf == io_r_idx_r1 ? gpr_15 : _GEN_14; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_16 = 5'h10 == io_r_idx_r1 ? gpr_16 : _GEN_15; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_17 = 5'h11 == io_r_idx_r1 ? gpr_17 : _GEN_16; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_18 = 5'h12 == io_r_idx_r1 ? gpr_18 : _GEN_17; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_19 = 5'h13 == io_r_idx_r1 ? gpr_19 : _GEN_18; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_20 = 5'h14 == io_r_idx_r1 ? gpr_20 : _GEN_19; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_21 = 5'h15 == io_r_idx_r1 ? gpr_21 : _GEN_20; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_22 = 5'h16 == io_r_idx_r1 ? gpr_22 : _GEN_21; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_23 = 5'h17 == io_r_idx_r1 ? gpr_23 : _GEN_22; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_24 = 5'h18 == io_r_idx_r1 ? gpr_24 : _GEN_23; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_25 = 5'h19 == io_r_idx_r1 ? gpr_25 : _GEN_24; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_26 = 5'h1a == io_r_idx_r1 ? gpr_26 : _GEN_25; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_27 = 5'h1b == io_r_idx_r1 ? gpr_27 : _GEN_26; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_28 = 5'h1c == io_r_idx_r1 ? gpr_28 : _GEN_27; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_29 = 5'h1d == io_r_idx_r1 ? gpr_29 : _GEN_28; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_30 = 5'h1e == io_r_idx_r1 ? gpr_30 : _GEN_29; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_31 = 5'h1f == io_r_idx_r1 ? gpr_31 : _GEN_30; // @[GPR.scala 26:{21,21}]
  wire [63:0] _GEN_33 = 5'h1 == io_r_idx_r2 ? gpr_1 : 64'h0; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_34 = 5'h2 == io_r_idx_r2 ? gpr_2 : _GEN_33; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_35 = 5'h3 == io_r_idx_r2 ? gpr_3 : _GEN_34; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_36 = 5'h4 == io_r_idx_r2 ? gpr_4 : _GEN_35; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_37 = 5'h5 == io_r_idx_r2 ? gpr_5 : _GEN_36; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_38 = 5'h6 == io_r_idx_r2 ? gpr_6 : _GEN_37; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_39 = 5'h7 == io_r_idx_r2 ? gpr_7 : _GEN_38; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_40 = 5'h8 == io_r_idx_r2 ? gpr_8 : _GEN_39; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_41 = 5'h9 == io_r_idx_r2 ? gpr_9 : _GEN_40; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_42 = 5'ha == io_r_idx_r2 ? gpr_10 : _GEN_41; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_43 = 5'hb == io_r_idx_r2 ? gpr_11 : _GEN_42; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_44 = 5'hc == io_r_idx_r2 ? gpr_12 : _GEN_43; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_45 = 5'hd == io_r_idx_r2 ? gpr_13 : _GEN_44; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_46 = 5'he == io_r_idx_r2 ? gpr_14 : _GEN_45; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_47 = 5'hf == io_r_idx_r2 ? gpr_15 : _GEN_46; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_48 = 5'h10 == io_r_idx_r2 ? gpr_16 : _GEN_47; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_49 = 5'h11 == io_r_idx_r2 ? gpr_17 : _GEN_48; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_50 = 5'h12 == io_r_idx_r2 ? gpr_18 : _GEN_49; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_51 = 5'h13 == io_r_idx_r2 ? gpr_19 : _GEN_50; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_52 = 5'h14 == io_r_idx_r2 ? gpr_20 : _GEN_51; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_53 = 5'h15 == io_r_idx_r2 ? gpr_21 : _GEN_52; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_54 = 5'h16 == io_r_idx_r2 ? gpr_22 : _GEN_53; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_55 = 5'h17 == io_r_idx_r2 ? gpr_23 : _GEN_54; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_56 = 5'h18 == io_r_idx_r2 ? gpr_24 : _GEN_55; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_57 = 5'h19 == io_r_idx_r2 ? gpr_25 : _GEN_56; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_58 = 5'h1a == io_r_idx_r2 ? gpr_26 : _GEN_57; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_59 = 5'h1b == io_r_idx_r2 ? gpr_27 : _GEN_58; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_60 = 5'h1c == io_r_idx_r2 ? gpr_28 : _GEN_59; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_61 = 5'h1d == io_r_idx_r2 ? gpr_29 : _GEN_60; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_62 = 5'h1e == io_r_idx_r2 ? gpr_30 : _GEN_61; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_63 = 5'h1f == io_r_idx_r2 ? gpr_31 : _GEN_62; // @[GPR.scala 27:{21,21}]
  wire [63:0] _GEN_65 = 5'h1 == io_w_idx_w ? gpr_1 : 64'h0; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_66 = 5'h2 == io_w_idx_w ? gpr_2 : _GEN_65; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_67 = 5'h3 == io_w_idx_w ? gpr_3 : _GEN_66; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_68 = 5'h4 == io_w_idx_w ? gpr_4 : _GEN_67; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_69 = 5'h5 == io_w_idx_w ? gpr_5 : _GEN_68; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_70 = 5'h6 == io_w_idx_w ? gpr_6 : _GEN_69; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_71 = 5'h7 == io_w_idx_w ? gpr_7 : _GEN_70; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_72 = 5'h8 == io_w_idx_w ? gpr_8 : _GEN_71; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_73 = 5'h9 == io_w_idx_w ? gpr_9 : _GEN_72; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_74 = 5'ha == io_w_idx_w ? gpr_10 : _GEN_73; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_75 = 5'hb == io_w_idx_w ? gpr_11 : _GEN_74; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_76 = 5'hc == io_w_idx_w ? gpr_12 : _GEN_75; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_77 = 5'hd == io_w_idx_w ? gpr_13 : _GEN_76; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_78 = 5'he == io_w_idx_w ? gpr_14 : _GEN_77; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_79 = 5'hf == io_w_idx_w ? gpr_15 : _GEN_78; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_80 = 5'h10 == io_w_idx_w ? gpr_16 : _GEN_79; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_81 = 5'h11 == io_w_idx_w ? gpr_17 : _GEN_80; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_82 = 5'h12 == io_w_idx_w ? gpr_18 : _GEN_81; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_83 = 5'h13 == io_w_idx_w ? gpr_19 : _GEN_82; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_84 = 5'h14 == io_w_idx_w ? gpr_20 : _GEN_83; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_85 = 5'h15 == io_w_idx_w ? gpr_21 : _GEN_84; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_86 = 5'h16 == io_w_idx_w ? gpr_22 : _GEN_85; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_87 = 5'h17 == io_w_idx_w ? gpr_23 : _GEN_86; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_88 = 5'h18 == io_w_idx_w ? gpr_24 : _GEN_87; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_89 = 5'h19 == io_w_idx_w ? gpr_25 : _GEN_88; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_90 = 5'h1a == io_w_idx_w ? gpr_26 : _GEN_89; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_91 = 5'h1b == io_w_idx_w ? gpr_27 : _GEN_90; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_92 = 5'h1c == io_w_idx_w ? gpr_28 : _GEN_91; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_93 = 5'h1d == io_w_idx_w ? gpr_29 : _GEN_92; // @[GPR.scala 28:{25,25}]
  wire [63:0] _GEN_94 = 5'h1e == io_w_idx_w ? gpr_30 : _GEN_93; // @[GPR.scala 28:{25,25}]
  print_gpr p ( // @[GPR.scala 31:17]
    .rf_0(p_rf_0),
    .rf_1(p_rf_1),
    .rf_2(p_rf_2),
    .rf_3(p_rf_3),
    .rf_4(p_rf_4),
    .rf_5(p_rf_5),
    .rf_6(p_rf_6),
    .rf_7(p_rf_7),
    .rf_8(p_rf_8),
    .rf_9(p_rf_9),
    .rf_10(p_rf_10),
    .rf_11(p_rf_11),
    .rf_12(p_rf_12),
    .rf_13(p_rf_13),
    .rf_14(p_rf_14),
    .rf_15(p_rf_15),
    .rf_16(p_rf_16),
    .rf_17(p_rf_17),
    .rf_18(p_rf_18),
    .rf_19(p_rf_19),
    .rf_20(p_rf_20),
    .rf_21(p_rf_21),
    .rf_22(p_rf_22),
    .rf_23(p_rf_23),
    .rf_24(p_rf_24),
    .rf_25(p_rf_25),
    .rf_26(p_rf_26),
    .rf_27(p_rf_27),
    .rf_28(p_rf_28),
    .rf_29(p_rf_29),
    .rf_30(p_rf_30),
    .rf_31(p_rf_31)
  );
  assign io_r_val_r1 = io_r_en_r1 ? _GEN_31 : 64'h0; // @[GPR.scala 26:21]
  assign io_r_val_r2 = io_r_en_r2 ? _GEN_63 : 64'h0; // @[GPR.scala 27:21]
  assign p_rf_0 = 64'h0; // @[GPR.scala 32:12]
  assign p_rf_1 = gpr_1; // @[GPR.scala 32:12]
  assign p_rf_2 = gpr_2; // @[GPR.scala 32:12]
  assign p_rf_3 = gpr_3; // @[GPR.scala 32:12]
  assign p_rf_4 = gpr_4; // @[GPR.scala 32:12]
  assign p_rf_5 = gpr_5; // @[GPR.scala 32:12]
  assign p_rf_6 = gpr_6; // @[GPR.scala 32:12]
  assign p_rf_7 = gpr_7; // @[GPR.scala 32:12]
  assign p_rf_8 = gpr_8; // @[GPR.scala 32:12]
  assign p_rf_9 = gpr_9; // @[GPR.scala 32:12]
  assign p_rf_10 = gpr_10; // @[GPR.scala 32:12]
  assign p_rf_11 = gpr_11; // @[GPR.scala 32:12]
  assign p_rf_12 = gpr_12; // @[GPR.scala 32:12]
  assign p_rf_13 = gpr_13; // @[GPR.scala 32:12]
  assign p_rf_14 = gpr_14; // @[GPR.scala 32:12]
  assign p_rf_15 = gpr_15; // @[GPR.scala 32:12]
  assign p_rf_16 = gpr_16; // @[GPR.scala 32:12]
  assign p_rf_17 = gpr_17; // @[GPR.scala 32:12]
  assign p_rf_18 = gpr_18; // @[GPR.scala 32:12]
  assign p_rf_19 = gpr_19; // @[GPR.scala 32:12]
  assign p_rf_20 = gpr_20; // @[GPR.scala 32:12]
  assign p_rf_21 = gpr_21; // @[GPR.scala 32:12]
  assign p_rf_22 = gpr_22; // @[GPR.scala 32:12]
  assign p_rf_23 = gpr_23; // @[GPR.scala 32:12]
  assign p_rf_24 = gpr_24; // @[GPR.scala 32:12]
  assign p_rf_25 = gpr_25; // @[GPR.scala 32:12]
  assign p_rf_26 = gpr_26; // @[GPR.scala 32:12]
  assign p_rf_27 = gpr_27; // @[GPR.scala 32:12]
  assign p_rf_28 = gpr_28; // @[GPR.scala 32:12]
  assign p_rf_29 = gpr_29; // @[GPR.scala 32:12]
  assign p_rf_30 = gpr_30; // @[GPR.scala 32:12]
  assign p_rf_31 = gpr_31; // @[GPR.scala 32:12]
  always @(posedge clock) begin
    if (reset) begin // @[GPR.scala 25:20]
      gpr_1 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_1 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_1 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_1 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_2 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h2 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_2 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_2 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_2 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_3 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h3 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_3 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_3 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_3 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_4 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h4 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_4 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_4 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_4 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_5 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h5 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_5 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_5 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_5 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_6 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h6 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_6 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_6 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_6 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_7 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h7 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_7 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_7 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_7 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_8 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h8 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_8 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_8 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_8 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_9 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h9 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_9 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_9 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_9 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_10 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'ha == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_10 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_10 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_10 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_11 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'hb == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_11 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_11 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_11 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_12 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'hc == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_12 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_12 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_12 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_13 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'hd == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_13 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_13 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_13 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_14 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'he == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_14 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_14 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_14 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_15 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'hf == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_15 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_15 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_15 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_16 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h10 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_16 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_16 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_16 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_17 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h11 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_17 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_17 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_17 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_18 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h12 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_18 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_18 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_18 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_19 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h13 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_19 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_19 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_19 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_20 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h14 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_20 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_20 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_20 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_21 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h15 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_21 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_21 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_21 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_22 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h16 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_22 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_22 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_22 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_23 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h17 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_23 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_23 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_23 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_24 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h18 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_24 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_24 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_24 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_25 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h19 == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_25 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_25 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_25 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_26 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1a == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_26 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_26 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_26 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_27 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1b == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_27 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_27 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_27 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_28 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1c == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_28 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_28 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_28 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_29 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1d == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_29 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_29 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_29 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_30 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1e == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_30 <= io_w_val_w;
      end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:25]
        gpr_30 <= gpr_31; // @[GPR.scala 28:25]
      end else begin
        gpr_30 <= _GEN_94;
      end
    end
    if (reset) begin // @[GPR.scala 25:20]
      gpr_31 <= 64'h0; // @[GPR.scala 25:20]
    end else if (5'h1f == io_w_idx_w) begin // @[GPR.scala 28:20]
      if (io_w_en_w) begin // @[GPR.scala 28:25]
        gpr_31 <= io_w_val_w;
      end else if (!(5'h1f == io_w_idx_w)) begin // @[GPR.scala 28:25]
        gpr_31 <= _GEN_94;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  gpr_1 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  gpr_2 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  gpr_3 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  gpr_4 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  gpr_5 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  gpr_6 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  gpr_7 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  gpr_8 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  gpr_9 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  gpr_10 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  gpr_11 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  gpr_12 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  gpr_13 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  gpr_14 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  gpr_15 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  gpr_16 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  gpr_17 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  gpr_18 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  gpr_19 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  gpr_20 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  gpr_21 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  gpr_22 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  gpr_23 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  gpr_24 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  gpr_25 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  gpr_26 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  gpr_27 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  gpr_28 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  gpr_29 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  gpr_30 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  gpr_31 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [11:0] io_r_idx_r,
  input         io_r_en_r,
  output [63:0] io_r_val_r,
  input         io_w_en_w,
  input  [11:0] io_w_idx_w,
  input  [63:0] io_w_val_w,
  input  [63:0] io_w_no,
  input  [63:0] io_w_epc
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] p_rf_0; // @[CSR.scala 48:17]
  wire [63:0] p_rf_1; // @[CSR.scala 48:17]
  wire [63:0] p_rf_2; // @[CSR.scala 48:17]
  wire [63:0] p_rf_3; // @[CSR.scala 48:17]
  reg [63:0] csr_0; // @[CSR.scala 24:20]
  reg [63:0] csr_1; // @[CSR.scala 24:20]
  reg [63:0] csr_2; // @[CSR.scala 24:20]
  reg [63:0] csr_3; // @[CSR.scala 24:20]
  wire [1:0] _map_r_T_4 = io_r_idx_r == 12'h342 ? 2'h3 : 2'h0; // @[CSR.scala 31:15]
  wire [1:0] _map_r_T_5 = io_r_idx_r == 12'h341 ? 2'h2 : _map_r_T_4; // @[CSR.scala 30:15]
  wire [1:0] _map_r_T_6 = io_r_idx_r == 12'h305 ? 2'h1 : _map_r_T_5; // @[CSR.scala 29:15]
  wire [1:0] map_r = io_r_idx_r == 12'h300 ? 2'h0 : _map_r_T_6; // @[CSR.scala 28:15]
  wire [1:0] _map_w_T_4 = io_w_idx_w == 12'h342 ? 2'h3 : 2'h0; // @[CSR.scala 37:15]
  wire [1:0] _map_w_T_5 = io_w_idx_w == 12'h341 ? 2'h2 : _map_w_T_4; // @[CSR.scala 36:15]
  wire [1:0] _map_w_T_6 = io_w_idx_w == 12'h305 ? 2'h1 : _map_w_T_5; // @[CSR.scala 35:15]
  wire [1:0] map_w = io_w_idx_w == 12'h300 ? 2'h0 : _map_w_T_6; // @[CSR.scala 34:15]
  wire  _csr_2_T = io_w_no == 64'h1; // @[CSR.scala 40:24]
  wire [63:0] _GEN_1 = 2'h1 == map_r ? csr_1 : csr_0; // @[CSR.scala 44:{20,20}]
  wire [63:0] _GEN_2 = 2'h2 == map_r ? csr_2 : _GEN_1; // @[CSR.scala 44:{20,20}]
  wire [63:0] _GEN_3 = 2'h3 == map_r ? csr_3 : _GEN_2; // @[CSR.scala 44:{20,20}]
  wire [63:0] _io_r_val_r_T_3 = io_r_en_r ? _GEN_3 : 64'h0; // @[CSR.scala 44:20]
  wire [63:0] _io_r_val_r_T_4 = io_w_no == 64'h2 ? csr_2 : _io_r_val_r_T_3; // @[CSR.scala 43:20]
  wire [63:0] _GEN_5 = 2'h1 == map_w ? csr_1 : csr_0; // @[CSR.scala 46:{20,20}]
  wire [63:0] _GEN_6 = 2'h2 == map_w ? csr_2 : _GEN_5; // @[CSR.scala 46:{20,20}]
  print_csr p ( // @[CSR.scala 48:17]
    .rf_0(p_rf_0),
    .rf_1(p_rf_1),
    .rf_2(p_rf_2),
    .rf_3(p_rf_3)
  );
  assign io_r_val_r = _csr_2_T ? csr_1 : _io_r_val_r_T_4; // @[CSR.scala 42:20]
  assign p_rf_0 = csr_0; // @[CSR.scala 49:12]
  assign p_rf_1 = csr_1; // @[CSR.scala 49:12]
  assign p_rf_2 = csr_2; // @[CSR.scala 49:12]
  assign p_rf_3 = csr_3; // @[CSR.scala 49:12]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 24:20]
      csr_0 <= 64'ha00001800; // @[CSR.scala 24:20]
    end else if (2'h0 == map_w) begin // @[CSR.scala 46:15]
      if (io_w_en_w) begin // @[CSR.scala 46:20]
        csr_0 <= io_w_val_w;
      end else if (2'h3 == map_w) begin // @[CSR.scala 46:20]
        csr_0 <= csr_3; // @[CSR.scala 46:20]
      end else begin
        csr_0 <= _GEN_6;
      end
    end
    if (reset) begin // @[CSR.scala 24:20]
      csr_1 <= 64'h0; // @[CSR.scala 24:20]
    end else if (2'h1 == map_w) begin // @[CSR.scala 46:15]
      if (io_w_en_w) begin // @[CSR.scala 46:20]
        csr_1 <= io_w_val_w;
      end else if (2'h3 == map_w) begin // @[CSR.scala 46:20]
        csr_1 <= csr_3; // @[CSR.scala 46:20]
      end else begin
        csr_1 <= _GEN_6;
      end
    end
    if (reset) begin // @[CSR.scala 24:20]
      csr_2 <= 64'h0; // @[CSR.scala 24:20]
    end else if (2'h2 == map_w) begin // @[CSR.scala 46:15]
      if (io_w_en_w) begin // @[CSR.scala 46:20]
        csr_2 <= io_w_val_w;
      end else if (2'h3 == map_w) begin // @[CSR.scala 46:20]
        csr_2 <= csr_3; // @[CSR.scala 46:20]
      end else begin
        csr_2 <= _GEN_6;
      end
    end else if (io_w_no == 64'h1) begin // @[CSR.scala 40:16]
      csr_2 <= io_w_epc;
    end
    if (reset) begin // @[CSR.scala 24:20]
      csr_3 <= 64'h0; // @[CSR.scala 24:20]
    end else if (2'h3 == map_w) begin // @[CSR.scala 46:15]
      if (io_w_en_w) begin // @[CSR.scala 46:20]
        csr_3 <= io_w_val_w;
      end else if (!(2'h3 == map_w)) begin // @[CSR.scala 46:20]
        csr_3 <= _GEN_6;
      end
    end else if (_csr_2_T) begin // @[CSR.scala 41:16]
      csr_3 <= 64'hb;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  csr_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  csr_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  csr_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  csr_3 = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ScoreBoard(
  input        clock,
  input        reset,
  input  [4:0] io_ID_lookidx1,
  input  [4:0] io_ID_lookidx2,
  input  [4:0] io_ID_setidx,
  output       io_ID_isBusy,
  input  [4:0] io_WB_clearidx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] busy; // @[ScoreBoard.scala 21:21]
  wire [62:0] _busy_T = 63'h1 << io_WB_clearidx; // @[ScoreBoard.scala 23:38]
  wire [31:0] _busy_T_2 = ~_busy_T[31:0]; // @[ScoreBoard.scala 25:24]
  wire [31:0] _busy_T_3 = busy & _busy_T_2; // @[ScoreBoard.scala 25:22]
  wire [62:0] _busy_T_4 = 63'h1 << io_ID_setidx; // @[ScoreBoard.scala 23:38]
  wire [31:0] _busy_T_6 = _busy_T_3 | _busy_T_4[31:0]; // @[ScoreBoard.scala 25:49]
  wire [31:0] _busy_T_8 = {_busy_T_6[31:1],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _io_ID_isBusy_T = busy >> io_ID_lookidx1; // @[ScoreBoard.scala 26:23]
  wire [31:0] _io_ID_isBusy_T_2 = busy >> io_ID_lookidx2; // @[ScoreBoard.scala 26:44]
  assign io_ID_isBusy = _io_ID_isBusy_T[0] | _io_ID_isBusy_T_2[0]; // @[ScoreBoard.scala 26:39]
  always @(posedge clock) begin
    if (reset) begin // @[ScoreBoard.scala 21:21]
      busy <= 32'h0; // @[ScoreBoard.scala 21:21]
    end else begin
      busy <= _busy_T_8; // @[ScoreBoard.scala 25:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LFSR_8(
  input        clock,
  input        reset,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] x; // @[LFSR_8.scala 9:16]
  wire  _x_T_6 = x[4] ^ x[3] ^ x[2] ^ x[0]; // @[LFSR_8.scala 10:25]
  wire [7:0] _x_T_8 = {_x_T_6,x[7:1]}; // @[Cat.scala 33:92]
  assign io_out = x; // @[LFSR_8.scala 11:9]
  always @(posedge clock) begin
    if (reset) begin // @[LFSR_8.scala 9:16]
      x <= 8'h1; // @[LFSR_8.scala 9:16]
    end else begin
      x <= _x_T_8; // @[LFSR_8.scala 10:4]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache(
  input          clock,
  input          reset,
  output         io_in_ar_ready,
  input          io_in_ar_valid,
  input  [31:0]  io_in_ar_bits_addr,
  input          io_in_r_ready,
  output         io_in_r_valid,
  output [63:0]  io_in_r_bits_data,
  output         io_in_aw_ready,
  input          io_in_aw_valid,
  input  [31:0]  io_in_aw_bits_addr,
  output         io_in_w_ready,
  input          io_in_w_valid,
  input  [63:0]  io_in_w_bits_data,
  input  [7:0]   io_in_w_bits_strb,
  input          io_in_b_ready,
  output         io_in_b_valid,
  input          io_mem_ar_ready,
  output         io_mem_ar_valid,
  output [31:0]  io_mem_ar_bits_addr,
  output         io_mem_r_ready,
  input          io_mem_r_valid,
  input  [63:0]  io_mem_r_bits_data,
  input          io_mem_aw_ready,
  output         io_mem_aw_valid,
  output [31:0]  io_mem_aw_bits_addr,
  input          io_mem_w_ready,
  output         io_mem_w_valid,
  output [63:0]  io_mem_w_bits_data,
  output         io_mem_w_bits_last,
  output         io_mem_b_ready,
  input          io_mem_b_valid,
  input  [127:0] io_ram_bits_Q,
  output         io_ram_bits_CEN,
  output         io_ram_bits_WEN,
  output [127:0] io_ram_bits_BWEN,
  output [7:0]   io_ram_bits_A,
  output [127:0] io_ram_bits_D,
  output [63:0]  io_hitrate
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [127:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [127:0] _RAND_517;
  reg [127:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
`endif // RANDOMIZE_REG_INIT
  reg [41:0] cache_tag [0:127]; // @[cache.scala 24:30]
  wire  cache_tag_tag_read_MPORT_en; // @[cache.scala 24:30]
  wire [6:0] cache_tag_tag_read_MPORT_addr; // @[cache.scala 24:30]
  wire [41:0] cache_tag_tag_read_MPORT_data; // @[cache.scala 24:30]
  wire [41:0] cache_tag_MPORT_data; // @[cache.scala 24:30]
  wire [6:0] cache_tag_MPORT_addr; // @[cache.scala 24:30]
  wire  cache_tag_MPORT_mask; // @[cache.scala 24:30]
  wire  cache_tag_MPORT_en; // @[cache.scala 24:30]
  reg  cache_tag_tag_read_MPORT_en_pipe_0;
  reg [6:0] cache_tag_tag_read_MPORT_addr_pipe_0;
  wire  lfsr8_clock; // @[cache.scala 61:21]
  wire  lfsr8_reset; // @[cache.scala 61:21]
  wire [7:0] lfsr8_io_out; // @[cache.scala 61:21]
  reg  valid_0_0; // @[cache.scala 25:22]
  reg  valid_0_1; // @[cache.scala 25:22]
  reg  valid_1_0; // @[cache.scala 25:22]
  reg  valid_1_1; // @[cache.scala 25:22]
  reg  valid_2_0; // @[cache.scala 25:22]
  reg  valid_2_1; // @[cache.scala 25:22]
  reg  valid_3_0; // @[cache.scala 25:22]
  reg  valid_3_1; // @[cache.scala 25:22]
  reg  valid_4_0; // @[cache.scala 25:22]
  reg  valid_4_1; // @[cache.scala 25:22]
  reg  valid_5_0; // @[cache.scala 25:22]
  reg  valid_5_1; // @[cache.scala 25:22]
  reg  valid_6_0; // @[cache.scala 25:22]
  reg  valid_6_1; // @[cache.scala 25:22]
  reg  valid_7_0; // @[cache.scala 25:22]
  reg  valid_7_1; // @[cache.scala 25:22]
  reg  valid_8_0; // @[cache.scala 25:22]
  reg  valid_8_1; // @[cache.scala 25:22]
  reg  valid_9_0; // @[cache.scala 25:22]
  reg  valid_9_1; // @[cache.scala 25:22]
  reg  valid_10_0; // @[cache.scala 25:22]
  reg  valid_10_1; // @[cache.scala 25:22]
  reg  valid_11_0; // @[cache.scala 25:22]
  reg  valid_11_1; // @[cache.scala 25:22]
  reg  valid_12_0; // @[cache.scala 25:22]
  reg  valid_12_1; // @[cache.scala 25:22]
  reg  valid_13_0; // @[cache.scala 25:22]
  reg  valid_13_1; // @[cache.scala 25:22]
  reg  valid_14_0; // @[cache.scala 25:22]
  reg  valid_14_1; // @[cache.scala 25:22]
  reg  valid_15_0; // @[cache.scala 25:22]
  reg  valid_15_1; // @[cache.scala 25:22]
  reg  valid_16_0; // @[cache.scala 25:22]
  reg  valid_16_1; // @[cache.scala 25:22]
  reg  valid_17_0; // @[cache.scala 25:22]
  reg  valid_17_1; // @[cache.scala 25:22]
  reg  valid_18_0; // @[cache.scala 25:22]
  reg  valid_18_1; // @[cache.scala 25:22]
  reg  valid_19_0; // @[cache.scala 25:22]
  reg  valid_19_1; // @[cache.scala 25:22]
  reg  valid_20_0; // @[cache.scala 25:22]
  reg  valid_20_1; // @[cache.scala 25:22]
  reg  valid_21_0; // @[cache.scala 25:22]
  reg  valid_21_1; // @[cache.scala 25:22]
  reg  valid_22_0; // @[cache.scala 25:22]
  reg  valid_22_1; // @[cache.scala 25:22]
  reg  valid_23_0; // @[cache.scala 25:22]
  reg  valid_23_1; // @[cache.scala 25:22]
  reg  valid_24_0; // @[cache.scala 25:22]
  reg  valid_24_1; // @[cache.scala 25:22]
  reg  valid_25_0; // @[cache.scala 25:22]
  reg  valid_25_1; // @[cache.scala 25:22]
  reg  valid_26_0; // @[cache.scala 25:22]
  reg  valid_26_1; // @[cache.scala 25:22]
  reg  valid_27_0; // @[cache.scala 25:22]
  reg  valid_27_1; // @[cache.scala 25:22]
  reg  valid_28_0; // @[cache.scala 25:22]
  reg  valid_28_1; // @[cache.scala 25:22]
  reg  valid_29_0; // @[cache.scala 25:22]
  reg  valid_29_1; // @[cache.scala 25:22]
  reg  valid_30_0; // @[cache.scala 25:22]
  reg  valid_30_1; // @[cache.scala 25:22]
  reg  valid_31_0; // @[cache.scala 25:22]
  reg  valid_31_1; // @[cache.scala 25:22]
  reg  valid_32_0; // @[cache.scala 25:22]
  reg  valid_32_1; // @[cache.scala 25:22]
  reg  valid_33_0; // @[cache.scala 25:22]
  reg  valid_33_1; // @[cache.scala 25:22]
  reg  valid_34_0; // @[cache.scala 25:22]
  reg  valid_34_1; // @[cache.scala 25:22]
  reg  valid_35_0; // @[cache.scala 25:22]
  reg  valid_35_1; // @[cache.scala 25:22]
  reg  valid_36_0; // @[cache.scala 25:22]
  reg  valid_36_1; // @[cache.scala 25:22]
  reg  valid_37_0; // @[cache.scala 25:22]
  reg  valid_37_1; // @[cache.scala 25:22]
  reg  valid_38_0; // @[cache.scala 25:22]
  reg  valid_38_1; // @[cache.scala 25:22]
  reg  valid_39_0; // @[cache.scala 25:22]
  reg  valid_39_1; // @[cache.scala 25:22]
  reg  valid_40_0; // @[cache.scala 25:22]
  reg  valid_40_1; // @[cache.scala 25:22]
  reg  valid_41_0; // @[cache.scala 25:22]
  reg  valid_41_1; // @[cache.scala 25:22]
  reg  valid_42_0; // @[cache.scala 25:22]
  reg  valid_42_1; // @[cache.scala 25:22]
  reg  valid_43_0; // @[cache.scala 25:22]
  reg  valid_43_1; // @[cache.scala 25:22]
  reg  valid_44_0; // @[cache.scala 25:22]
  reg  valid_44_1; // @[cache.scala 25:22]
  reg  valid_45_0; // @[cache.scala 25:22]
  reg  valid_45_1; // @[cache.scala 25:22]
  reg  valid_46_0; // @[cache.scala 25:22]
  reg  valid_46_1; // @[cache.scala 25:22]
  reg  valid_47_0; // @[cache.scala 25:22]
  reg  valid_47_1; // @[cache.scala 25:22]
  reg  valid_48_0; // @[cache.scala 25:22]
  reg  valid_48_1; // @[cache.scala 25:22]
  reg  valid_49_0; // @[cache.scala 25:22]
  reg  valid_49_1; // @[cache.scala 25:22]
  reg  valid_50_0; // @[cache.scala 25:22]
  reg  valid_50_1; // @[cache.scala 25:22]
  reg  valid_51_0; // @[cache.scala 25:22]
  reg  valid_51_1; // @[cache.scala 25:22]
  reg  valid_52_0; // @[cache.scala 25:22]
  reg  valid_52_1; // @[cache.scala 25:22]
  reg  valid_53_0; // @[cache.scala 25:22]
  reg  valid_53_1; // @[cache.scala 25:22]
  reg  valid_54_0; // @[cache.scala 25:22]
  reg  valid_54_1; // @[cache.scala 25:22]
  reg  valid_55_0; // @[cache.scala 25:22]
  reg  valid_55_1; // @[cache.scala 25:22]
  reg  valid_56_0; // @[cache.scala 25:22]
  reg  valid_56_1; // @[cache.scala 25:22]
  reg  valid_57_0; // @[cache.scala 25:22]
  reg  valid_57_1; // @[cache.scala 25:22]
  reg  valid_58_0; // @[cache.scala 25:22]
  reg  valid_58_1; // @[cache.scala 25:22]
  reg  valid_59_0; // @[cache.scala 25:22]
  reg  valid_59_1; // @[cache.scala 25:22]
  reg  valid_60_0; // @[cache.scala 25:22]
  reg  valid_60_1; // @[cache.scala 25:22]
  reg  valid_61_0; // @[cache.scala 25:22]
  reg  valid_61_1; // @[cache.scala 25:22]
  reg  valid_62_0; // @[cache.scala 25:22]
  reg  valid_62_1; // @[cache.scala 25:22]
  reg  valid_63_0; // @[cache.scala 25:22]
  reg  valid_63_1; // @[cache.scala 25:22]
  reg  valid_64_0; // @[cache.scala 25:22]
  reg  valid_64_1; // @[cache.scala 25:22]
  reg  valid_65_0; // @[cache.scala 25:22]
  reg  valid_65_1; // @[cache.scala 25:22]
  reg  valid_66_0; // @[cache.scala 25:22]
  reg  valid_66_1; // @[cache.scala 25:22]
  reg  valid_67_0; // @[cache.scala 25:22]
  reg  valid_67_1; // @[cache.scala 25:22]
  reg  valid_68_0; // @[cache.scala 25:22]
  reg  valid_68_1; // @[cache.scala 25:22]
  reg  valid_69_0; // @[cache.scala 25:22]
  reg  valid_69_1; // @[cache.scala 25:22]
  reg  valid_70_0; // @[cache.scala 25:22]
  reg  valid_70_1; // @[cache.scala 25:22]
  reg  valid_71_0; // @[cache.scala 25:22]
  reg  valid_71_1; // @[cache.scala 25:22]
  reg  valid_72_0; // @[cache.scala 25:22]
  reg  valid_72_1; // @[cache.scala 25:22]
  reg  valid_73_0; // @[cache.scala 25:22]
  reg  valid_73_1; // @[cache.scala 25:22]
  reg  valid_74_0; // @[cache.scala 25:22]
  reg  valid_74_1; // @[cache.scala 25:22]
  reg  valid_75_0; // @[cache.scala 25:22]
  reg  valid_75_1; // @[cache.scala 25:22]
  reg  valid_76_0; // @[cache.scala 25:22]
  reg  valid_76_1; // @[cache.scala 25:22]
  reg  valid_77_0; // @[cache.scala 25:22]
  reg  valid_77_1; // @[cache.scala 25:22]
  reg  valid_78_0; // @[cache.scala 25:22]
  reg  valid_78_1; // @[cache.scala 25:22]
  reg  valid_79_0; // @[cache.scala 25:22]
  reg  valid_79_1; // @[cache.scala 25:22]
  reg  valid_80_0; // @[cache.scala 25:22]
  reg  valid_80_1; // @[cache.scala 25:22]
  reg  valid_81_0; // @[cache.scala 25:22]
  reg  valid_81_1; // @[cache.scala 25:22]
  reg  valid_82_0; // @[cache.scala 25:22]
  reg  valid_82_1; // @[cache.scala 25:22]
  reg  valid_83_0; // @[cache.scala 25:22]
  reg  valid_83_1; // @[cache.scala 25:22]
  reg  valid_84_0; // @[cache.scala 25:22]
  reg  valid_84_1; // @[cache.scala 25:22]
  reg  valid_85_0; // @[cache.scala 25:22]
  reg  valid_85_1; // @[cache.scala 25:22]
  reg  valid_86_0; // @[cache.scala 25:22]
  reg  valid_86_1; // @[cache.scala 25:22]
  reg  valid_87_0; // @[cache.scala 25:22]
  reg  valid_87_1; // @[cache.scala 25:22]
  reg  valid_88_0; // @[cache.scala 25:22]
  reg  valid_88_1; // @[cache.scala 25:22]
  reg  valid_89_0; // @[cache.scala 25:22]
  reg  valid_89_1; // @[cache.scala 25:22]
  reg  valid_90_0; // @[cache.scala 25:22]
  reg  valid_90_1; // @[cache.scala 25:22]
  reg  valid_91_0; // @[cache.scala 25:22]
  reg  valid_91_1; // @[cache.scala 25:22]
  reg  valid_92_0; // @[cache.scala 25:22]
  reg  valid_92_1; // @[cache.scala 25:22]
  reg  valid_93_0; // @[cache.scala 25:22]
  reg  valid_93_1; // @[cache.scala 25:22]
  reg  valid_94_0; // @[cache.scala 25:22]
  reg  valid_94_1; // @[cache.scala 25:22]
  reg  valid_95_0; // @[cache.scala 25:22]
  reg  valid_95_1; // @[cache.scala 25:22]
  reg  valid_96_0; // @[cache.scala 25:22]
  reg  valid_96_1; // @[cache.scala 25:22]
  reg  valid_97_0; // @[cache.scala 25:22]
  reg  valid_97_1; // @[cache.scala 25:22]
  reg  valid_98_0; // @[cache.scala 25:22]
  reg  valid_98_1; // @[cache.scala 25:22]
  reg  valid_99_0; // @[cache.scala 25:22]
  reg  valid_99_1; // @[cache.scala 25:22]
  reg  valid_100_0; // @[cache.scala 25:22]
  reg  valid_100_1; // @[cache.scala 25:22]
  reg  valid_101_0; // @[cache.scala 25:22]
  reg  valid_101_1; // @[cache.scala 25:22]
  reg  valid_102_0; // @[cache.scala 25:22]
  reg  valid_102_1; // @[cache.scala 25:22]
  reg  valid_103_0; // @[cache.scala 25:22]
  reg  valid_103_1; // @[cache.scala 25:22]
  reg  valid_104_0; // @[cache.scala 25:22]
  reg  valid_104_1; // @[cache.scala 25:22]
  reg  valid_105_0; // @[cache.scala 25:22]
  reg  valid_105_1; // @[cache.scala 25:22]
  reg  valid_106_0; // @[cache.scala 25:22]
  reg  valid_106_1; // @[cache.scala 25:22]
  reg  valid_107_0; // @[cache.scala 25:22]
  reg  valid_107_1; // @[cache.scala 25:22]
  reg  valid_108_0; // @[cache.scala 25:22]
  reg  valid_108_1; // @[cache.scala 25:22]
  reg  valid_109_0; // @[cache.scala 25:22]
  reg  valid_109_1; // @[cache.scala 25:22]
  reg  valid_110_0; // @[cache.scala 25:22]
  reg  valid_110_1; // @[cache.scala 25:22]
  reg  valid_111_0; // @[cache.scala 25:22]
  reg  valid_111_1; // @[cache.scala 25:22]
  reg  valid_112_0; // @[cache.scala 25:22]
  reg  valid_112_1; // @[cache.scala 25:22]
  reg  valid_113_0; // @[cache.scala 25:22]
  reg  valid_113_1; // @[cache.scala 25:22]
  reg  valid_114_0; // @[cache.scala 25:22]
  reg  valid_114_1; // @[cache.scala 25:22]
  reg  valid_115_0; // @[cache.scala 25:22]
  reg  valid_115_1; // @[cache.scala 25:22]
  reg  valid_116_0; // @[cache.scala 25:22]
  reg  valid_116_1; // @[cache.scala 25:22]
  reg  valid_117_0; // @[cache.scala 25:22]
  reg  valid_117_1; // @[cache.scala 25:22]
  reg  valid_118_0; // @[cache.scala 25:22]
  reg  valid_118_1; // @[cache.scala 25:22]
  reg  valid_119_0; // @[cache.scala 25:22]
  reg  valid_119_1; // @[cache.scala 25:22]
  reg  valid_120_0; // @[cache.scala 25:22]
  reg  valid_120_1; // @[cache.scala 25:22]
  reg  valid_121_0; // @[cache.scala 25:22]
  reg  valid_121_1; // @[cache.scala 25:22]
  reg  valid_122_0; // @[cache.scala 25:22]
  reg  valid_122_1; // @[cache.scala 25:22]
  reg  valid_123_0; // @[cache.scala 25:22]
  reg  valid_123_1; // @[cache.scala 25:22]
  reg  valid_124_0; // @[cache.scala 25:22]
  reg  valid_124_1; // @[cache.scala 25:22]
  reg  valid_125_0; // @[cache.scala 25:22]
  reg  valid_125_1; // @[cache.scala 25:22]
  reg  valid_126_0; // @[cache.scala 25:22]
  reg  valid_126_1; // @[cache.scala 25:22]
  reg  valid_127_0; // @[cache.scala 25:22]
  reg  valid_127_1; // @[cache.scala 25:22]
  reg  dirty_0_0; // @[cache.scala 26:22]
  reg  dirty_0_1; // @[cache.scala 26:22]
  reg  dirty_1_0; // @[cache.scala 26:22]
  reg  dirty_1_1; // @[cache.scala 26:22]
  reg  dirty_2_0; // @[cache.scala 26:22]
  reg  dirty_2_1; // @[cache.scala 26:22]
  reg  dirty_3_0; // @[cache.scala 26:22]
  reg  dirty_3_1; // @[cache.scala 26:22]
  reg  dirty_4_0; // @[cache.scala 26:22]
  reg  dirty_4_1; // @[cache.scala 26:22]
  reg  dirty_5_0; // @[cache.scala 26:22]
  reg  dirty_5_1; // @[cache.scala 26:22]
  reg  dirty_6_0; // @[cache.scala 26:22]
  reg  dirty_6_1; // @[cache.scala 26:22]
  reg  dirty_7_0; // @[cache.scala 26:22]
  reg  dirty_7_1; // @[cache.scala 26:22]
  reg  dirty_8_0; // @[cache.scala 26:22]
  reg  dirty_8_1; // @[cache.scala 26:22]
  reg  dirty_9_0; // @[cache.scala 26:22]
  reg  dirty_9_1; // @[cache.scala 26:22]
  reg  dirty_10_0; // @[cache.scala 26:22]
  reg  dirty_10_1; // @[cache.scala 26:22]
  reg  dirty_11_0; // @[cache.scala 26:22]
  reg  dirty_11_1; // @[cache.scala 26:22]
  reg  dirty_12_0; // @[cache.scala 26:22]
  reg  dirty_12_1; // @[cache.scala 26:22]
  reg  dirty_13_0; // @[cache.scala 26:22]
  reg  dirty_13_1; // @[cache.scala 26:22]
  reg  dirty_14_0; // @[cache.scala 26:22]
  reg  dirty_14_1; // @[cache.scala 26:22]
  reg  dirty_15_0; // @[cache.scala 26:22]
  reg  dirty_15_1; // @[cache.scala 26:22]
  reg  dirty_16_0; // @[cache.scala 26:22]
  reg  dirty_16_1; // @[cache.scala 26:22]
  reg  dirty_17_0; // @[cache.scala 26:22]
  reg  dirty_17_1; // @[cache.scala 26:22]
  reg  dirty_18_0; // @[cache.scala 26:22]
  reg  dirty_18_1; // @[cache.scala 26:22]
  reg  dirty_19_0; // @[cache.scala 26:22]
  reg  dirty_19_1; // @[cache.scala 26:22]
  reg  dirty_20_0; // @[cache.scala 26:22]
  reg  dirty_20_1; // @[cache.scala 26:22]
  reg  dirty_21_0; // @[cache.scala 26:22]
  reg  dirty_21_1; // @[cache.scala 26:22]
  reg  dirty_22_0; // @[cache.scala 26:22]
  reg  dirty_22_1; // @[cache.scala 26:22]
  reg  dirty_23_0; // @[cache.scala 26:22]
  reg  dirty_23_1; // @[cache.scala 26:22]
  reg  dirty_24_0; // @[cache.scala 26:22]
  reg  dirty_24_1; // @[cache.scala 26:22]
  reg  dirty_25_0; // @[cache.scala 26:22]
  reg  dirty_25_1; // @[cache.scala 26:22]
  reg  dirty_26_0; // @[cache.scala 26:22]
  reg  dirty_26_1; // @[cache.scala 26:22]
  reg  dirty_27_0; // @[cache.scala 26:22]
  reg  dirty_27_1; // @[cache.scala 26:22]
  reg  dirty_28_0; // @[cache.scala 26:22]
  reg  dirty_28_1; // @[cache.scala 26:22]
  reg  dirty_29_0; // @[cache.scala 26:22]
  reg  dirty_29_1; // @[cache.scala 26:22]
  reg  dirty_30_0; // @[cache.scala 26:22]
  reg  dirty_30_1; // @[cache.scala 26:22]
  reg  dirty_31_0; // @[cache.scala 26:22]
  reg  dirty_31_1; // @[cache.scala 26:22]
  reg  dirty_32_0; // @[cache.scala 26:22]
  reg  dirty_32_1; // @[cache.scala 26:22]
  reg  dirty_33_0; // @[cache.scala 26:22]
  reg  dirty_33_1; // @[cache.scala 26:22]
  reg  dirty_34_0; // @[cache.scala 26:22]
  reg  dirty_34_1; // @[cache.scala 26:22]
  reg  dirty_35_0; // @[cache.scala 26:22]
  reg  dirty_35_1; // @[cache.scala 26:22]
  reg  dirty_36_0; // @[cache.scala 26:22]
  reg  dirty_36_1; // @[cache.scala 26:22]
  reg  dirty_37_0; // @[cache.scala 26:22]
  reg  dirty_37_1; // @[cache.scala 26:22]
  reg  dirty_38_0; // @[cache.scala 26:22]
  reg  dirty_38_1; // @[cache.scala 26:22]
  reg  dirty_39_0; // @[cache.scala 26:22]
  reg  dirty_39_1; // @[cache.scala 26:22]
  reg  dirty_40_0; // @[cache.scala 26:22]
  reg  dirty_40_1; // @[cache.scala 26:22]
  reg  dirty_41_0; // @[cache.scala 26:22]
  reg  dirty_41_1; // @[cache.scala 26:22]
  reg  dirty_42_0; // @[cache.scala 26:22]
  reg  dirty_42_1; // @[cache.scala 26:22]
  reg  dirty_43_0; // @[cache.scala 26:22]
  reg  dirty_43_1; // @[cache.scala 26:22]
  reg  dirty_44_0; // @[cache.scala 26:22]
  reg  dirty_44_1; // @[cache.scala 26:22]
  reg  dirty_45_0; // @[cache.scala 26:22]
  reg  dirty_45_1; // @[cache.scala 26:22]
  reg  dirty_46_0; // @[cache.scala 26:22]
  reg  dirty_46_1; // @[cache.scala 26:22]
  reg  dirty_47_0; // @[cache.scala 26:22]
  reg  dirty_47_1; // @[cache.scala 26:22]
  reg  dirty_48_0; // @[cache.scala 26:22]
  reg  dirty_48_1; // @[cache.scala 26:22]
  reg  dirty_49_0; // @[cache.scala 26:22]
  reg  dirty_49_1; // @[cache.scala 26:22]
  reg  dirty_50_0; // @[cache.scala 26:22]
  reg  dirty_50_1; // @[cache.scala 26:22]
  reg  dirty_51_0; // @[cache.scala 26:22]
  reg  dirty_51_1; // @[cache.scala 26:22]
  reg  dirty_52_0; // @[cache.scala 26:22]
  reg  dirty_52_1; // @[cache.scala 26:22]
  reg  dirty_53_0; // @[cache.scala 26:22]
  reg  dirty_53_1; // @[cache.scala 26:22]
  reg  dirty_54_0; // @[cache.scala 26:22]
  reg  dirty_54_1; // @[cache.scala 26:22]
  reg  dirty_55_0; // @[cache.scala 26:22]
  reg  dirty_55_1; // @[cache.scala 26:22]
  reg  dirty_56_0; // @[cache.scala 26:22]
  reg  dirty_56_1; // @[cache.scala 26:22]
  reg  dirty_57_0; // @[cache.scala 26:22]
  reg  dirty_57_1; // @[cache.scala 26:22]
  reg  dirty_58_0; // @[cache.scala 26:22]
  reg  dirty_58_1; // @[cache.scala 26:22]
  reg  dirty_59_0; // @[cache.scala 26:22]
  reg  dirty_59_1; // @[cache.scala 26:22]
  reg  dirty_60_0; // @[cache.scala 26:22]
  reg  dirty_60_1; // @[cache.scala 26:22]
  reg  dirty_61_0; // @[cache.scala 26:22]
  reg  dirty_61_1; // @[cache.scala 26:22]
  reg  dirty_62_0; // @[cache.scala 26:22]
  reg  dirty_62_1; // @[cache.scala 26:22]
  reg  dirty_63_0; // @[cache.scala 26:22]
  reg  dirty_63_1; // @[cache.scala 26:22]
  reg  dirty_64_0; // @[cache.scala 26:22]
  reg  dirty_64_1; // @[cache.scala 26:22]
  reg  dirty_65_0; // @[cache.scala 26:22]
  reg  dirty_65_1; // @[cache.scala 26:22]
  reg  dirty_66_0; // @[cache.scala 26:22]
  reg  dirty_66_1; // @[cache.scala 26:22]
  reg  dirty_67_0; // @[cache.scala 26:22]
  reg  dirty_67_1; // @[cache.scala 26:22]
  reg  dirty_68_0; // @[cache.scala 26:22]
  reg  dirty_68_1; // @[cache.scala 26:22]
  reg  dirty_69_0; // @[cache.scala 26:22]
  reg  dirty_69_1; // @[cache.scala 26:22]
  reg  dirty_70_0; // @[cache.scala 26:22]
  reg  dirty_70_1; // @[cache.scala 26:22]
  reg  dirty_71_0; // @[cache.scala 26:22]
  reg  dirty_71_1; // @[cache.scala 26:22]
  reg  dirty_72_0; // @[cache.scala 26:22]
  reg  dirty_72_1; // @[cache.scala 26:22]
  reg  dirty_73_0; // @[cache.scala 26:22]
  reg  dirty_73_1; // @[cache.scala 26:22]
  reg  dirty_74_0; // @[cache.scala 26:22]
  reg  dirty_74_1; // @[cache.scala 26:22]
  reg  dirty_75_0; // @[cache.scala 26:22]
  reg  dirty_75_1; // @[cache.scala 26:22]
  reg  dirty_76_0; // @[cache.scala 26:22]
  reg  dirty_76_1; // @[cache.scala 26:22]
  reg  dirty_77_0; // @[cache.scala 26:22]
  reg  dirty_77_1; // @[cache.scala 26:22]
  reg  dirty_78_0; // @[cache.scala 26:22]
  reg  dirty_78_1; // @[cache.scala 26:22]
  reg  dirty_79_0; // @[cache.scala 26:22]
  reg  dirty_79_1; // @[cache.scala 26:22]
  reg  dirty_80_0; // @[cache.scala 26:22]
  reg  dirty_80_1; // @[cache.scala 26:22]
  reg  dirty_81_0; // @[cache.scala 26:22]
  reg  dirty_81_1; // @[cache.scala 26:22]
  reg  dirty_82_0; // @[cache.scala 26:22]
  reg  dirty_82_1; // @[cache.scala 26:22]
  reg  dirty_83_0; // @[cache.scala 26:22]
  reg  dirty_83_1; // @[cache.scala 26:22]
  reg  dirty_84_0; // @[cache.scala 26:22]
  reg  dirty_84_1; // @[cache.scala 26:22]
  reg  dirty_85_0; // @[cache.scala 26:22]
  reg  dirty_85_1; // @[cache.scala 26:22]
  reg  dirty_86_0; // @[cache.scala 26:22]
  reg  dirty_86_1; // @[cache.scala 26:22]
  reg  dirty_87_0; // @[cache.scala 26:22]
  reg  dirty_87_1; // @[cache.scala 26:22]
  reg  dirty_88_0; // @[cache.scala 26:22]
  reg  dirty_88_1; // @[cache.scala 26:22]
  reg  dirty_89_0; // @[cache.scala 26:22]
  reg  dirty_89_1; // @[cache.scala 26:22]
  reg  dirty_90_0; // @[cache.scala 26:22]
  reg  dirty_90_1; // @[cache.scala 26:22]
  reg  dirty_91_0; // @[cache.scala 26:22]
  reg  dirty_91_1; // @[cache.scala 26:22]
  reg  dirty_92_0; // @[cache.scala 26:22]
  reg  dirty_92_1; // @[cache.scala 26:22]
  reg  dirty_93_0; // @[cache.scala 26:22]
  reg  dirty_93_1; // @[cache.scala 26:22]
  reg  dirty_94_0; // @[cache.scala 26:22]
  reg  dirty_94_1; // @[cache.scala 26:22]
  reg  dirty_95_0; // @[cache.scala 26:22]
  reg  dirty_95_1; // @[cache.scala 26:22]
  reg  dirty_96_0; // @[cache.scala 26:22]
  reg  dirty_96_1; // @[cache.scala 26:22]
  reg  dirty_97_0; // @[cache.scala 26:22]
  reg  dirty_97_1; // @[cache.scala 26:22]
  reg  dirty_98_0; // @[cache.scala 26:22]
  reg  dirty_98_1; // @[cache.scala 26:22]
  reg  dirty_99_0; // @[cache.scala 26:22]
  reg  dirty_99_1; // @[cache.scala 26:22]
  reg  dirty_100_0; // @[cache.scala 26:22]
  reg  dirty_100_1; // @[cache.scala 26:22]
  reg  dirty_101_0; // @[cache.scala 26:22]
  reg  dirty_101_1; // @[cache.scala 26:22]
  reg  dirty_102_0; // @[cache.scala 26:22]
  reg  dirty_102_1; // @[cache.scala 26:22]
  reg  dirty_103_0; // @[cache.scala 26:22]
  reg  dirty_103_1; // @[cache.scala 26:22]
  reg  dirty_104_0; // @[cache.scala 26:22]
  reg  dirty_104_1; // @[cache.scala 26:22]
  reg  dirty_105_0; // @[cache.scala 26:22]
  reg  dirty_105_1; // @[cache.scala 26:22]
  reg  dirty_106_0; // @[cache.scala 26:22]
  reg  dirty_106_1; // @[cache.scala 26:22]
  reg  dirty_107_0; // @[cache.scala 26:22]
  reg  dirty_107_1; // @[cache.scala 26:22]
  reg  dirty_108_0; // @[cache.scala 26:22]
  reg  dirty_108_1; // @[cache.scala 26:22]
  reg  dirty_109_0; // @[cache.scala 26:22]
  reg  dirty_109_1; // @[cache.scala 26:22]
  reg  dirty_110_0; // @[cache.scala 26:22]
  reg  dirty_110_1; // @[cache.scala 26:22]
  reg  dirty_111_0; // @[cache.scala 26:22]
  reg  dirty_111_1; // @[cache.scala 26:22]
  reg  dirty_112_0; // @[cache.scala 26:22]
  reg  dirty_112_1; // @[cache.scala 26:22]
  reg  dirty_113_0; // @[cache.scala 26:22]
  reg  dirty_113_1; // @[cache.scala 26:22]
  reg  dirty_114_0; // @[cache.scala 26:22]
  reg  dirty_114_1; // @[cache.scala 26:22]
  reg  dirty_115_0; // @[cache.scala 26:22]
  reg  dirty_115_1; // @[cache.scala 26:22]
  reg  dirty_116_0; // @[cache.scala 26:22]
  reg  dirty_116_1; // @[cache.scala 26:22]
  reg  dirty_117_0; // @[cache.scala 26:22]
  reg  dirty_117_1; // @[cache.scala 26:22]
  reg  dirty_118_0; // @[cache.scala 26:22]
  reg  dirty_118_1; // @[cache.scala 26:22]
  reg  dirty_119_0; // @[cache.scala 26:22]
  reg  dirty_119_1; // @[cache.scala 26:22]
  reg  dirty_120_0; // @[cache.scala 26:22]
  reg  dirty_120_1; // @[cache.scala 26:22]
  reg  dirty_121_0; // @[cache.scala 26:22]
  reg  dirty_121_1; // @[cache.scala 26:22]
  reg  dirty_122_0; // @[cache.scala 26:22]
  reg  dirty_122_1; // @[cache.scala 26:22]
  reg  dirty_123_0; // @[cache.scala 26:22]
  reg  dirty_123_1; // @[cache.scala 26:22]
  reg  dirty_124_0; // @[cache.scala 26:22]
  reg  dirty_124_1; // @[cache.scala 26:22]
  reg  dirty_125_0; // @[cache.scala 26:22]
  reg  dirty_125_1; // @[cache.scala 26:22]
  reg  dirty_126_0; // @[cache.scala 26:22]
  reg  dirty_126_1; // @[cache.scala 26:22]
  reg  dirty_127_0; // @[cache.scala 26:22]
  reg  dirty_127_1; // @[cache.scala 26:22]
  reg [127:0] buf_; // @[cache.scala 27:20]
  reg [31:0] addr; // @[cache.scala 29:21]
  reg [127:0] wdata; // @[cache.scala 30:22]
  reg [127:0] wstrb; // @[cache.scala 31:22]
  wire [6:0] offset = {addr[3:0], 3'h0}; // @[cache.scala 32:42]
  wire [6:0] idx = addr[10:4]; // @[cache.scala 33:17]
  wire [20:0] tag = addr[31:11]; // @[cache.scala 34:17]
  reg [7:0] way2; // @[cache.scala 37:21]
  reg [3:0] state; // @[cache.scala 40:22]
  reg [3:0] state_r; // @[cache.scala 41:24]
  reg [3:0] state_w; // @[cache.scala 42:24]
  wire [7:0] _idxh_T = {idx, 1'h0}; // @[cache.scala 44:18]
  wire [41:0] tag_read = cache_tag_tag_read_MPORT_data; // @[cache.scala 56:22 57:12]
  wire  _GEN_5 = 7'h1 == idx ? valid_1_0 : valid_0_0; // @[cache.scala 58:{66,66}]
  wire  _GEN_6 = 7'h2 == idx ? valid_2_0 : _GEN_5; // @[cache.scala 58:{66,66}]
  wire  _GEN_7 = 7'h3 == idx ? valid_3_0 : _GEN_6; // @[cache.scala 58:{66,66}]
  wire  _GEN_8 = 7'h4 == idx ? valid_4_0 : _GEN_7; // @[cache.scala 58:{66,66}]
  wire  _GEN_9 = 7'h5 == idx ? valid_5_0 : _GEN_8; // @[cache.scala 58:{66,66}]
  wire  _GEN_10 = 7'h6 == idx ? valid_6_0 : _GEN_9; // @[cache.scala 58:{66,66}]
  wire  _GEN_11 = 7'h7 == idx ? valid_7_0 : _GEN_10; // @[cache.scala 58:{66,66}]
  wire  _GEN_12 = 7'h8 == idx ? valid_8_0 : _GEN_11; // @[cache.scala 58:{66,66}]
  wire  _GEN_13 = 7'h9 == idx ? valid_9_0 : _GEN_12; // @[cache.scala 58:{66,66}]
  wire  _GEN_14 = 7'ha == idx ? valid_10_0 : _GEN_13; // @[cache.scala 58:{66,66}]
  wire  _GEN_15 = 7'hb == idx ? valid_11_0 : _GEN_14; // @[cache.scala 58:{66,66}]
  wire  _GEN_16 = 7'hc == idx ? valid_12_0 : _GEN_15; // @[cache.scala 58:{66,66}]
  wire  _GEN_17 = 7'hd == idx ? valid_13_0 : _GEN_16; // @[cache.scala 58:{66,66}]
  wire  _GEN_18 = 7'he == idx ? valid_14_0 : _GEN_17; // @[cache.scala 58:{66,66}]
  wire  _GEN_19 = 7'hf == idx ? valid_15_0 : _GEN_18; // @[cache.scala 58:{66,66}]
  wire  _GEN_20 = 7'h10 == idx ? valid_16_0 : _GEN_19; // @[cache.scala 58:{66,66}]
  wire  _GEN_21 = 7'h11 == idx ? valid_17_0 : _GEN_20; // @[cache.scala 58:{66,66}]
  wire  _GEN_22 = 7'h12 == idx ? valid_18_0 : _GEN_21; // @[cache.scala 58:{66,66}]
  wire  _GEN_23 = 7'h13 == idx ? valid_19_0 : _GEN_22; // @[cache.scala 58:{66,66}]
  wire  _GEN_24 = 7'h14 == idx ? valid_20_0 : _GEN_23; // @[cache.scala 58:{66,66}]
  wire  _GEN_25 = 7'h15 == idx ? valid_21_0 : _GEN_24; // @[cache.scala 58:{66,66}]
  wire  _GEN_26 = 7'h16 == idx ? valid_22_0 : _GEN_25; // @[cache.scala 58:{66,66}]
  wire  _GEN_27 = 7'h17 == idx ? valid_23_0 : _GEN_26; // @[cache.scala 58:{66,66}]
  wire  _GEN_28 = 7'h18 == idx ? valid_24_0 : _GEN_27; // @[cache.scala 58:{66,66}]
  wire  _GEN_29 = 7'h19 == idx ? valid_25_0 : _GEN_28; // @[cache.scala 58:{66,66}]
  wire  _GEN_30 = 7'h1a == idx ? valid_26_0 : _GEN_29; // @[cache.scala 58:{66,66}]
  wire  _GEN_31 = 7'h1b == idx ? valid_27_0 : _GEN_30; // @[cache.scala 58:{66,66}]
  wire  _GEN_32 = 7'h1c == idx ? valid_28_0 : _GEN_31; // @[cache.scala 58:{66,66}]
  wire  _GEN_33 = 7'h1d == idx ? valid_29_0 : _GEN_32; // @[cache.scala 58:{66,66}]
  wire  _GEN_34 = 7'h1e == idx ? valid_30_0 : _GEN_33; // @[cache.scala 58:{66,66}]
  wire  _GEN_35 = 7'h1f == idx ? valid_31_0 : _GEN_34; // @[cache.scala 58:{66,66}]
  wire  _GEN_36 = 7'h20 == idx ? valid_32_0 : _GEN_35; // @[cache.scala 58:{66,66}]
  wire  _GEN_37 = 7'h21 == idx ? valid_33_0 : _GEN_36; // @[cache.scala 58:{66,66}]
  wire  _GEN_38 = 7'h22 == idx ? valid_34_0 : _GEN_37; // @[cache.scala 58:{66,66}]
  wire  _GEN_39 = 7'h23 == idx ? valid_35_0 : _GEN_38; // @[cache.scala 58:{66,66}]
  wire  _GEN_40 = 7'h24 == idx ? valid_36_0 : _GEN_39; // @[cache.scala 58:{66,66}]
  wire  _GEN_41 = 7'h25 == idx ? valid_37_0 : _GEN_40; // @[cache.scala 58:{66,66}]
  wire  _GEN_42 = 7'h26 == idx ? valid_38_0 : _GEN_41; // @[cache.scala 58:{66,66}]
  wire  _GEN_43 = 7'h27 == idx ? valid_39_0 : _GEN_42; // @[cache.scala 58:{66,66}]
  wire  _GEN_44 = 7'h28 == idx ? valid_40_0 : _GEN_43; // @[cache.scala 58:{66,66}]
  wire  _GEN_45 = 7'h29 == idx ? valid_41_0 : _GEN_44; // @[cache.scala 58:{66,66}]
  wire  _GEN_46 = 7'h2a == idx ? valid_42_0 : _GEN_45; // @[cache.scala 58:{66,66}]
  wire  _GEN_47 = 7'h2b == idx ? valid_43_0 : _GEN_46; // @[cache.scala 58:{66,66}]
  wire  _GEN_48 = 7'h2c == idx ? valid_44_0 : _GEN_47; // @[cache.scala 58:{66,66}]
  wire  _GEN_49 = 7'h2d == idx ? valid_45_0 : _GEN_48; // @[cache.scala 58:{66,66}]
  wire  _GEN_50 = 7'h2e == idx ? valid_46_0 : _GEN_49; // @[cache.scala 58:{66,66}]
  wire  _GEN_51 = 7'h2f == idx ? valid_47_0 : _GEN_50; // @[cache.scala 58:{66,66}]
  wire  _GEN_52 = 7'h30 == idx ? valid_48_0 : _GEN_51; // @[cache.scala 58:{66,66}]
  wire  _GEN_53 = 7'h31 == idx ? valid_49_0 : _GEN_52; // @[cache.scala 58:{66,66}]
  wire  _GEN_54 = 7'h32 == idx ? valid_50_0 : _GEN_53; // @[cache.scala 58:{66,66}]
  wire  _GEN_55 = 7'h33 == idx ? valid_51_0 : _GEN_54; // @[cache.scala 58:{66,66}]
  wire  _GEN_56 = 7'h34 == idx ? valid_52_0 : _GEN_55; // @[cache.scala 58:{66,66}]
  wire  _GEN_57 = 7'h35 == idx ? valid_53_0 : _GEN_56; // @[cache.scala 58:{66,66}]
  wire  _GEN_58 = 7'h36 == idx ? valid_54_0 : _GEN_57; // @[cache.scala 58:{66,66}]
  wire  _GEN_59 = 7'h37 == idx ? valid_55_0 : _GEN_58; // @[cache.scala 58:{66,66}]
  wire  _GEN_60 = 7'h38 == idx ? valid_56_0 : _GEN_59; // @[cache.scala 58:{66,66}]
  wire  _GEN_61 = 7'h39 == idx ? valid_57_0 : _GEN_60; // @[cache.scala 58:{66,66}]
  wire  _GEN_62 = 7'h3a == idx ? valid_58_0 : _GEN_61; // @[cache.scala 58:{66,66}]
  wire  _GEN_63 = 7'h3b == idx ? valid_59_0 : _GEN_62; // @[cache.scala 58:{66,66}]
  wire  _GEN_64 = 7'h3c == idx ? valid_60_0 : _GEN_63; // @[cache.scala 58:{66,66}]
  wire  _GEN_65 = 7'h3d == idx ? valid_61_0 : _GEN_64; // @[cache.scala 58:{66,66}]
  wire  _GEN_66 = 7'h3e == idx ? valid_62_0 : _GEN_65; // @[cache.scala 58:{66,66}]
  wire  _GEN_67 = 7'h3f == idx ? valid_63_0 : _GEN_66; // @[cache.scala 58:{66,66}]
  wire  _GEN_68 = 7'h40 == idx ? valid_64_0 : _GEN_67; // @[cache.scala 58:{66,66}]
  wire  _GEN_69 = 7'h41 == idx ? valid_65_0 : _GEN_68; // @[cache.scala 58:{66,66}]
  wire  _GEN_70 = 7'h42 == idx ? valid_66_0 : _GEN_69; // @[cache.scala 58:{66,66}]
  wire  _GEN_71 = 7'h43 == idx ? valid_67_0 : _GEN_70; // @[cache.scala 58:{66,66}]
  wire  _GEN_72 = 7'h44 == idx ? valid_68_0 : _GEN_71; // @[cache.scala 58:{66,66}]
  wire  _GEN_73 = 7'h45 == idx ? valid_69_0 : _GEN_72; // @[cache.scala 58:{66,66}]
  wire  _GEN_74 = 7'h46 == idx ? valid_70_0 : _GEN_73; // @[cache.scala 58:{66,66}]
  wire  _GEN_75 = 7'h47 == idx ? valid_71_0 : _GEN_74; // @[cache.scala 58:{66,66}]
  wire  _GEN_76 = 7'h48 == idx ? valid_72_0 : _GEN_75; // @[cache.scala 58:{66,66}]
  wire  _GEN_77 = 7'h49 == idx ? valid_73_0 : _GEN_76; // @[cache.scala 58:{66,66}]
  wire  _GEN_78 = 7'h4a == idx ? valid_74_0 : _GEN_77; // @[cache.scala 58:{66,66}]
  wire  _GEN_79 = 7'h4b == idx ? valid_75_0 : _GEN_78; // @[cache.scala 58:{66,66}]
  wire  _GEN_80 = 7'h4c == idx ? valid_76_0 : _GEN_79; // @[cache.scala 58:{66,66}]
  wire  _GEN_81 = 7'h4d == idx ? valid_77_0 : _GEN_80; // @[cache.scala 58:{66,66}]
  wire  _GEN_82 = 7'h4e == idx ? valid_78_0 : _GEN_81; // @[cache.scala 58:{66,66}]
  wire  _GEN_83 = 7'h4f == idx ? valid_79_0 : _GEN_82; // @[cache.scala 58:{66,66}]
  wire  _GEN_84 = 7'h50 == idx ? valid_80_0 : _GEN_83; // @[cache.scala 58:{66,66}]
  wire  _GEN_85 = 7'h51 == idx ? valid_81_0 : _GEN_84; // @[cache.scala 58:{66,66}]
  wire  _GEN_86 = 7'h52 == idx ? valid_82_0 : _GEN_85; // @[cache.scala 58:{66,66}]
  wire  _GEN_87 = 7'h53 == idx ? valid_83_0 : _GEN_86; // @[cache.scala 58:{66,66}]
  wire  _GEN_88 = 7'h54 == idx ? valid_84_0 : _GEN_87; // @[cache.scala 58:{66,66}]
  wire  _GEN_89 = 7'h55 == idx ? valid_85_0 : _GEN_88; // @[cache.scala 58:{66,66}]
  wire  _GEN_90 = 7'h56 == idx ? valid_86_0 : _GEN_89; // @[cache.scala 58:{66,66}]
  wire  _GEN_91 = 7'h57 == idx ? valid_87_0 : _GEN_90; // @[cache.scala 58:{66,66}]
  wire  _GEN_92 = 7'h58 == idx ? valid_88_0 : _GEN_91; // @[cache.scala 58:{66,66}]
  wire  _GEN_93 = 7'h59 == idx ? valid_89_0 : _GEN_92; // @[cache.scala 58:{66,66}]
  wire  _GEN_94 = 7'h5a == idx ? valid_90_0 : _GEN_93; // @[cache.scala 58:{66,66}]
  wire  _GEN_95 = 7'h5b == idx ? valid_91_0 : _GEN_94; // @[cache.scala 58:{66,66}]
  wire  _GEN_96 = 7'h5c == idx ? valid_92_0 : _GEN_95; // @[cache.scala 58:{66,66}]
  wire  _GEN_97 = 7'h5d == idx ? valid_93_0 : _GEN_96; // @[cache.scala 58:{66,66}]
  wire  _GEN_98 = 7'h5e == idx ? valid_94_0 : _GEN_97; // @[cache.scala 58:{66,66}]
  wire  _GEN_99 = 7'h5f == idx ? valid_95_0 : _GEN_98; // @[cache.scala 58:{66,66}]
  wire  _GEN_100 = 7'h60 == idx ? valid_96_0 : _GEN_99; // @[cache.scala 58:{66,66}]
  wire  _GEN_101 = 7'h61 == idx ? valid_97_0 : _GEN_100; // @[cache.scala 58:{66,66}]
  wire  _GEN_102 = 7'h62 == idx ? valid_98_0 : _GEN_101; // @[cache.scala 58:{66,66}]
  wire  _GEN_103 = 7'h63 == idx ? valid_99_0 : _GEN_102; // @[cache.scala 58:{66,66}]
  wire  _GEN_104 = 7'h64 == idx ? valid_100_0 : _GEN_103; // @[cache.scala 58:{66,66}]
  wire  _GEN_105 = 7'h65 == idx ? valid_101_0 : _GEN_104; // @[cache.scala 58:{66,66}]
  wire  _GEN_106 = 7'h66 == idx ? valid_102_0 : _GEN_105; // @[cache.scala 58:{66,66}]
  wire  _GEN_107 = 7'h67 == idx ? valid_103_0 : _GEN_106; // @[cache.scala 58:{66,66}]
  wire  _GEN_108 = 7'h68 == idx ? valid_104_0 : _GEN_107; // @[cache.scala 58:{66,66}]
  wire  _GEN_109 = 7'h69 == idx ? valid_105_0 : _GEN_108; // @[cache.scala 58:{66,66}]
  wire  _GEN_110 = 7'h6a == idx ? valid_106_0 : _GEN_109; // @[cache.scala 58:{66,66}]
  wire  _GEN_111 = 7'h6b == idx ? valid_107_0 : _GEN_110; // @[cache.scala 58:{66,66}]
  wire  _GEN_112 = 7'h6c == idx ? valid_108_0 : _GEN_111; // @[cache.scala 58:{66,66}]
  wire  _GEN_113 = 7'h6d == idx ? valid_109_0 : _GEN_112; // @[cache.scala 58:{66,66}]
  wire  _GEN_114 = 7'h6e == idx ? valid_110_0 : _GEN_113; // @[cache.scala 58:{66,66}]
  wire  _GEN_115 = 7'h6f == idx ? valid_111_0 : _GEN_114; // @[cache.scala 58:{66,66}]
  wire  _GEN_116 = 7'h70 == idx ? valid_112_0 : _GEN_115; // @[cache.scala 58:{66,66}]
  wire  _GEN_117 = 7'h71 == idx ? valid_113_0 : _GEN_116; // @[cache.scala 58:{66,66}]
  wire  _GEN_118 = 7'h72 == idx ? valid_114_0 : _GEN_117; // @[cache.scala 58:{66,66}]
  wire  _GEN_119 = 7'h73 == idx ? valid_115_0 : _GEN_118; // @[cache.scala 58:{66,66}]
  wire  _GEN_120 = 7'h74 == idx ? valid_116_0 : _GEN_119; // @[cache.scala 58:{66,66}]
  wire  _GEN_121 = 7'h75 == idx ? valid_117_0 : _GEN_120; // @[cache.scala 58:{66,66}]
  wire  _GEN_122 = 7'h76 == idx ? valid_118_0 : _GEN_121; // @[cache.scala 58:{66,66}]
  wire  _GEN_123 = 7'h77 == idx ? valid_119_0 : _GEN_122; // @[cache.scala 58:{66,66}]
  wire  _GEN_124 = 7'h78 == idx ? valid_120_0 : _GEN_123; // @[cache.scala 58:{66,66}]
  wire  _GEN_125 = 7'h79 == idx ? valid_121_0 : _GEN_124; // @[cache.scala 58:{66,66}]
  wire  _GEN_126 = 7'h7a == idx ? valid_122_0 : _GEN_125; // @[cache.scala 58:{66,66}]
  wire  _GEN_127 = 7'h7b == idx ? valid_123_0 : _GEN_126; // @[cache.scala 58:{66,66}]
  wire  _GEN_128 = 7'h7c == idx ? valid_124_0 : _GEN_127; // @[cache.scala 58:{66,66}]
  wire  _GEN_129 = 7'h7d == idx ? valid_125_0 : _GEN_128; // @[cache.scala 58:{66,66}]
  wire  _GEN_130 = 7'h7e == idx ? valid_126_0 : _GEN_129; // @[cache.scala 58:{66,66}]
  wire  _GEN_131 = 7'h7f == idx ? valid_127_0 : _GEN_130; // @[cache.scala 58:{66,66}]
  wire  _GEN_133 = 7'h1 == idx ? valid_1_1 : valid_0_1; // @[cache.scala 59:{66,66}]
  wire  _GEN_134 = 7'h2 == idx ? valid_2_1 : _GEN_133; // @[cache.scala 59:{66,66}]
  wire  _GEN_135 = 7'h3 == idx ? valid_3_1 : _GEN_134; // @[cache.scala 59:{66,66}]
  wire  _GEN_136 = 7'h4 == idx ? valid_4_1 : _GEN_135; // @[cache.scala 59:{66,66}]
  wire  _GEN_137 = 7'h5 == idx ? valid_5_1 : _GEN_136; // @[cache.scala 59:{66,66}]
  wire  _GEN_138 = 7'h6 == idx ? valid_6_1 : _GEN_137; // @[cache.scala 59:{66,66}]
  wire  _GEN_139 = 7'h7 == idx ? valid_7_1 : _GEN_138; // @[cache.scala 59:{66,66}]
  wire  _GEN_140 = 7'h8 == idx ? valid_8_1 : _GEN_139; // @[cache.scala 59:{66,66}]
  wire  _GEN_141 = 7'h9 == idx ? valid_9_1 : _GEN_140; // @[cache.scala 59:{66,66}]
  wire  _GEN_142 = 7'ha == idx ? valid_10_1 : _GEN_141; // @[cache.scala 59:{66,66}]
  wire  _GEN_143 = 7'hb == idx ? valid_11_1 : _GEN_142; // @[cache.scala 59:{66,66}]
  wire  _GEN_144 = 7'hc == idx ? valid_12_1 : _GEN_143; // @[cache.scala 59:{66,66}]
  wire  _GEN_145 = 7'hd == idx ? valid_13_1 : _GEN_144; // @[cache.scala 59:{66,66}]
  wire  _GEN_146 = 7'he == idx ? valid_14_1 : _GEN_145; // @[cache.scala 59:{66,66}]
  wire  _GEN_147 = 7'hf == idx ? valid_15_1 : _GEN_146; // @[cache.scala 59:{66,66}]
  wire  _GEN_148 = 7'h10 == idx ? valid_16_1 : _GEN_147; // @[cache.scala 59:{66,66}]
  wire  _GEN_149 = 7'h11 == idx ? valid_17_1 : _GEN_148; // @[cache.scala 59:{66,66}]
  wire  _GEN_150 = 7'h12 == idx ? valid_18_1 : _GEN_149; // @[cache.scala 59:{66,66}]
  wire  _GEN_151 = 7'h13 == idx ? valid_19_1 : _GEN_150; // @[cache.scala 59:{66,66}]
  wire  _GEN_152 = 7'h14 == idx ? valid_20_1 : _GEN_151; // @[cache.scala 59:{66,66}]
  wire  _GEN_153 = 7'h15 == idx ? valid_21_1 : _GEN_152; // @[cache.scala 59:{66,66}]
  wire  _GEN_154 = 7'h16 == idx ? valid_22_1 : _GEN_153; // @[cache.scala 59:{66,66}]
  wire  _GEN_155 = 7'h17 == idx ? valid_23_1 : _GEN_154; // @[cache.scala 59:{66,66}]
  wire  _GEN_156 = 7'h18 == idx ? valid_24_1 : _GEN_155; // @[cache.scala 59:{66,66}]
  wire  _GEN_157 = 7'h19 == idx ? valid_25_1 : _GEN_156; // @[cache.scala 59:{66,66}]
  wire  _GEN_158 = 7'h1a == idx ? valid_26_1 : _GEN_157; // @[cache.scala 59:{66,66}]
  wire  _GEN_159 = 7'h1b == idx ? valid_27_1 : _GEN_158; // @[cache.scala 59:{66,66}]
  wire  _GEN_160 = 7'h1c == idx ? valid_28_1 : _GEN_159; // @[cache.scala 59:{66,66}]
  wire  _GEN_161 = 7'h1d == idx ? valid_29_1 : _GEN_160; // @[cache.scala 59:{66,66}]
  wire  _GEN_162 = 7'h1e == idx ? valid_30_1 : _GEN_161; // @[cache.scala 59:{66,66}]
  wire  _GEN_163 = 7'h1f == idx ? valid_31_1 : _GEN_162; // @[cache.scala 59:{66,66}]
  wire  _GEN_164 = 7'h20 == idx ? valid_32_1 : _GEN_163; // @[cache.scala 59:{66,66}]
  wire  _GEN_165 = 7'h21 == idx ? valid_33_1 : _GEN_164; // @[cache.scala 59:{66,66}]
  wire  _GEN_166 = 7'h22 == idx ? valid_34_1 : _GEN_165; // @[cache.scala 59:{66,66}]
  wire  _GEN_167 = 7'h23 == idx ? valid_35_1 : _GEN_166; // @[cache.scala 59:{66,66}]
  wire  _GEN_168 = 7'h24 == idx ? valid_36_1 : _GEN_167; // @[cache.scala 59:{66,66}]
  wire  _GEN_169 = 7'h25 == idx ? valid_37_1 : _GEN_168; // @[cache.scala 59:{66,66}]
  wire  _GEN_170 = 7'h26 == idx ? valid_38_1 : _GEN_169; // @[cache.scala 59:{66,66}]
  wire  _GEN_171 = 7'h27 == idx ? valid_39_1 : _GEN_170; // @[cache.scala 59:{66,66}]
  wire  _GEN_172 = 7'h28 == idx ? valid_40_1 : _GEN_171; // @[cache.scala 59:{66,66}]
  wire  _GEN_173 = 7'h29 == idx ? valid_41_1 : _GEN_172; // @[cache.scala 59:{66,66}]
  wire  _GEN_174 = 7'h2a == idx ? valid_42_1 : _GEN_173; // @[cache.scala 59:{66,66}]
  wire  _GEN_175 = 7'h2b == idx ? valid_43_1 : _GEN_174; // @[cache.scala 59:{66,66}]
  wire  _GEN_176 = 7'h2c == idx ? valid_44_1 : _GEN_175; // @[cache.scala 59:{66,66}]
  wire  _GEN_177 = 7'h2d == idx ? valid_45_1 : _GEN_176; // @[cache.scala 59:{66,66}]
  wire  _GEN_178 = 7'h2e == idx ? valid_46_1 : _GEN_177; // @[cache.scala 59:{66,66}]
  wire  _GEN_179 = 7'h2f == idx ? valid_47_1 : _GEN_178; // @[cache.scala 59:{66,66}]
  wire  _GEN_180 = 7'h30 == idx ? valid_48_1 : _GEN_179; // @[cache.scala 59:{66,66}]
  wire  _GEN_181 = 7'h31 == idx ? valid_49_1 : _GEN_180; // @[cache.scala 59:{66,66}]
  wire  _GEN_182 = 7'h32 == idx ? valid_50_1 : _GEN_181; // @[cache.scala 59:{66,66}]
  wire  _GEN_183 = 7'h33 == idx ? valid_51_1 : _GEN_182; // @[cache.scala 59:{66,66}]
  wire  _GEN_184 = 7'h34 == idx ? valid_52_1 : _GEN_183; // @[cache.scala 59:{66,66}]
  wire  _GEN_185 = 7'h35 == idx ? valid_53_1 : _GEN_184; // @[cache.scala 59:{66,66}]
  wire  _GEN_186 = 7'h36 == idx ? valid_54_1 : _GEN_185; // @[cache.scala 59:{66,66}]
  wire  _GEN_187 = 7'h37 == idx ? valid_55_1 : _GEN_186; // @[cache.scala 59:{66,66}]
  wire  _GEN_188 = 7'h38 == idx ? valid_56_1 : _GEN_187; // @[cache.scala 59:{66,66}]
  wire  _GEN_189 = 7'h39 == idx ? valid_57_1 : _GEN_188; // @[cache.scala 59:{66,66}]
  wire  _GEN_190 = 7'h3a == idx ? valid_58_1 : _GEN_189; // @[cache.scala 59:{66,66}]
  wire  _GEN_191 = 7'h3b == idx ? valid_59_1 : _GEN_190; // @[cache.scala 59:{66,66}]
  wire  _GEN_192 = 7'h3c == idx ? valid_60_1 : _GEN_191; // @[cache.scala 59:{66,66}]
  wire  _GEN_193 = 7'h3d == idx ? valid_61_1 : _GEN_192; // @[cache.scala 59:{66,66}]
  wire  _GEN_194 = 7'h3e == idx ? valid_62_1 : _GEN_193; // @[cache.scala 59:{66,66}]
  wire  _GEN_195 = 7'h3f == idx ? valid_63_1 : _GEN_194; // @[cache.scala 59:{66,66}]
  wire  _GEN_196 = 7'h40 == idx ? valid_64_1 : _GEN_195; // @[cache.scala 59:{66,66}]
  wire  _GEN_197 = 7'h41 == idx ? valid_65_1 : _GEN_196; // @[cache.scala 59:{66,66}]
  wire  _GEN_198 = 7'h42 == idx ? valid_66_1 : _GEN_197; // @[cache.scala 59:{66,66}]
  wire  _GEN_199 = 7'h43 == idx ? valid_67_1 : _GEN_198; // @[cache.scala 59:{66,66}]
  wire  _GEN_200 = 7'h44 == idx ? valid_68_1 : _GEN_199; // @[cache.scala 59:{66,66}]
  wire  _GEN_201 = 7'h45 == idx ? valid_69_1 : _GEN_200; // @[cache.scala 59:{66,66}]
  wire  _GEN_202 = 7'h46 == idx ? valid_70_1 : _GEN_201; // @[cache.scala 59:{66,66}]
  wire  _GEN_203 = 7'h47 == idx ? valid_71_1 : _GEN_202; // @[cache.scala 59:{66,66}]
  wire  _GEN_204 = 7'h48 == idx ? valid_72_1 : _GEN_203; // @[cache.scala 59:{66,66}]
  wire  _GEN_205 = 7'h49 == idx ? valid_73_1 : _GEN_204; // @[cache.scala 59:{66,66}]
  wire  _GEN_206 = 7'h4a == idx ? valid_74_1 : _GEN_205; // @[cache.scala 59:{66,66}]
  wire  _GEN_207 = 7'h4b == idx ? valid_75_1 : _GEN_206; // @[cache.scala 59:{66,66}]
  wire  _GEN_208 = 7'h4c == idx ? valid_76_1 : _GEN_207; // @[cache.scala 59:{66,66}]
  wire  _GEN_209 = 7'h4d == idx ? valid_77_1 : _GEN_208; // @[cache.scala 59:{66,66}]
  wire  _GEN_210 = 7'h4e == idx ? valid_78_1 : _GEN_209; // @[cache.scala 59:{66,66}]
  wire  _GEN_211 = 7'h4f == idx ? valid_79_1 : _GEN_210; // @[cache.scala 59:{66,66}]
  wire  _GEN_212 = 7'h50 == idx ? valid_80_1 : _GEN_211; // @[cache.scala 59:{66,66}]
  wire  _GEN_213 = 7'h51 == idx ? valid_81_1 : _GEN_212; // @[cache.scala 59:{66,66}]
  wire  _GEN_214 = 7'h52 == idx ? valid_82_1 : _GEN_213; // @[cache.scala 59:{66,66}]
  wire  _GEN_215 = 7'h53 == idx ? valid_83_1 : _GEN_214; // @[cache.scala 59:{66,66}]
  wire  _GEN_216 = 7'h54 == idx ? valid_84_1 : _GEN_215; // @[cache.scala 59:{66,66}]
  wire  _GEN_217 = 7'h55 == idx ? valid_85_1 : _GEN_216; // @[cache.scala 59:{66,66}]
  wire  _GEN_218 = 7'h56 == idx ? valid_86_1 : _GEN_217; // @[cache.scala 59:{66,66}]
  wire  _GEN_219 = 7'h57 == idx ? valid_87_1 : _GEN_218; // @[cache.scala 59:{66,66}]
  wire  _GEN_220 = 7'h58 == idx ? valid_88_1 : _GEN_219; // @[cache.scala 59:{66,66}]
  wire  _GEN_221 = 7'h59 == idx ? valid_89_1 : _GEN_220; // @[cache.scala 59:{66,66}]
  wire  _GEN_222 = 7'h5a == idx ? valid_90_1 : _GEN_221; // @[cache.scala 59:{66,66}]
  wire  _GEN_223 = 7'h5b == idx ? valid_91_1 : _GEN_222; // @[cache.scala 59:{66,66}]
  wire  _GEN_224 = 7'h5c == idx ? valid_92_1 : _GEN_223; // @[cache.scala 59:{66,66}]
  wire  _GEN_225 = 7'h5d == idx ? valid_93_1 : _GEN_224; // @[cache.scala 59:{66,66}]
  wire  _GEN_226 = 7'h5e == idx ? valid_94_1 : _GEN_225; // @[cache.scala 59:{66,66}]
  wire  _GEN_227 = 7'h5f == idx ? valid_95_1 : _GEN_226; // @[cache.scala 59:{66,66}]
  wire  _GEN_228 = 7'h60 == idx ? valid_96_1 : _GEN_227; // @[cache.scala 59:{66,66}]
  wire  _GEN_229 = 7'h61 == idx ? valid_97_1 : _GEN_228; // @[cache.scala 59:{66,66}]
  wire  _GEN_230 = 7'h62 == idx ? valid_98_1 : _GEN_229; // @[cache.scala 59:{66,66}]
  wire  _GEN_231 = 7'h63 == idx ? valid_99_1 : _GEN_230; // @[cache.scala 59:{66,66}]
  wire  _GEN_232 = 7'h64 == idx ? valid_100_1 : _GEN_231; // @[cache.scala 59:{66,66}]
  wire  _GEN_233 = 7'h65 == idx ? valid_101_1 : _GEN_232; // @[cache.scala 59:{66,66}]
  wire  _GEN_234 = 7'h66 == idx ? valid_102_1 : _GEN_233; // @[cache.scala 59:{66,66}]
  wire  _GEN_235 = 7'h67 == idx ? valid_103_1 : _GEN_234; // @[cache.scala 59:{66,66}]
  wire  _GEN_236 = 7'h68 == idx ? valid_104_1 : _GEN_235; // @[cache.scala 59:{66,66}]
  wire  _GEN_237 = 7'h69 == idx ? valid_105_1 : _GEN_236; // @[cache.scala 59:{66,66}]
  wire  _GEN_238 = 7'h6a == idx ? valid_106_1 : _GEN_237; // @[cache.scala 59:{66,66}]
  wire  _GEN_239 = 7'h6b == idx ? valid_107_1 : _GEN_238; // @[cache.scala 59:{66,66}]
  wire  _GEN_240 = 7'h6c == idx ? valid_108_1 : _GEN_239; // @[cache.scala 59:{66,66}]
  wire  _GEN_241 = 7'h6d == idx ? valid_109_1 : _GEN_240; // @[cache.scala 59:{66,66}]
  wire  _GEN_242 = 7'h6e == idx ? valid_110_1 : _GEN_241; // @[cache.scala 59:{66,66}]
  wire  _GEN_243 = 7'h6f == idx ? valid_111_1 : _GEN_242; // @[cache.scala 59:{66,66}]
  wire  _GEN_244 = 7'h70 == idx ? valid_112_1 : _GEN_243; // @[cache.scala 59:{66,66}]
  wire  _GEN_245 = 7'h71 == idx ? valid_113_1 : _GEN_244; // @[cache.scala 59:{66,66}]
  wire  _GEN_246 = 7'h72 == idx ? valid_114_1 : _GEN_245; // @[cache.scala 59:{66,66}]
  wire  _GEN_247 = 7'h73 == idx ? valid_115_1 : _GEN_246; // @[cache.scala 59:{66,66}]
  wire  _GEN_248 = 7'h74 == idx ? valid_116_1 : _GEN_247; // @[cache.scala 59:{66,66}]
  wire  _GEN_249 = 7'h75 == idx ? valid_117_1 : _GEN_248; // @[cache.scala 59:{66,66}]
  wire  _GEN_250 = 7'h76 == idx ? valid_118_1 : _GEN_249; // @[cache.scala 59:{66,66}]
  wire  _GEN_251 = 7'h77 == idx ? valid_119_1 : _GEN_250; // @[cache.scala 59:{66,66}]
  wire  _GEN_252 = 7'h78 == idx ? valid_120_1 : _GEN_251; // @[cache.scala 59:{66,66}]
  wire  _GEN_253 = 7'h79 == idx ? valid_121_1 : _GEN_252; // @[cache.scala 59:{66,66}]
  wire  _GEN_254 = 7'h7a == idx ? valid_122_1 : _GEN_253; // @[cache.scala 59:{66,66}]
  wire  _GEN_255 = 7'h7b == idx ? valid_123_1 : _GEN_254; // @[cache.scala 59:{66,66}]
  wire  _GEN_256 = 7'h7c == idx ? valid_124_1 : _GEN_255; // @[cache.scala 59:{66,66}]
  wire  _GEN_257 = 7'h7d == idx ? valid_125_1 : _GEN_256; // @[cache.scala 59:{66,66}]
  wire  _GEN_258 = 7'h7e == idx ? valid_126_1 : _GEN_257; // @[cache.scala 59:{66,66}]
  wire  _GEN_259 = 7'h7f == idx ? valid_127_1 : _GEN_258; // @[cache.scala 59:{66,66}]
  wire [7:0] _hit_way_T_8 = tag_read[41:21] == tag & _GEN_259 ? 8'h1 : 8'hff; // @[cache.scala 59:18]
  wire [7:0] hit_way = tag_read[20:0] == tag & _GEN_131 ? 8'h0 : _hit_way_T_8; // @[cache.scala 58:18]
  wire [7:0] idxh = _idxh_T | hit_way; // @[cache.scala 44:25]
  wire [7:0] idxw = _idxh_T | way2; // @[cache.scala 45:25]
  reg  rmode; // @[cache.scala 51:22]
  reg  wmode; // @[cache.scala 52:22]
  wire  _rmode_T = state == 4'h0; // @[cache.scala 53:23]
  wire  _rmode_T_1 = io_in_ar_ready & io_in_ar_valid; // @[Decoupled.scala 52:35]
  wire  _rmode_T_2 = state == 4'h0 & _rmode_T_1; // @[cache.scala 53:35]
  wire  _rmode_T_4 = state == 4'h0 ? 1'h0 : rmode; // @[cache.scala 53:58]
  wire  _wmode_T_1 = io_in_aw_ready & io_in_aw_valid; // @[Decoupled.scala 52:35]
  wire  _wmode_T_2 = _rmode_T & _wmode_T_1; // @[cache.scala 54:35]
  wire  _wmode_T_4 = _rmode_T ? 1'h0 : wmode; // @[cache.scala 54:58]
  wire  _tag_way_T = way2 == 8'h0; // @[cache.scala 65:23]
  wire [20:0] tag_way = way2 == 8'h0 ? tag_read[20:0] : tag_read[41:21]; // @[cache.scala 65:17]
  wire [3:0] _state_T_3 = _wmode_T_1 | _rmode_T_1 ? 4'h1 : 4'h0; // @[cache.scala 68:20]
  wire [3:0] _state_T_5 = hit_way == 8'hff ? 4'h4 : 4'h3; // @[cache.scala 70:19]
  wire  _GEN_2057 = 7'h0 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_261 = 7'h0 == idx & way2[0] ? dirty_0_1 : dirty_0_0; // @[cache.scala 72:{64,64}]
  wire  _GEN_2058 = 7'h1 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_2059 = ~way2[0]; // @[cache.scala 72:{64,64}]
  wire  _GEN_262 = 7'h1 == idx & ~way2[0] ? dirty_1_0 : _GEN_261; // @[cache.scala 72:{64,64}]
  wire  _GEN_263 = 7'h1 == idx & way2[0] ? dirty_1_1 : _GEN_262; // @[cache.scala 72:{64,64}]
  wire  _GEN_2061 = 7'h2 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_264 = 7'h2 == idx & ~way2[0] ? dirty_2_0 : _GEN_263; // @[cache.scala 72:{64,64}]
  wire  _GEN_265 = 7'h2 == idx & way2[0] ? dirty_2_1 : _GEN_264; // @[cache.scala 72:{64,64}]
  wire  _GEN_2064 = 7'h3 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_266 = 7'h3 == idx & ~way2[0] ? dirty_3_0 : _GEN_265; // @[cache.scala 72:{64,64}]
  wire  _GEN_267 = 7'h3 == idx & way2[0] ? dirty_3_1 : _GEN_266; // @[cache.scala 72:{64,64}]
  wire  _GEN_2067 = 7'h4 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_268 = 7'h4 == idx & ~way2[0] ? dirty_4_0 : _GEN_267; // @[cache.scala 72:{64,64}]
  wire  _GEN_269 = 7'h4 == idx & way2[0] ? dirty_4_1 : _GEN_268; // @[cache.scala 72:{64,64}]
  wire  _GEN_2070 = 7'h5 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_270 = 7'h5 == idx & ~way2[0] ? dirty_5_0 : _GEN_269; // @[cache.scala 72:{64,64}]
  wire  _GEN_271 = 7'h5 == idx & way2[0] ? dirty_5_1 : _GEN_270; // @[cache.scala 72:{64,64}]
  wire  _GEN_2073 = 7'h6 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_272 = 7'h6 == idx & ~way2[0] ? dirty_6_0 : _GEN_271; // @[cache.scala 72:{64,64}]
  wire  _GEN_273 = 7'h6 == idx & way2[0] ? dirty_6_1 : _GEN_272; // @[cache.scala 72:{64,64}]
  wire  _GEN_2076 = 7'h7 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_274 = 7'h7 == idx & ~way2[0] ? dirty_7_0 : _GEN_273; // @[cache.scala 72:{64,64}]
  wire  _GEN_275 = 7'h7 == idx & way2[0] ? dirty_7_1 : _GEN_274; // @[cache.scala 72:{64,64}]
  wire  _GEN_2079 = 7'h8 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_276 = 7'h8 == idx & ~way2[0] ? dirty_8_0 : _GEN_275; // @[cache.scala 72:{64,64}]
  wire  _GEN_277 = 7'h8 == idx & way2[0] ? dirty_8_1 : _GEN_276; // @[cache.scala 72:{64,64}]
  wire  _GEN_2082 = 7'h9 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_278 = 7'h9 == idx & ~way2[0] ? dirty_9_0 : _GEN_277; // @[cache.scala 72:{64,64}]
  wire  _GEN_279 = 7'h9 == idx & way2[0] ? dirty_9_1 : _GEN_278; // @[cache.scala 72:{64,64}]
  wire  _GEN_2085 = 7'ha == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_280 = 7'ha == idx & ~way2[0] ? dirty_10_0 : _GEN_279; // @[cache.scala 72:{64,64}]
  wire  _GEN_281 = 7'ha == idx & way2[0] ? dirty_10_1 : _GEN_280; // @[cache.scala 72:{64,64}]
  wire  _GEN_2088 = 7'hb == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_282 = 7'hb == idx & ~way2[0] ? dirty_11_0 : _GEN_281; // @[cache.scala 72:{64,64}]
  wire  _GEN_283 = 7'hb == idx & way2[0] ? dirty_11_1 : _GEN_282; // @[cache.scala 72:{64,64}]
  wire  _GEN_2091 = 7'hc == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_284 = 7'hc == idx & ~way2[0] ? dirty_12_0 : _GEN_283; // @[cache.scala 72:{64,64}]
  wire  _GEN_285 = 7'hc == idx & way2[0] ? dirty_12_1 : _GEN_284; // @[cache.scala 72:{64,64}]
  wire  _GEN_2094 = 7'hd == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_286 = 7'hd == idx & ~way2[0] ? dirty_13_0 : _GEN_285; // @[cache.scala 72:{64,64}]
  wire  _GEN_287 = 7'hd == idx & way2[0] ? dirty_13_1 : _GEN_286; // @[cache.scala 72:{64,64}]
  wire  _GEN_2097 = 7'he == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_288 = 7'he == idx & ~way2[0] ? dirty_14_0 : _GEN_287; // @[cache.scala 72:{64,64}]
  wire  _GEN_289 = 7'he == idx & way2[0] ? dirty_14_1 : _GEN_288; // @[cache.scala 72:{64,64}]
  wire  _GEN_2100 = 7'hf == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_290 = 7'hf == idx & ~way2[0] ? dirty_15_0 : _GEN_289; // @[cache.scala 72:{64,64}]
  wire  _GEN_291 = 7'hf == idx & way2[0] ? dirty_15_1 : _GEN_290; // @[cache.scala 72:{64,64}]
  wire  _GEN_2103 = 7'h10 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_292 = 7'h10 == idx & ~way2[0] ? dirty_16_0 : _GEN_291; // @[cache.scala 72:{64,64}]
  wire  _GEN_293 = 7'h10 == idx & way2[0] ? dirty_16_1 : _GEN_292; // @[cache.scala 72:{64,64}]
  wire  _GEN_2106 = 7'h11 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_294 = 7'h11 == idx & ~way2[0] ? dirty_17_0 : _GEN_293; // @[cache.scala 72:{64,64}]
  wire  _GEN_295 = 7'h11 == idx & way2[0] ? dirty_17_1 : _GEN_294; // @[cache.scala 72:{64,64}]
  wire  _GEN_2109 = 7'h12 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_296 = 7'h12 == idx & ~way2[0] ? dirty_18_0 : _GEN_295; // @[cache.scala 72:{64,64}]
  wire  _GEN_297 = 7'h12 == idx & way2[0] ? dirty_18_1 : _GEN_296; // @[cache.scala 72:{64,64}]
  wire  _GEN_2112 = 7'h13 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_298 = 7'h13 == idx & ~way2[0] ? dirty_19_0 : _GEN_297; // @[cache.scala 72:{64,64}]
  wire  _GEN_299 = 7'h13 == idx & way2[0] ? dirty_19_1 : _GEN_298; // @[cache.scala 72:{64,64}]
  wire  _GEN_2115 = 7'h14 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_300 = 7'h14 == idx & ~way2[0] ? dirty_20_0 : _GEN_299; // @[cache.scala 72:{64,64}]
  wire  _GEN_301 = 7'h14 == idx & way2[0] ? dirty_20_1 : _GEN_300; // @[cache.scala 72:{64,64}]
  wire  _GEN_2118 = 7'h15 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_302 = 7'h15 == idx & ~way2[0] ? dirty_21_0 : _GEN_301; // @[cache.scala 72:{64,64}]
  wire  _GEN_303 = 7'h15 == idx & way2[0] ? dirty_21_1 : _GEN_302; // @[cache.scala 72:{64,64}]
  wire  _GEN_2121 = 7'h16 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_304 = 7'h16 == idx & ~way2[0] ? dirty_22_0 : _GEN_303; // @[cache.scala 72:{64,64}]
  wire  _GEN_305 = 7'h16 == idx & way2[0] ? dirty_22_1 : _GEN_304; // @[cache.scala 72:{64,64}]
  wire  _GEN_2124 = 7'h17 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_306 = 7'h17 == idx & ~way2[0] ? dirty_23_0 : _GEN_305; // @[cache.scala 72:{64,64}]
  wire  _GEN_307 = 7'h17 == idx & way2[0] ? dirty_23_1 : _GEN_306; // @[cache.scala 72:{64,64}]
  wire  _GEN_2127 = 7'h18 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_308 = 7'h18 == idx & ~way2[0] ? dirty_24_0 : _GEN_307; // @[cache.scala 72:{64,64}]
  wire  _GEN_309 = 7'h18 == idx & way2[0] ? dirty_24_1 : _GEN_308; // @[cache.scala 72:{64,64}]
  wire  _GEN_2130 = 7'h19 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_310 = 7'h19 == idx & ~way2[0] ? dirty_25_0 : _GEN_309; // @[cache.scala 72:{64,64}]
  wire  _GEN_311 = 7'h19 == idx & way2[0] ? dirty_25_1 : _GEN_310; // @[cache.scala 72:{64,64}]
  wire  _GEN_2133 = 7'h1a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_312 = 7'h1a == idx & ~way2[0] ? dirty_26_0 : _GEN_311; // @[cache.scala 72:{64,64}]
  wire  _GEN_313 = 7'h1a == idx & way2[0] ? dirty_26_1 : _GEN_312; // @[cache.scala 72:{64,64}]
  wire  _GEN_2136 = 7'h1b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_314 = 7'h1b == idx & ~way2[0] ? dirty_27_0 : _GEN_313; // @[cache.scala 72:{64,64}]
  wire  _GEN_315 = 7'h1b == idx & way2[0] ? dirty_27_1 : _GEN_314; // @[cache.scala 72:{64,64}]
  wire  _GEN_2139 = 7'h1c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_316 = 7'h1c == idx & ~way2[0] ? dirty_28_0 : _GEN_315; // @[cache.scala 72:{64,64}]
  wire  _GEN_317 = 7'h1c == idx & way2[0] ? dirty_28_1 : _GEN_316; // @[cache.scala 72:{64,64}]
  wire  _GEN_2142 = 7'h1d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_318 = 7'h1d == idx & ~way2[0] ? dirty_29_0 : _GEN_317; // @[cache.scala 72:{64,64}]
  wire  _GEN_319 = 7'h1d == idx & way2[0] ? dirty_29_1 : _GEN_318; // @[cache.scala 72:{64,64}]
  wire  _GEN_2145 = 7'h1e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_320 = 7'h1e == idx & ~way2[0] ? dirty_30_0 : _GEN_319; // @[cache.scala 72:{64,64}]
  wire  _GEN_321 = 7'h1e == idx & way2[0] ? dirty_30_1 : _GEN_320; // @[cache.scala 72:{64,64}]
  wire  _GEN_2148 = 7'h1f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_322 = 7'h1f == idx & ~way2[0] ? dirty_31_0 : _GEN_321; // @[cache.scala 72:{64,64}]
  wire  _GEN_323 = 7'h1f == idx & way2[0] ? dirty_31_1 : _GEN_322; // @[cache.scala 72:{64,64}]
  wire  _GEN_2151 = 7'h20 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_324 = 7'h20 == idx & ~way2[0] ? dirty_32_0 : _GEN_323; // @[cache.scala 72:{64,64}]
  wire  _GEN_325 = 7'h20 == idx & way2[0] ? dirty_32_1 : _GEN_324; // @[cache.scala 72:{64,64}]
  wire  _GEN_2154 = 7'h21 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_326 = 7'h21 == idx & ~way2[0] ? dirty_33_0 : _GEN_325; // @[cache.scala 72:{64,64}]
  wire  _GEN_327 = 7'h21 == idx & way2[0] ? dirty_33_1 : _GEN_326; // @[cache.scala 72:{64,64}]
  wire  _GEN_2157 = 7'h22 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_328 = 7'h22 == idx & ~way2[0] ? dirty_34_0 : _GEN_327; // @[cache.scala 72:{64,64}]
  wire  _GEN_329 = 7'h22 == idx & way2[0] ? dirty_34_1 : _GEN_328; // @[cache.scala 72:{64,64}]
  wire  _GEN_2160 = 7'h23 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_330 = 7'h23 == idx & ~way2[0] ? dirty_35_0 : _GEN_329; // @[cache.scala 72:{64,64}]
  wire  _GEN_331 = 7'h23 == idx & way2[0] ? dirty_35_1 : _GEN_330; // @[cache.scala 72:{64,64}]
  wire  _GEN_2163 = 7'h24 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_332 = 7'h24 == idx & ~way2[0] ? dirty_36_0 : _GEN_331; // @[cache.scala 72:{64,64}]
  wire  _GEN_333 = 7'h24 == idx & way2[0] ? dirty_36_1 : _GEN_332; // @[cache.scala 72:{64,64}]
  wire  _GEN_2166 = 7'h25 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_334 = 7'h25 == idx & ~way2[0] ? dirty_37_0 : _GEN_333; // @[cache.scala 72:{64,64}]
  wire  _GEN_335 = 7'h25 == idx & way2[0] ? dirty_37_1 : _GEN_334; // @[cache.scala 72:{64,64}]
  wire  _GEN_2169 = 7'h26 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_336 = 7'h26 == idx & ~way2[0] ? dirty_38_0 : _GEN_335; // @[cache.scala 72:{64,64}]
  wire  _GEN_337 = 7'h26 == idx & way2[0] ? dirty_38_1 : _GEN_336; // @[cache.scala 72:{64,64}]
  wire  _GEN_2172 = 7'h27 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_338 = 7'h27 == idx & ~way2[0] ? dirty_39_0 : _GEN_337; // @[cache.scala 72:{64,64}]
  wire  _GEN_339 = 7'h27 == idx & way2[0] ? dirty_39_1 : _GEN_338; // @[cache.scala 72:{64,64}]
  wire  _GEN_2175 = 7'h28 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_340 = 7'h28 == idx & ~way2[0] ? dirty_40_0 : _GEN_339; // @[cache.scala 72:{64,64}]
  wire  _GEN_341 = 7'h28 == idx & way2[0] ? dirty_40_1 : _GEN_340; // @[cache.scala 72:{64,64}]
  wire  _GEN_2178 = 7'h29 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_342 = 7'h29 == idx & ~way2[0] ? dirty_41_0 : _GEN_341; // @[cache.scala 72:{64,64}]
  wire  _GEN_343 = 7'h29 == idx & way2[0] ? dirty_41_1 : _GEN_342; // @[cache.scala 72:{64,64}]
  wire  _GEN_2181 = 7'h2a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_344 = 7'h2a == idx & ~way2[0] ? dirty_42_0 : _GEN_343; // @[cache.scala 72:{64,64}]
  wire  _GEN_345 = 7'h2a == idx & way2[0] ? dirty_42_1 : _GEN_344; // @[cache.scala 72:{64,64}]
  wire  _GEN_2184 = 7'h2b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_346 = 7'h2b == idx & ~way2[0] ? dirty_43_0 : _GEN_345; // @[cache.scala 72:{64,64}]
  wire  _GEN_347 = 7'h2b == idx & way2[0] ? dirty_43_1 : _GEN_346; // @[cache.scala 72:{64,64}]
  wire  _GEN_2187 = 7'h2c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_348 = 7'h2c == idx & ~way2[0] ? dirty_44_0 : _GEN_347; // @[cache.scala 72:{64,64}]
  wire  _GEN_349 = 7'h2c == idx & way2[0] ? dirty_44_1 : _GEN_348; // @[cache.scala 72:{64,64}]
  wire  _GEN_2190 = 7'h2d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_350 = 7'h2d == idx & ~way2[0] ? dirty_45_0 : _GEN_349; // @[cache.scala 72:{64,64}]
  wire  _GEN_351 = 7'h2d == idx & way2[0] ? dirty_45_1 : _GEN_350; // @[cache.scala 72:{64,64}]
  wire  _GEN_2193 = 7'h2e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_352 = 7'h2e == idx & ~way2[0] ? dirty_46_0 : _GEN_351; // @[cache.scala 72:{64,64}]
  wire  _GEN_353 = 7'h2e == idx & way2[0] ? dirty_46_1 : _GEN_352; // @[cache.scala 72:{64,64}]
  wire  _GEN_2196 = 7'h2f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_354 = 7'h2f == idx & ~way2[0] ? dirty_47_0 : _GEN_353; // @[cache.scala 72:{64,64}]
  wire  _GEN_355 = 7'h2f == idx & way2[0] ? dirty_47_1 : _GEN_354; // @[cache.scala 72:{64,64}]
  wire  _GEN_2199 = 7'h30 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_356 = 7'h30 == idx & ~way2[0] ? dirty_48_0 : _GEN_355; // @[cache.scala 72:{64,64}]
  wire  _GEN_357 = 7'h30 == idx & way2[0] ? dirty_48_1 : _GEN_356; // @[cache.scala 72:{64,64}]
  wire  _GEN_2202 = 7'h31 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_358 = 7'h31 == idx & ~way2[0] ? dirty_49_0 : _GEN_357; // @[cache.scala 72:{64,64}]
  wire  _GEN_359 = 7'h31 == idx & way2[0] ? dirty_49_1 : _GEN_358; // @[cache.scala 72:{64,64}]
  wire  _GEN_2205 = 7'h32 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_360 = 7'h32 == idx & ~way2[0] ? dirty_50_0 : _GEN_359; // @[cache.scala 72:{64,64}]
  wire  _GEN_361 = 7'h32 == idx & way2[0] ? dirty_50_1 : _GEN_360; // @[cache.scala 72:{64,64}]
  wire  _GEN_2208 = 7'h33 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_362 = 7'h33 == idx & ~way2[0] ? dirty_51_0 : _GEN_361; // @[cache.scala 72:{64,64}]
  wire  _GEN_363 = 7'h33 == idx & way2[0] ? dirty_51_1 : _GEN_362; // @[cache.scala 72:{64,64}]
  wire  _GEN_2211 = 7'h34 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_364 = 7'h34 == idx & ~way2[0] ? dirty_52_0 : _GEN_363; // @[cache.scala 72:{64,64}]
  wire  _GEN_365 = 7'h34 == idx & way2[0] ? dirty_52_1 : _GEN_364; // @[cache.scala 72:{64,64}]
  wire  _GEN_2214 = 7'h35 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_366 = 7'h35 == idx & ~way2[0] ? dirty_53_0 : _GEN_365; // @[cache.scala 72:{64,64}]
  wire  _GEN_367 = 7'h35 == idx & way2[0] ? dirty_53_1 : _GEN_366; // @[cache.scala 72:{64,64}]
  wire  _GEN_2217 = 7'h36 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_368 = 7'h36 == idx & ~way2[0] ? dirty_54_0 : _GEN_367; // @[cache.scala 72:{64,64}]
  wire  _GEN_369 = 7'h36 == idx & way2[0] ? dirty_54_1 : _GEN_368; // @[cache.scala 72:{64,64}]
  wire  _GEN_2220 = 7'h37 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_370 = 7'h37 == idx & ~way2[0] ? dirty_55_0 : _GEN_369; // @[cache.scala 72:{64,64}]
  wire  _GEN_371 = 7'h37 == idx & way2[0] ? dirty_55_1 : _GEN_370; // @[cache.scala 72:{64,64}]
  wire  _GEN_2223 = 7'h38 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_372 = 7'h38 == idx & ~way2[0] ? dirty_56_0 : _GEN_371; // @[cache.scala 72:{64,64}]
  wire  _GEN_373 = 7'h38 == idx & way2[0] ? dirty_56_1 : _GEN_372; // @[cache.scala 72:{64,64}]
  wire  _GEN_2226 = 7'h39 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_374 = 7'h39 == idx & ~way2[0] ? dirty_57_0 : _GEN_373; // @[cache.scala 72:{64,64}]
  wire  _GEN_375 = 7'h39 == idx & way2[0] ? dirty_57_1 : _GEN_374; // @[cache.scala 72:{64,64}]
  wire  _GEN_2229 = 7'h3a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_376 = 7'h3a == idx & ~way2[0] ? dirty_58_0 : _GEN_375; // @[cache.scala 72:{64,64}]
  wire  _GEN_377 = 7'h3a == idx & way2[0] ? dirty_58_1 : _GEN_376; // @[cache.scala 72:{64,64}]
  wire  _GEN_2232 = 7'h3b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_378 = 7'h3b == idx & ~way2[0] ? dirty_59_0 : _GEN_377; // @[cache.scala 72:{64,64}]
  wire  _GEN_379 = 7'h3b == idx & way2[0] ? dirty_59_1 : _GEN_378; // @[cache.scala 72:{64,64}]
  wire  _GEN_2235 = 7'h3c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_380 = 7'h3c == idx & ~way2[0] ? dirty_60_0 : _GEN_379; // @[cache.scala 72:{64,64}]
  wire  _GEN_381 = 7'h3c == idx & way2[0] ? dirty_60_1 : _GEN_380; // @[cache.scala 72:{64,64}]
  wire  _GEN_2238 = 7'h3d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_382 = 7'h3d == idx & ~way2[0] ? dirty_61_0 : _GEN_381; // @[cache.scala 72:{64,64}]
  wire  _GEN_383 = 7'h3d == idx & way2[0] ? dirty_61_1 : _GEN_382; // @[cache.scala 72:{64,64}]
  wire  _GEN_2241 = 7'h3e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_384 = 7'h3e == idx & ~way2[0] ? dirty_62_0 : _GEN_383; // @[cache.scala 72:{64,64}]
  wire  _GEN_385 = 7'h3e == idx & way2[0] ? dirty_62_1 : _GEN_384; // @[cache.scala 72:{64,64}]
  wire  _GEN_2244 = 7'h3f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_386 = 7'h3f == idx & ~way2[0] ? dirty_63_0 : _GEN_385; // @[cache.scala 72:{64,64}]
  wire  _GEN_387 = 7'h3f == idx & way2[0] ? dirty_63_1 : _GEN_386; // @[cache.scala 72:{64,64}]
  wire  _GEN_2247 = 7'h40 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_388 = 7'h40 == idx & ~way2[0] ? dirty_64_0 : _GEN_387; // @[cache.scala 72:{64,64}]
  wire  _GEN_389 = 7'h40 == idx & way2[0] ? dirty_64_1 : _GEN_388; // @[cache.scala 72:{64,64}]
  wire  _GEN_2250 = 7'h41 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_390 = 7'h41 == idx & ~way2[0] ? dirty_65_0 : _GEN_389; // @[cache.scala 72:{64,64}]
  wire  _GEN_391 = 7'h41 == idx & way2[0] ? dirty_65_1 : _GEN_390; // @[cache.scala 72:{64,64}]
  wire  _GEN_2253 = 7'h42 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_392 = 7'h42 == idx & ~way2[0] ? dirty_66_0 : _GEN_391; // @[cache.scala 72:{64,64}]
  wire  _GEN_393 = 7'h42 == idx & way2[0] ? dirty_66_1 : _GEN_392; // @[cache.scala 72:{64,64}]
  wire  _GEN_2256 = 7'h43 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_394 = 7'h43 == idx & ~way2[0] ? dirty_67_0 : _GEN_393; // @[cache.scala 72:{64,64}]
  wire  _GEN_395 = 7'h43 == idx & way2[0] ? dirty_67_1 : _GEN_394; // @[cache.scala 72:{64,64}]
  wire  _GEN_2259 = 7'h44 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_396 = 7'h44 == idx & ~way2[0] ? dirty_68_0 : _GEN_395; // @[cache.scala 72:{64,64}]
  wire  _GEN_397 = 7'h44 == idx & way2[0] ? dirty_68_1 : _GEN_396; // @[cache.scala 72:{64,64}]
  wire  _GEN_2262 = 7'h45 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_398 = 7'h45 == idx & ~way2[0] ? dirty_69_0 : _GEN_397; // @[cache.scala 72:{64,64}]
  wire  _GEN_399 = 7'h45 == idx & way2[0] ? dirty_69_1 : _GEN_398; // @[cache.scala 72:{64,64}]
  wire  _GEN_2265 = 7'h46 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_400 = 7'h46 == idx & ~way2[0] ? dirty_70_0 : _GEN_399; // @[cache.scala 72:{64,64}]
  wire  _GEN_401 = 7'h46 == idx & way2[0] ? dirty_70_1 : _GEN_400; // @[cache.scala 72:{64,64}]
  wire  _GEN_2268 = 7'h47 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_402 = 7'h47 == idx & ~way2[0] ? dirty_71_0 : _GEN_401; // @[cache.scala 72:{64,64}]
  wire  _GEN_403 = 7'h47 == idx & way2[0] ? dirty_71_1 : _GEN_402; // @[cache.scala 72:{64,64}]
  wire  _GEN_2271 = 7'h48 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_404 = 7'h48 == idx & ~way2[0] ? dirty_72_0 : _GEN_403; // @[cache.scala 72:{64,64}]
  wire  _GEN_405 = 7'h48 == idx & way2[0] ? dirty_72_1 : _GEN_404; // @[cache.scala 72:{64,64}]
  wire  _GEN_2274 = 7'h49 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_406 = 7'h49 == idx & ~way2[0] ? dirty_73_0 : _GEN_405; // @[cache.scala 72:{64,64}]
  wire  _GEN_407 = 7'h49 == idx & way2[0] ? dirty_73_1 : _GEN_406; // @[cache.scala 72:{64,64}]
  wire  _GEN_2277 = 7'h4a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_408 = 7'h4a == idx & ~way2[0] ? dirty_74_0 : _GEN_407; // @[cache.scala 72:{64,64}]
  wire  _GEN_409 = 7'h4a == idx & way2[0] ? dirty_74_1 : _GEN_408; // @[cache.scala 72:{64,64}]
  wire  _GEN_2280 = 7'h4b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_410 = 7'h4b == idx & ~way2[0] ? dirty_75_0 : _GEN_409; // @[cache.scala 72:{64,64}]
  wire  _GEN_411 = 7'h4b == idx & way2[0] ? dirty_75_1 : _GEN_410; // @[cache.scala 72:{64,64}]
  wire  _GEN_2283 = 7'h4c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_412 = 7'h4c == idx & ~way2[0] ? dirty_76_0 : _GEN_411; // @[cache.scala 72:{64,64}]
  wire  _GEN_413 = 7'h4c == idx & way2[0] ? dirty_76_1 : _GEN_412; // @[cache.scala 72:{64,64}]
  wire  _GEN_2286 = 7'h4d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_414 = 7'h4d == idx & ~way2[0] ? dirty_77_0 : _GEN_413; // @[cache.scala 72:{64,64}]
  wire  _GEN_415 = 7'h4d == idx & way2[0] ? dirty_77_1 : _GEN_414; // @[cache.scala 72:{64,64}]
  wire  _GEN_2289 = 7'h4e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_416 = 7'h4e == idx & ~way2[0] ? dirty_78_0 : _GEN_415; // @[cache.scala 72:{64,64}]
  wire  _GEN_417 = 7'h4e == idx & way2[0] ? dirty_78_1 : _GEN_416; // @[cache.scala 72:{64,64}]
  wire  _GEN_2292 = 7'h4f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_418 = 7'h4f == idx & ~way2[0] ? dirty_79_0 : _GEN_417; // @[cache.scala 72:{64,64}]
  wire  _GEN_419 = 7'h4f == idx & way2[0] ? dirty_79_1 : _GEN_418; // @[cache.scala 72:{64,64}]
  wire  _GEN_2295 = 7'h50 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_420 = 7'h50 == idx & ~way2[0] ? dirty_80_0 : _GEN_419; // @[cache.scala 72:{64,64}]
  wire  _GEN_421 = 7'h50 == idx & way2[0] ? dirty_80_1 : _GEN_420; // @[cache.scala 72:{64,64}]
  wire  _GEN_2298 = 7'h51 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_422 = 7'h51 == idx & ~way2[0] ? dirty_81_0 : _GEN_421; // @[cache.scala 72:{64,64}]
  wire  _GEN_423 = 7'h51 == idx & way2[0] ? dirty_81_1 : _GEN_422; // @[cache.scala 72:{64,64}]
  wire  _GEN_2301 = 7'h52 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_424 = 7'h52 == idx & ~way2[0] ? dirty_82_0 : _GEN_423; // @[cache.scala 72:{64,64}]
  wire  _GEN_425 = 7'h52 == idx & way2[0] ? dirty_82_1 : _GEN_424; // @[cache.scala 72:{64,64}]
  wire  _GEN_2304 = 7'h53 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_426 = 7'h53 == idx & ~way2[0] ? dirty_83_0 : _GEN_425; // @[cache.scala 72:{64,64}]
  wire  _GEN_427 = 7'h53 == idx & way2[0] ? dirty_83_1 : _GEN_426; // @[cache.scala 72:{64,64}]
  wire  _GEN_2307 = 7'h54 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_428 = 7'h54 == idx & ~way2[0] ? dirty_84_0 : _GEN_427; // @[cache.scala 72:{64,64}]
  wire  _GEN_429 = 7'h54 == idx & way2[0] ? dirty_84_1 : _GEN_428; // @[cache.scala 72:{64,64}]
  wire  _GEN_2310 = 7'h55 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_430 = 7'h55 == idx & ~way2[0] ? dirty_85_0 : _GEN_429; // @[cache.scala 72:{64,64}]
  wire  _GEN_431 = 7'h55 == idx & way2[0] ? dirty_85_1 : _GEN_430; // @[cache.scala 72:{64,64}]
  wire  _GEN_2313 = 7'h56 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_432 = 7'h56 == idx & ~way2[0] ? dirty_86_0 : _GEN_431; // @[cache.scala 72:{64,64}]
  wire  _GEN_433 = 7'h56 == idx & way2[0] ? dirty_86_1 : _GEN_432; // @[cache.scala 72:{64,64}]
  wire  _GEN_2316 = 7'h57 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_434 = 7'h57 == idx & ~way2[0] ? dirty_87_0 : _GEN_433; // @[cache.scala 72:{64,64}]
  wire  _GEN_435 = 7'h57 == idx & way2[0] ? dirty_87_1 : _GEN_434; // @[cache.scala 72:{64,64}]
  wire  _GEN_2319 = 7'h58 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_436 = 7'h58 == idx & ~way2[0] ? dirty_88_0 : _GEN_435; // @[cache.scala 72:{64,64}]
  wire  _GEN_437 = 7'h58 == idx & way2[0] ? dirty_88_1 : _GEN_436; // @[cache.scala 72:{64,64}]
  wire  _GEN_2322 = 7'h59 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_438 = 7'h59 == idx & ~way2[0] ? dirty_89_0 : _GEN_437; // @[cache.scala 72:{64,64}]
  wire  _GEN_439 = 7'h59 == idx & way2[0] ? dirty_89_1 : _GEN_438; // @[cache.scala 72:{64,64}]
  wire  _GEN_2325 = 7'h5a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_440 = 7'h5a == idx & ~way2[0] ? dirty_90_0 : _GEN_439; // @[cache.scala 72:{64,64}]
  wire  _GEN_441 = 7'h5a == idx & way2[0] ? dirty_90_1 : _GEN_440; // @[cache.scala 72:{64,64}]
  wire  _GEN_2328 = 7'h5b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_442 = 7'h5b == idx & ~way2[0] ? dirty_91_0 : _GEN_441; // @[cache.scala 72:{64,64}]
  wire  _GEN_443 = 7'h5b == idx & way2[0] ? dirty_91_1 : _GEN_442; // @[cache.scala 72:{64,64}]
  wire  _GEN_2331 = 7'h5c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_444 = 7'h5c == idx & ~way2[0] ? dirty_92_0 : _GEN_443; // @[cache.scala 72:{64,64}]
  wire  _GEN_445 = 7'h5c == idx & way2[0] ? dirty_92_1 : _GEN_444; // @[cache.scala 72:{64,64}]
  wire  _GEN_2334 = 7'h5d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_446 = 7'h5d == idx & ~way2[0] ? dirty_93_0 : _GEN_445; // @[cache.scala 72:{64,64}]
  wire  _GEN_447 = 7'h5d == idx & way2[0] ? dirty_93_1 : _GEN_446; // @[cache.scala 72:{64,64}]
  wire  _GEN_2337 = 7'h5e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_448 = 7'h5e == idx & ~way2[0] ? dirty_94_0 : _GEN_447; // @[cache.scala 72:{64,64}]
  wire  _GEN_449 = 7'h5e == idx & way2[0] ? dirty_94_1 : _GEN_448; // @[cache.scala 72:{64,64}]
  wire  _GEN_2340 = 7'h5f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_450 = 7'h5f == idx & ~way2[0] ? dirty_95_0 : _GEN_449; // @[cache.scala 72:{64,64}]
  wire  _GEN_451 = 7'h5f == idx & way2[0] ? dirty_95_1 : _GEN_450; // @[cache.scala 72:{64,64}]
  wire  _GEN_2343 = 7'h60 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_452 = 7'h60 == idx & ~way2[0] ? dirty_96_0 : _GEN_451; // @[cache.scala 72:{64,64}]
  wire  _GEN_453 = 7'h60 == idx & way2[0] ? dirty_96_1 : _GEN_452; // @[cache.scala 72:{64,64}]
  wire  _GEN_2346 = 7'h61 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_454 = 7'h61 == idx & ~way2[0] ? dirty_97_0 : _GEN_453; // @[cache.scala 72:{64,64}]
  wire  _GEN_455 = 7'h61 == idx & way2[0] ? dirty_97_1 : _GEN_454; // @[cache.scala 72:{64,64}]
  wire  _GEN_2349 = 7'h62 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_456 = 7'h62 == idx & ~way2[0] ? dirty_98_0 : _GEN_455; // @[cache.scala 72:{64,64}]
  wire  _GEN_457 = 7'h62 == idx & way2[0] ? dirty_98_1 : _GEN_456; // @[cache.scala 72:{64,64}]
  wire  _GEN_2352 = 7'h63 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_458 = 7'h63 == idx & ~way2[0] ? dirty_99_0 : _GEN_457; // @[cache.scala 72:{64,64}]
  wire  _GEN_459 = 7'h63 == idx & way2[0] ? dirty_99_1 : _GEN_458; // @[cache.scala 72:{64,64}]
  wire  _GEN_2355 = 7'h64 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_460 = 7'h64 == idx & ~way2[0] ? dirty_100_0 : _GEN_459; // @[cache.scala 72:{64,64}]
  wire  _GEN_461 = 7'h64 == idx & way2[0] ? dirty_100_1 : _GEN_460; // @[cache.scala 72:{64,64}]
  wire  _GEN_2358 = 7'h65 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_462 = 7'h65 == idx & ~way2[0] ? dirty_101_0 : _GEN_461; // @[cache.scala 72:{64,64}]
  wire  _GEN_463 = 7'h65 == idx & way2[0] ? dirty_101_1 : _GEN_462; // @[cache.scala 72:{64,64}]
  wire  _GEN_2361 = 7'h66 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_464 = 7'h66 == idx & ~way2[0] ? dirty_102_0 : _GEN_463; // @[cache.scala 72:{64,64}]
  wire  _GEN_465 = 7'h66 == idx & way2[0] ? dirty_102_1 : _GEN_464; // @[cache.scala 72:{64,64}]
  wire  _GEN_2364 = 7'h67 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_466 = 7'h67 == idx & ~way2[0] ? dirty_103_0 : _GEN_465; // @[cache.scala 72:{64,64}]
  wire  _GEN_467 = 7'h67 == idx & way2[0] ? dirty_103_1 : _GEN_466; // @[cache.scala 72:{64,64}]
  wire  _GEN_2367 = 7'h68 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_468 = 7'h68 == idx & ~way2[0] ? dirty_104_0 : _GEN_467; // @[cache.scala 72:{64,64}]
  wire  _GEN_469 = 7'h68 == idx & way2[0] ? dirty_104_1 : _GEN_468; // @[cache.scala 72:{64,64}]
  wire  _GEN_2370 = 7'h69 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_470 = 7'h69 == idx & ~way2[0] ? dirty_105_0 : _GEN_469; // @[cache.scala 72:{64,64}]
  wire  _GEN_471 = 7'h69 == idx & way2[0] ? dirty_105_1 : _GEN_470; // @[cache.scala 72:{64,64}]
  wire  _GEN_2373 = 7'h6a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_472 = 7'h6a == idx & ~way2[0] ? dirty_106_0 : _GEN_471; // @[cache.scala 72:{64,64}]
  wire  _GEN_473 = 7'h6a == idx & way2[0] ? dirty_106_1 : _GEN_472; // @[cache.scala 72:{64,64}]
  wire  _GEN_2376 = 7'h6b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_474 = 7'h6b == idx & ~way2[0] ? dirty_107_0 : _GEN_473; // @[cache.scala 72:{64,64}]
  wire  _GEN_475 = 7'h6b == idx & way2[0] ? dirty_107_1 : _GEN_474; // @[cache.scala 72:{64,64}]
  wire  _GEN_2379 = 7'h6c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_476 = 7'h6c == idx & ~way2[0] ? dirty_108_0 : _GEN_475; // @[cache.scala 72:{64,64}]
  wire  _GEN_477 = 7'h6c == idx & way2[0] ? dirty_108_1 : _GEN_476; // @[cache.scala 72:{64,64}]
  wire  _GEN_2382 = 7'h6d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_478 = 7'h6d == idx & ~way2[0] ? dirty_109_0 : _GEN_477; // @[cache.scala 72:{64,64}]
  wire  _GEN_479 = 7'h6d == idx & way2[0] ? dirty_109_1 : _GEN_478; // @[cache.scala 72:{64,64}]
  wire  _GEN_2385 = 7'h6e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_480 = 7'h6e == idx & ~way2[0] ? dirty_110_0 : _GEN_479; // @[cache.scala 72:{64,64}]
  wire  _GEN_481 = 7'h6e == idx & way2[0] ? dirty_110_1 : _GEN_480; // @[cache.scala 72:{64,64}]
  wire  _GEN_2388 = 7'h6f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_482 = 7'h6f == idx & ~way2[0] ? dirty_111_0 : _GEN_481; // @[cache.scala 72:{64,64}]
  wire  _GEN_483 = 7'h6f == idx & way2[0] ? dirty_111_1 : _GEN_482; // @[cache.scala 72:{64,64}]
  wire  _GEN_2391 = 7'h70 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_484 = 7'h70 == idx & ~way2[0] ? dirty_112_0 : _GEN_483; // @[cache.scala 72:{64,64}]
  wire  _GEN_485 = 7'h70 == idx & way2[0] ? dirty_112_1 : _GEN_484; // @[cache.scala 72:{64,64}]
  wire  _GEN_2394 = 7'h71 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_486 = 7'h71 == idx & ~way2[0] ? dirty_113_0 : _GEN_485; // @[cache.scala 72:{64,64}]
  wire  _GEN_487 = 7'h71 == idx & way2[0] ? dirty_113_1 : _GEN_486; // @[cache.scala 72:{64,64}]
  wire  _GEN_2397 = 7'h72 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_488 = 7'h72 == idx & ~way2[0] ? dirty_114_0 : _GEN_487; // @[cache.scala 72:{64,64}]
  wire  _GEN_489 = 7'h72 == idx & way2[0] ? dirty_114_1 : _GEN_488; // @[cache.scala 72:{64,64}]
  wire  _GEN_2400 = 7'h73 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_490 = 7'h73 == idx & ~way2[0] ? dirty_115_0 : _GEN_489; // @[cache.scala 72:{64,64}]
  wire  _GEN_491 = 7'h73 == idx & way2[0] ? dirty_115_1 : _GEN_490; // @[cache.scala 72:{64,64}]
  wire  _GEN_2403 = 7'h74 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_492 = 7'h74 == idx & ~way2[0] ? dirty_116_0 : _GEN_491; // @[cache.scala 72:{64,64}]
  wire  _GEN_493 = 7'h74 == idx & way2[0] ? dirty_116_1 : _GEN_492; // @[cache.scala 72:{64,64}]
  wire  _GEN_2406 = 7'h75 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_494 = 7'h75 == idx & ~way2[0] ? dirty_117_0 : _GEN_493; // @[cache.scala 72:{64,64}]
  wire  _GEN_495 = 7'h75 == idx & way2[0] ? dirty_117_1 : _GEN_494; // @[cache.scala 72:{64,64}]
  wire  _GEN_2409 = 7'h76 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_496 = 7'h76 == idx & ~way2[0] ? dirty_118_0 : _GEN_495; // @[cache.scala 72:{64,64}]
  wire  _GEN_497 = 7'h76 == idx & way2[0] ? dirty_118_1 : _GEN_496; // @[cache.scala 72:{64,64}]
  wire  _GEN_2412 = 7'h77 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_498 = 7'h77 == idx & ~way2[0] ? dirty_119_0 : _GEN_497; // @[cache.scala 72:{64,64}]
  wire  _GEN_499 = 7'h77 == idx & way2[0] ? dirty_119_1 : _GEN_498; // @[cache.scala 72:{64,64}]
  wire  _GEN_2415 = 7'h78 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_500 = 7'h78 == idx & ~way2[0] ? dirty_120_0 : _GEN_499; // @[cache.scala 72:{64,64}]
  wire  _GEN_501 = 7'h78 == idx & way2[0] ? dirty_120_1 : _GEN_500; // @[cache.scala 72:{64,64}]
  wire  _GEN_2418 = 7'h79 == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_502 = 7'h79 == idx & ~way2[0] ? dirty_121_0 : _GEN_501; // @[cache.scala 72:{64,64}]
  wire  _GEN_503 = 7'h79 == idx & way2[0] ? dirty_121_1 : _GEN_502; // @[cache.scala 72:{64,64}]
  wire  _GEN_2421 = 7'h7a == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_504 = 7'h7a == idx & ~way2[0] ? dirty_122_0 : _GEN_503; // @[cache.scala 72:{64,64}]
  wire  _GEN_505 = 7'h7a == idx & way2[0] ? dirty_122_1 : _GEN_504; // @[cache.scala 72:{64,64}]
  wire  _GEN_2424 = 7'h7b == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_506 = 7'h7b == idx & ~way2[0] ? dirty_123_0 : _GEN_505; // @[cache.scala 72:{64,64}]
  wire  _GEN_507 = 7'h7b == idx & way2[0] ? dirty_123_1 : _GEN_506; // @[cache.scala 72:{64,64}]
  wire  _GEN_2427 = 7'h7c == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_508 = 7'h7c == idx & ~way2[0] ? dirty_124_0 : _GEN_507; // @[cache.scala 72:{64,64}]
  wire  _GEN_509 = 7'h7c == idx & way2[0] ? dirty_124_1 : _GEN_508; // @[cache.scala 72:{64,64}]
  wire  _GEN_2430 = 7'h7d == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_510 = 7'h7d == idx & ~way2[0] ? dirty_125_0 : _GEN_509; // @[cache.scala 72:{64,64}]
  wire  _GEN_511 = 7'h7d == idx & way2[0] ? dirty_125_1 : _GEN_510; // @[cache.scala 72:{64,64}]
  wire  _GEN_2433 = 7'h7e == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_512 = 7'h7e == idx & ~way2[0] ? dirty_126_0 : _GEN_511; // @[cache.scala 72:{64,64}]
  wire  _GEN_513 = 7'h7e == idx & way2[0] ? dirty_126_1 : _GEN_512; // @[cache.scala 72:{64,64}]
  wire  _GEN_2436 = 7'h7f == idx; // @[cache.scala 72:{64,64}]
  wire  _GEN_514 = 7'h7f == idx & ~way2[0] ? dirty_127_0 : _GEN_513; // @[cache.scala 72:{64,64}]
  wire  _GEN_515 = 7'h7f == idx & way2[0] ? dirty_127_1 : _GEN_514; // @[cache.scala 72:{64,64}]
  wire [3:0] _state_T_17 = 4'h0 == state ? _state_T_3 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _state_T_19 = 4'h1 == state ? 4'h2 : _state_T_17; // @[Mux.scala 81:58]
  wire [3:0] _state_T_21 = 4'h2 == state ? _state_T_5 : _state_T_19; // @[Mux.scala 81:58]
  wire  _wdata_T = state == 4'h1; // @[cache.scala 78:22]
  wire  _wdata_T_1 = io_in_w_ready & io_in_w_valid; // @[Decoupled.scala 52:35]
  wire  _wdata_T_2 = state == 4'h1 & _wdata_T_1; // @[cache.scala 78:34]
  wire  _io_in_r_bits_data_T = state == 4'h3; // @[cache.scala 81:34]
  wire [127:0] _io_in_r_bits_data_T_1 = io_ram_bits_Q >> offset; // @[cache.scala 81:58]
  wire  _io_in_r_bits_data_T_3 = state == 4'h5; // @[cache.scala 82:34]
  wire [127:0] _io_in_r_bits_data_T_4 = buf_ >> offset; // @[cache.scala 82:52]
  wire [127:0] _io_in_r_bits_data_T_5 = state == 4'h5 ? _io_in_r_bits_data_T_4 : 128'h0; // @[cache.scala 82:27]
  wire [127:0] _io_in_r_bits_data_T_6 = state == 4'h3 ? {{64'd0}, _io_in_r_bits_data_T_1[63:0]} : _io_in_r_bits_data_T_5
    ; // @[cache.scala 81:27]
  wire  _state_r_T = state == 4'h4; // @[cache.scala 99:27]
  wire  _state_r_T_1 = io_mem_ar_ready & io_mem_ar_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _state_r_T_3 = state == 4'h4 & _state_r_T_1 ? 4'h6 : 4'h0; // @[cache.scala 99:20]
  wire  _state_r_T_4 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _state_r_T_5 = _state_r_T_4 ? 4'h7 : 4'h6; // @[cache.scala 100:26]
  wire [3:0] _state_r_T_11 = 4'h0 == state_r ? _state_r_T_3 : 4'h0; // @[Mux.scala 81:58]
  wire  _state_w_T_1 = io_mem_aw_ready & io_mem_aw_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _state_w_T_3 = _state_r_T & _state_w_T_1 ? 4'h1 : 4'h0; // @[cache.scala 109:20]
  wire  _state_w_T_4 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _state_w_T_5 = _state_w_T_4 ? 4'h7 : 4'h6; // @[cache.scala 111:26]
  wire  _state_w_T_6 = io_mem_b_ready & io_mem_b_valid; // @[Decoupled.scala 52:35]
  wire [3:0] _state_w_T_11 = 4'h0 == state_w ? _state_w_T_3 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _state_w_T_13 = 4'h1 == state_w ? 4'h6 : _state_w_T_11; // @[Mux.scala 81:58]
  wire [27:0] _io_mem_aw_bits_addr_T = {tag_way, 7'h0}; // @[cache.scala 116:35]
  wire [27:0] _GEN_2821 = {{21'd0}, idx}; // @[cache.scala 116:48]
  wire [27:0] _io_mem_aw_bits_addr_T_1 = _io_mem_aw_bits_addr_T | _GEN_2821; // @[cache.scala 116:48]
  wire  _io_mem_w_bits_data_T = state_w == 4'h7; // @[cache.scala 125:37]
  wire [34:0] _GEN_3204 = {{3'd0}, addr}; // @[cache.scala 131:31]
  wire [34:0] _io_mem_ar_bits_addr_T_2 = _GEN_3204 & 35'h7fffffff8; // @[cache.scala 131:31]
  wire  _io_mem_ar_valid_T = state_r == 4'h0; // @[cache.scala 132:30]
  reg  rcnt; // @[cache.scala 138:21]
  wire  _buf_T_1 = ~_state_r_T_4; // @[cache.scala 144:5]
  wire [127:0] _buf_T_5 = {buf_[127:64],io_mem_r_bits_data}; // @[Cat.scala 33:92]
  wire [127:0] _buf_T_7 = {io_mem_r_bits_data,buf_[63:0]}; // @[Cat.scala 33:92]
  reg [41:0] taggg; // @[cache.scala 150:22]
  wire [41:0] _tagg_T_2 = {taggg[41:21],tag}; // @[Cat.scala 33:92]
  wire [41:0] _tagg_T_4 = {tag,taggg[20:0]}; // @[Cat.scala 33:92]
  wire  _GEN_1034 = _GEN_2057 & way2[0] ? valid_0_1 : valid_0_0; // @[cache.scala 154:{26,26}]
  wire  _GEN_1035 = _GEN_2058 & _GEN_2059 ? valid_1_0 : _GEN_1034; // @[cache.scala 154:{26,26}]
  wire  _GEN_1036 = _GEN_2058 & way2[0] ? valid_1_1 : _GEN_1035; // @[cache.scala 154:{26,26}]
  wire  _GEN_1037 = _GEN_2061 & _GEN_2059 ? valid_2_0 : _GEN_1036; // @[cache.scala 154:{26,26}]
  wire  _GEN_1038 = _GEN_2061 & way2[0] ? valid_2_1 : _GEN_1037; // @[cache.scala 154:{26,26}]
  wire  _GEN_1039 = _GEN_2064 & _GEN_2059 ? valid_3_0 : _GEN_1038; // @[cache.scala 154:{26,26}]
  wire  _GEN_1040 = _GEN_2064 & way2[0] ? valid_3_1 : _GEN_1039; // @[cache.scala 154:{26,26}]
  wire  _GEN_1041 = _GEN_2067 & _GEN_2059 ? valid_4_0 : _GEN_1040; // @[cache.scala 154:{26,26}]
  wire  _GEN_1042 = _GEN_2067 & way2[0] ? valid_4_1 : _GEN_1041; // @[cache.scala 154:{26,26}]
  wire  _GEN_1043 = _GEN_2070 & _GEN_2059 ? valid_5_0 : _GEN_1042; // @[cache.scala 154:{26,26}]
  wire  _GEN_1044 = _GEN_2070 & way2[0] ? valid_5_1 : _GEN_1043; // @[cache.scala 154:{26,26}]
  wire  _GEN_1045 = _GEN_2073 & _GEN_2059 ? valid_6_0 : _GEN_1044; // @[cache.scala 154:{26,26}]
  wire  _GEN_1046 = _GEN_2073 & way2[0] ? valid_6_1 : _GEN_1045; // @[cache.scala 154:{26,26}]
  wire  _GEN_1047 = _GEN_2076 & _GEN_2059 ? valid_7_0 : _GEN_1046; // @[cache.scala 154:{26,26}]
  wire  _GEN_1048 = _GEN_2076 & way2[0] ? valid_7_1 : _GEN_1047; // @[cache.scala 154:{26,26}]
  wire  _GEN_1049 = _GEN_2079 & _GEN_2059 ? valid_8_0 : _GEN_1048; // @[cache.scala 154:{26,26}]
  wire  _GEN_1050 = _GEN_2079 & way2[0] ? valid_8_1 : _GEN_1049; // @[cache.scala 154:{26,26}]
  wire  _GEN_1051 = _GEN_2082 & _GEN_2059 ? valid_9_0 : _GEN_1050; // @[cache.scala 154:{26,26}]
  wire  _GEN_1052 = _GEN_2082 & way2[0] ? valid_9_1 : _GEN_1051; // @[cache.scala 154:{26,26}]
  wire  _GEN_1053 = _GEN_2085 & _GEN_2059 ? valid_10_0 : _GEN_1052; // @[cache.scala 154:{26,26}]
  wire  _GEN_1054 = _GEN_2085 & way2[0] ? valid_10_1 : _GEN_1053; // @[cache.scala 154:{26,26}]
  wire  _GEN_1055 = _GEN_2088 & _GEN_2059 ? valid_11_0 : _GEN_1054; // @[cache.scala 154:{26,26}]
  wire  _GEN_1056 = _GEN_2088 & way2[0] ? valid_11_1 : _GEN_1055; // @[cache.scala 154:{26,26}]
  wire  _GEN_1057 = _GEN_2091 & _GEN_2059 ? valid_12_0 : _GEN_1056; // @[cache.scala 154:{26,26}]
  wire  _GEN_1058 = _GEN_2091 & way2[0] ? valid_12_1 : _GEN_1057; // @[cache.scala 154:{26,26}]
  wire  _GEN_1059 = _GEN_2094 & _GEN_2059 ? valid_13_0 : _GEN_1058; // @[cache.scala 154:{26,26}]
  wire  _GEN_1060 = _GEN_2094 & way2[0] ? valid_13_1 : _GEN_1059; // @[cache.scala 154:{26,26}]
  wire  _GEN_1061 = _GEN_2097 & _GEN_2059 ? valid_14_0 : _GEN_1060; // @[cache.scala 154:{26,26}]
  wire  _GEN_1062 = _GEN_2097 & way2[0] ? valid_14_1 : _GEN_1061; // @[cache.scala 154:{26,26}]
  wire  _GEN_1063 = _GEN_2100 & _GEN_2059 ? valid_15_0 : _GEN_1062; // @[cache.scala 154:{26,26}]
  wire  _GEN_1064 = _GEN_2100 & way2[0] ? valid_15_1 : _GEN_1063; // @[cache.scala 154:{26,26}]
  wire  _GEN_1065 = _GEN_2103 & _GEN_2059 ? valid_16_0 : _GEN_1064; // @[cache.scala 154:{26,26}]
  wire  _GEN_1066 = _GEN_2103 & way2[0] ? valid_16_1 : _GEN_1065; // @[cache.scala 154:{26,26}]
  wire  _GEN_1067 = _GEN_2106 & _GEN_2059 ? valid_17_0 : _GEN_1066; // @[cache.scala 154:{26,26}]
  wire  _GEN_1068 = _GEN_2106 & way2[0] ? valid_17_1 : _GEN_1067; // @[cache.scala 154:{26,26}]
  wire  _GEN_1069 = _GEN_2109 & _GEN_2059 ? valid_18_0 : _GEN_1068; // @[cache.scala 154:{26,26}]
  wire  _GEN_1070 = _GEN_2109 & way2[0] ? valid_18_1 : _GEN_1069; // @[cache.scala 154:{26,26}]
  wire  _GEN_1071 = _GEN_2112 & _GEN_2059 ? valid_19_0 : _GEN_1070; // @[cache.scala 154:{26,26}]
  wire  _GEN_1072 = _GEN_2112 & way2[0] ? valid_19_1 : _GEN_1071; // @[cache.scala 154:{26,26}]
  wire  _GEN_1073 = _GEN_2115 & _GEN_2059 ? valid_20_0 : _GEN_1072; // @[cache.scala 154:{26,26}]
  wire  _GEN_1074 = _GEN_2115 & way2[0] ? valid_20_1 : _GEN_1073; // @[cache.scala 154:{26,26}]
  wire  _GEN_1075 = _GEN_2118 & _GEN_2059 ? valid_21_0 : _GEN_1074; // @[cache.scala 154:{26,26}]
  wire  _GEN_1076 = _GEN_2118 & way2[0] ? valid_21_1 : _GEN_1075; // @[cache.scala 154:{26,26}]
  wire  _GEN_1077 = _GEN_2121 & _GEN_2059 ? valid_22_0 : _GEN_1076; // @[cache.scala 154:{26,26}]
  wire  _GEN_1078 = _GEN_2121 & way2[0] ? valid_22_1 : _GEN_1077; // @[cache.scala 154:{26,26}]
  wire  _GEN_1079 = _GEN_2124 & _GEN_2059 ? valid_23_0 : _GEN_1078; // @[cache.scala 154:{26,26}]
  wire  _GEN_1080 = _GEN_2124 & way2[0] ? valid_23_1 : _GEN_1079; // @[cache.scala 154:{26,26}]
  wire  _GEN_1081 = _GEN_2127 & _GEN_2059 ? valid_24_0 : _GEN_1080; // @[cache.scala 154:{26,26}]
  wire  _GEN_1082 = _GEN_2127 & way2[0] ? valid_24_1 : _GEN_1081; // @[cache.scala 154:{26,26}]
  wire  _GEN_1083 = _GEN_2130 & _GEN_2059 ? valid_25_0 : _GEN_1082; // @[cache.scala 154:{26,26}]
  wire  _GEN_1084 = _GEN_2130 & way2[0] ? valid_25_1 : _GEN_1083; // @[cache.scala 154:{26,26}]
  wire  _GEN_1085 = _GEN_2133 & _GEN_2059 ? valid_26_0 : _GEN_1084; // @[cache.scala 154:{26,26}]
  wire  _GEN_1086 = _GEN_2133 & way2[0] ? valid_26_1 : _GEN_1085; // @[cache.scala 154:{26,26}]
  wire  _GEN_1087 = _GEN_2136 & _GEN_2059 ? valid_27_0 : _GEN_1086; // @[cache.scala 154:{26,26}]
  wire  _GEN_1088 = _GEN_2136 & way2[0] ? valid_27_1 : _GEN_1087; // @[cache.scala 154:{26,26}]
  wire  _GEN_1089 = _GEN_2139 & _GEN_2059 ? valid_28_0 : _GEN_1088; // @[cache.scala 154:{26,26}]
  wire  _GEN_1090 = _GEN_2139 & way2[0] ? valid_28_1 : _GEN_1089; // @[cache.scala 154:{26,26}]
  wire  _GEN_1091 = _GEN_2142 & _GEN_2059 ? valid_29_0 : _GEN_1090; // @[cache.scala 154:{26,26}]
  wire  _GEN_1092 = _GEN_2142 & way2[0] ? valid_29_1 : _GEN_1091; // @[cache.scala 154:{26,26}]
  wire  _GEN_1093 = _GEN_2145 & _GEN_2059 ? valid_30_0 : _GEN_1092; // @[cache.scala 154:{26,26}]
  wire  _GEN_1094 = _GEN_2145 & way2[0] ? valid_30_1 : _GEN_1093; // @[cache.scala 154:{26,26}]
  wire  _GEN_1095 = _GEN_2148 & _GEN_2059 ? valid_31_0 : _GEN_1094; // @[cache.scala 154:{26,26}]
  wire  _GEN_1096 = _GEN_2148 & way2[0] ? valid_31_1 : _GEN_1095; // @[cache.scala 154:{26,26}]
  wire  _GEN_1097 = _GEN_2151 & _GEN_2059 ? valid_32_0 : _GEN_1096; // @[cache.scala 154:{26,26}]
  wire  _GEN_1098 = _GEN_2151 & way2[0] ? valid_32_1 : _GEN_1097; // @[cache.scala 154:{26,26}]
  wire  _GEN_1099 = _GEN_2154 & _GEN_2059 ? valid_33_0 : _GEN_1098; // @[cache.scala 154:{26,26}]
  wire  _GEN_1100 = _GEN_2154 & way2[0] ? valid_33_1 : _GEN_1099; // @[cache.scala 154:{26,26}]
  wire  _GEN_1101 = _GEN_2157 & _GEN_2059 ? valid_34_0 : _GEN_1100; // @[cache.scala 154:{26,26}]
  wire  _GEN_1102 = _GEN_2157 & way2[0] ? valid_34_1 : _GEN_1101; // @[cache.scala 154:{26,26}]
  wire  _GEN_1103 = _GEN_2160 & _GEN_2059 ? valid_35_0 : _GEN_1102; // @[cache.scala 154:{26,26}]
  wire  _GEN_1104 = _GEN_2160 & way2[0] ? valid_35_1 : _GEN_1103; // @[cache.scala 154:{26,26}]
  wire  _GEN_1105 = _GEN_2163 & _GEN_2059 ? valid_36_0 : _GEN_1104; // @[cache.scala 154:{26,26}]
  wire  _GEN_1106 = _GEN_2163 & way2[0] ? valid_36_1 : _GEN_1105; // @[cache.scala 154:{26,26}]
  wire  _GEN_1107 = _GEN_2166 & _GEN_2059 ? valid_37_0 : _GEN_1106; // @[cache.scala 154:{26,26}]
  wire  _GEN_1108 = _GEN_2166 & way2[0] ? valid_37_1 : _GEN_1107; // @[cache.scala 154:{26,26}]
  wire  _GEN_1109 = _GEN_2169 & _GEN_2059 ? valid_38_0 : _GEN_1108; // @[cache.scala 154:{26,26}]
  wire  _GEN_1110 = _GEN_2169 & way2[0] ? valid_38_1 : _GEN_1109; // @[cache.scala 154:{26,26}]
  wire  _GEN_1111 = _GEN_2172 & _GEN_2059 ? valid_39_0 : _GEN_1110; // @[cache.scala 154:{26,26}]
  wire  _GEN_1112 = _GEN_2172 & way2[0] ? valid_39_1 : _GEN_1111; // @[cache.scala 154:{26,26}]
  wire  _GEN_1113 = _GEN_2175 & _GEN_2059 ? valid_40_0 : _GEN_1112; // @[cache.scala 154:{26,26}]
  wire  _GEN_1114 = _GEN_2175 & way2[0] ? valid_40_1 : _GEN_1113; // @[cache.scala 154:{26,26}]
  wire  _GEN_1115 = _GEN_2178 & _GEN_2059 ? valid_41_0 : _GEN_1114; // @[cache.scala 154:{26,26}]
  wire  _GEN_1116 = _GEN_2178 & way2[0] ? valid_41_1 : _GEN_1115; // @[cache.scala 154:{26,26}]
  wire  _GEN_1117 = _GEN_2181 & _GEN_2059 ? valid_42_0 : _GEN_1116; // @[cache.scala 154:{26,26}]
  wire  _GEN_1118 = _GEN_2181 & way2[0] ? valid_42_1 : _GEN_1117; // @[cache.scala 154:{26,26}]
  wire  _GEN_1119 = _GEN_2184 & _GEN_2059 ? valid_43_0 : _GEN_1118; // @[cache.scala 154:{26,26}]
  wire  _GEN_1120 = _GEN_2184 & way2[0] ? valid_43_1 : _GEN_1119; // @[cache.scala 154:{26,26}]
  wire  _GEN_1121 = _GEN_2187 & _GEN_2059 ? valid_44_0 : _GEN_1120; // @[cache.scala 154:{26,26}]
  wire  _GEN_1122 = _GEN_2187 & way2[0] ? valid_44_1 : _GEN_1121; // @[cache.scala 154:{26,26}]
  wire  _GEN_1123 = _GEN_2190 & _GEN_2059 ? valid_45_0 : _GEN_1122; // @[cache.scala 154:{26,26}]
  wire  _GEN_1124 = _GEN_2190 & way2[0] ? valid_45_1 : _GEN_1123; // @[cache.scala 154:{26,26}]
  wire  _GEN_1125 = _GEN_2193 & _GEN_2059 ? valid_46_0 : _GEN_1124; // @[cache.scala 154:{26,26}]
  wire  _GEN_1126 = _GEN_2193 & way2[0] ? valid_46_1 : _GEN_1125; // @[cache.scala 154:{26,26}]
  wire  _GEN_1127 = _GEN_2196 & _GEN_2059 ? valid_47_0 : _GEN_1126; // @[cache.scala 154:{26,26}]
  wire  _GEN_1128 = _GEN_2196 & way2[0] ? valid_47_1 : _GEN_1127; // @[cache.scala 154:{26,26}]
  wire  _GEN_1129 = _GEN_2199 & _GEN_2059 ? valid_48_0 : _GEN_1128; // @[cache.scala 154:{26,26}]
  wire  _GEN_1130 = _GEN_2199 & way2[0] ? valid_48_1 : _GEN_1129; // @[cache.scala 154:{26,26}]
  wire  _GEN_1131 = _GEN_2202 & _GEN_2059 ? valid_49_0 : _GEN_1130; // @[cache.scala 154:{26,26}]
  wire  _GEN_1132 = _GEN_2202 & way2[0] ? valid_49_1 : _GEN_1131; // @[cache.scala 154:{26,26}]
  wire  _GEN_1133 = _GEN_2205 & _GEN_2059 ? valid_50_0 : _GEN_1132; // @[cache.scala 154:{26,26}]
  wire  _GEN_1134 = _GEN_2205 & way2[0] ? valid_50_1 : _GEN_1133; // @[cache.scala 154:{26,26}]
  wire  _GEN_1135 = _GEN_2208 & _GEN_2059 ? valid_51_0 : _GEN_1134; // @[cache.scala 154:{26,26}]
  wire  _GEN_1136 = _GEN_2208 & way2[0] ? valid_51_1 : _GEN_1135; // @[cache.scala 154:{26,26}]
  wire  _GEN_1137 = _GEN_2211 & _GEN_2059 ? valid_52_0 : _GEN_1136; // @[cache.scala 154:{26,26}]
  wire  _GEN_1138 = _GEN_2211 & way2[0] ? valid_52_1 : _GEN_1137; // @[cache.scala 154:{26,26}]
  wire  _GEN_1139 = _GEN_2214 & _GEN_2059 ? valid_53_0 : _GEN_1138; // @[cache.scala 154:{26,26}]
  wire  _GEN_1140 = _GEN_2214 & way2[0] ? valid_53_1 : _GEN_1139; // @[cache.scala 154:{26,26}]
  wire  _GEN_1141 = _GEN_2217 & _GEN_2059 ? valid_54_0 : _GEN_1140; // @[cache.scala 154:{26,26}]
  wire  _GEN_1142 = _GEN_2217 & way2[0] ? valid_54_1 : _GEN_1141; // @[cache.scala 154:{26,26}]
  wire  _GEN_1143 = _GEN_2220 & _GEN_2059 ? valid_55_0 : _GEN_1142; // @[cache.scala 154:{26,26}]
  wire  _GEN_1144 = _GEN_2220 & way2[0] ? valid_55_1 : _GEN_1143; // @[cache.scala 154:{26,26}]
  wire  _GEN_1145 = _GEN_2223 & _GEN_2059 ? valid_56_0 : _GEN_1144; // @[cache.scala 154:{26,26}]
  wire  _GEN_1146 = _GEN_2223 & way2[0] ? valid_56_1 : _GEN_1145; // @[cache.scala 154:{26,26}]
  wire  _GEN_1147 = _GEN_2226 & _GEN_2059 ? valid_57_0 : _GEN_1146; // @[cache.scala 154:{26,26}]
  wire  _GEN_1148 = _GEN_2226 & way2[0] ? valid_57_1 : _GEN_1147; // @[cache.scala 154:{26,26}]
  wire  _GEN_1149 = _GEN_2229 & _GEN_2059 ? valid_58_0 : _GEN_1148; // @[cache.scala 154:{26,26}]
  wire  _GEN_1150 = _GEN_2229 & way2[0] ? valid_58_1 : _GEN_1149; // @[cache.scala 154:{26,26}]
  wire  _GEN_1151 = _GEN_2232 & _GEN_2059 ? valid_59_0 : _GEN_1150; // @[cache.scala 154:{26,26}]
  wire  _GEN_1152 = _GEN_2232 & way2[0] ? valid_59_1 : _GEN_1151; // @[cache.scala 154:{26,26}]
  wire  _GEN_1153 = _GEN_2235 & _GEN_2059 ? valid_60_0 : _GEN_1152; // @[cache.scala 154:{26,26}]
  wire  _GEN_1154 = _GEN_2235 & way2[0] ? valid_60_1 : _GEN_1153; // @[cache.scala 154:{26,26}]
  wire  _GEN_1155 = _GEN_2238 & _GEN_2059 ? valid_61_0 : _GEN_1154; // @[cache.scala 154:{26,26}]
  wire  _GEN_1156 = _GEN_2238 & way2[0] ? valid_61_1 : _GEN_1155; // @[cache.scala 154:{26,26}]
  wire  _GEN_1157 = _GEN_2241 & _GEN_2059 ? valid_62_0 : _GEN_1156; // @[cache.scala 154:{26,26}]
  wire  _GEN_1158 = _GEN_2241 & way2[0] ? valid_62_1 : _GEN_1157; // @[cache.scala 154:{26,26}]
  wire  _GEN_1159 = _GEN_2244 & _GEN_2059 ? valid_63_0 : _GEN_1158; // @[cache.scala 154:{26,26}]
  wire  _GEN_1160 = _GEN_2244 & way2[0] ? valid_63_1 : _GEN_1159; // @[cache.scala 154:{26,26}]
  wire  _GEN_1161 = _GEN_2247 & _GEN_2059 ? valid_64_0 : _GEN_1160; // @[cache.scala 154:{26,26}]
  wire  _GEN_1162 = _GEN_2247 & way2[0] ? valid_64_1 : _GEN_1161; // @[cache.scala 154:{26,26}]
  wire  _GEN_1163 = _GEN_2250 & _GEN_2059 ? valid_65_0 : _GEN_1162; // @[cache.scala 154:{26,26}]
  wire  _GEN_1164 = _GEN_2250 & way2[0] ? valid_65_1 : _GEN_1163; // @[cache.scala 154:{26,26}]
  wire  _GEN_1165 = _GEN_2253 & _GEN_2059 ? valid_66_0 : _GEN_1164; // @[cache.scala 154:{26,26}]
  wire  _GEN_1166 = _GEN_2253 & way2[0] ? valid_66_1 : _GEN_1165; // @[cache.scala 154:{26,26}]
  wire  _GEN_1167 = _GEN_2256 & _GEN_2059 ? valid_67_0 : _GEN_1166; // @[cache.scala 154:{26,26}]
  wire  _GEN_1168 = _GEN_2256 & way2[0] ? valid_67_1 : _GEN_1167; // @[cache.scala 154:{26,26}]
  wire  _GEN_1169 = _GEN_2259 & _GEN_2059 ? valid_68_0 : _GEN_1168; // @[cache.scala 154:{26,26}]
  wire  _GEN_1170 = _GEN_2259 & way2[0] ? valid_68_1 : _GEN_1169; // @[cache.scala 154:{26,26}]
  wire  _GEN_1171 = _GEN_2262 & _GEN_2059 ? valid_69_0 : _GEN_1170; // @[cache.scala 154:{26,26}]
  wire  _GEN_1172 = _GEN_2262 & way2[0] ? valid_69_1 : _GEN_1171; // @[cache.scala 154:{26,26}]
  wire  _GEN_1173 = _GEN_2265 & _GEN_2059 ? valid_70_0 : _GEN_1172; // @[cache.scala 154:{26,26}]
  wire  _GEN_1174 = _GEN_2265 & way2[0] ? valid_70_1 : _GEN_1173; // @[cache.scala 154:{26,26}]
  wire  _GEN_1175 = _GEN_2268 & _GEN_2059 ? valid_71_0 : _GEN_1174; // @[cache.scala 154:{26,26}]
  wire  _GEN_1176 = _GEN_2268 & way2[0] ? valid_71_1 : _GEN_1175; // @[cache.scala 154:{26,26}]
  wire  _GEN_1177 = _GEN_2271 & _GEN_2059 ? valid_72_0 : _GEN_1176; // @[cache.scala 154:{26,26}]
  wire  _GEN_1178 = _GEN_2271 & way2[0] ? valid_72_1 : _GEN_1177; // @[cache.scala 154:{26,26}]
  wire  _GEN_1179 = _GEN_2274 & _GEN_2059 ? valid_73_0 : _GEN_1178; // @[cache.scala 154:{26,26}]
  wire  _GEN_1180 = _GEN_2274 & way2[0] ? valid_73_1 : _GEN_1179; // @[cache.scala 154:{26,26}]
  wire  _GEN_1181 = _GEN_2277 & _GEN_2059 ? valid_74_0 : _GEN_1180; // @[cache.scala 154:{26,26}]
  wire  _GEN_1182 = _GEN_2277 & way2[0] ? valid_74_1 : _GEN_1181; // @[cache.scala 154:{26,26}]
  wire  _GEN_1183 = _GEN_2280 & _GEN_2059 ? valid_75_0 : _GEN_1182; // @[cache.scala 154:{26,26}]
  wire  _GEN_1184 = _GEN_2280 & way2[0] ? valid_75_1 : _GEN_1183; // @[cache.scala 154:{26,26}]
  wire  _GEN_1185 = _GEN_2283 & _GEN_2059 ? valid_76_0 : _GEN_1184; // @[cache.scala 154:{26,26}]
  wire  _GEN_1186 = _GEN_2283 & way2[0] ? valid_76_1 : _GEN_1185; // @[cache.scala 154:{26,26}]
  wire  _GEN_1187 = _GEN_2286 & _GEN_2059 ? valid_77_0 : _GEN_1186; // @[cache.scala 154:{26,26}]
  wire  _GEN_1188 = _GEN_2286 & way2[0] ? valid_77_1 : _GEN_1187; // @[cache.scala 154:{26,26}]
  wire  _GEN_1189 = _GEN_2289 & _GEN_2059 ? valid_78_0 : _GEN_1188; // @[cache.scala 154:{26,26}]
  wire  _GEN_1190 = _GEN_2289 & way2[0] ? valid_78_1 : _GEN_1189; // @[cache.scala 154:{26,26}]
  wire  _GEN_1191 = _GEN_2292 & _GEN_2059 ? valid_79_0 : _GEN_1190; // @[cache.scala 154:{26,26}]
  wire  _GEN_1192 = _GEN_2292 & way2[0] ? valid_79_1 : _GEN_1191; // @[cache.scala 154:{26,26}]
  wire  _GEN_1193 = _GEN_2295 & _GEN_2059 ? valid_80_0 : _GEN_1192; // @[cache.scala 154:{26,26}]
  wire  _GEN_1194 = _GEN_2295 & way2[0] ? valid_80_1 : _GEN_1193; // @[cache.scala 154:{26,26}]
  wire  _GEN_1195 = _GEN_2298 & _GEN_2059 ? valid_81_0 : _GEN_1194; // @[cache.scala 154:{26,26}]
  wire  _GEN_1196 = _GEN_2298 & way2[0] ? valid_81_1 : _GEN_1195; // @[cache.scala 154:{26,26}]
  wire  _GEN_1197 = _GEN_2301 & _GEN_2059 ? valid_82_0 : _GEN_1196; // @[cache.scala 154:{26,26}]
  wire  _GEN_1198 = _GEN_2301 & way2[0] ? valid_82_1 : _GEN_1197; // @[cache.scala 154:{26,26}]
  wire  _GEN_1199 = _GEN_2304 & _GEN_2059 ? valid_83_0 : _GEN_1198; // @[cache.scala 154:{26,26}]
  wire  _GEN_1200 = _GEN_2304 & way2[0] ? valid_83_1 : _GEN_1199; // @[cache.scala 154:{26,26}]
  wire  _GEN_1201 = _GEN_2307 & _GEN_2059 ? valid_84_0 : _GEN_1200; // @[cache.scala 154:{26,26}]
  wire  _GEN_1202 = _GEN_2307 & way2[0] ? valid_84_1 : _GEN_1201; // @[cache.scala 154:{26,26}]
  wire  _GEN_1203 = _GEN_2310 & _GEN_2059 ? valid_85_0 : _GEN_1202; // @[cache.scala 154:{26,26}]
  wire  _GEN_1204 = _GEN_2310 & way2[0] ? valid_85_1 : _GEN_1203; // @[cache.scala 154:{26,26}]
  wire  _GEN_1205 = _GEN_2313 & _GEN_2059 ? valid_86_0 : _GEN_1204; // @[cache.scala 154:{26,26}]
  wire  _GEN_1206 = _GEN_2313 & way2[0] ? valid_86_1 : _GEN_1205; // @[cache.scala 154:{26,26}]
  wire  _GEN_1207 = _GEN_2316 & _GEN_2059 ? valid_87_0 : _GEN_1206; // @[cache.scala 154:{26,26}]
  wire  _GEN_1208 = _GEN_2316 & way2[0] ? valid_87_1 : _GEN_1207; // @[cache.scala 154:{26,26}]
  wire  _GEN_1209 = _GEN_2319 & _GEN_2059 ? valid_88_0 : _GEN_1208; // @[cache.scala 154:{26,26}]
  wire  _GEN_1210 = _GEN_2319 & way2[0] ? valid_88_1 : _GEN_1209; // @[cache.scala 154:{26,26}]
  wire  _GEN_1211 = _GEN_2322 & _GEN_2059 ? valid_89_0 : _GEN_1210; // @[cache.scala 154:{26,26}]
  wire  _GEN_1212 = _GEN_2322 & way2[0] ? valid_89_1 : _GEN_1211; // @[cache.scala 154:{26,26}]
  wire  _GEN_1213 = _GEN_2325 & _GEN_2059 ? valid_90_0 : _GEN_1212; // @[cache.scala 154:{26,26}]
  wire  _GEN_1214 = _GEN_2325 & way2[0] ? valid_90_1 : _GEN_1213; // @[cache.scala 154:{26,26}]
  wire  _GEN_1215 = _GEN_2328 & _GEN_2059 ? valid_91_0 : _GEN_1214; // @[cache.scala 154:{26,26}]
  wire  _GEN_1216 = _GEN_2328 & way2[0] ? valid_91_1 : _GEN_1215; // @[cache.scala 154:{26,26}]
  wire  _GEN_1217 = _GEN_2331 & _GEN_2059 ? valid_92_0 : _GEN_1216; // @[cache.scala 154:{26,26}]
  wire  _GEN_1218 = _GEN_2331 & way2[0] ? valid_92_1 : _GEN_1217; // @[cache.scala 154:{26,26}]
  wire  _GEN_1219 = _GEN_2334 & _GEN_2059 ? valid_93_0 : _GEN_1218; // @[cache.scala 154:{26,26}]
  wire  _GEN_1220 = _GEN_2334 & way2[0] ? valid_93_1 : _GEN_1219; // @[cache.scala 154:{26,26}]
  wire  _GEN_1221 = _GEN_2337 & _GEN_2059 ? valid_94_0 : _GEN_1220; // @[cache.scala 154:{26,26}]
  wire  _GEN_1222 = _GEN_2337 & way2[0] ? valid_94_1 : _GEN_1221; // @[cache.scala 154:{26,26}]
  wire  _GEN_1223 = _GEN_2340 & _GEN_2059 ? valid_95_0 : _GEN_1222; // @[cache.scala 154:{26,26}]
  wire  _GEN_1224 = _GEN_2340 & way2[0] ? valid_95_1 : _GEN_1223; // @[cache.scala 154:{26,26}]
  wire  _GEN_1225 = _GEN_2343 & _GEN_2059 ? valid_96_0 : _GEN_1224; // @[cache.scala 154:{26,26}]
  wire  _GEN_1226 = _GEN_2343 & way2[0] ? valid_96_1 : _GEN_1225; // @[cache.scala 154:{26,26}]
  wire  _GEN_1227 = _GEN_2346 & _GEN_2059 ? valid_97_0 : _GEN_1226; // @[cache.scala 154:{26,26}]
  wire  _GEN_1228 = _GEN_2346 & way2[0] ? valid_97_1 : _GEN_1227; // @[cache.scala 154:{26,26}]
  wire  _GEN_1229 = _GEN_2349 & _GEN_2059 ? valid_98_0 : _GEN_1228; // @[cache.scala 154:{26,26}]
  wire  _GEN_1230 = _GEN_2349 & way2[0] ? valid_98_1 : _GEN_1229; // @[cache.scala 154:{26,26}]
  wire  _GEN_1231 = _GEN_2352 & _GEN_2059 ? valid_99_0 : _GEN_1230; // @[cache.scala 154:{26,26}]
  wire  _GEN_1232 = _GEN_2352 & way2[0] ? valid_99_1 : _GEN_1231; // @[cache.scala 154:{26,26}]
  wire  _GEN_1233 = _GEN_2355 & _GEN_2059 ? valid_100_0 : _GEN_1232; // @[cache.scala 154:{26,26}]
  wire  _GEN_1234 = _GEN_2355 & way2[0] ? valid_100_1 : _GEN_1233; // @[cache.scala 154:{26,26}]
  wire  _GEN_1235 = _GEN_2358 & _GEN_2059 ? valid_101_0 : _GEN_1234; // @[cache.scala 154:{26,26}]
  wire  _GEN_1236 = _GEN_2358 & way2[0] ? valid_101_1 : _GEN_1235; // @[cache.scala 154:{26,26}]
  wire  _GEN_1237 = _GEN_2361 & _GEN_2059 ? valid_102_0 : _GEN_1236; // @[cache.scala 154:{26,26}]
  wire  _GEN_1238 = _GEN_2361 & way2[0] ? valid_102_1 : _GEN_1237; // @[cache.scala 154:{26,26}]
  wire  _GEN_1239 = _GEN_2364 & _GEN_2059 ? valid_103_0 : _GEN_1238; // @[cache.scala 154:{26,26}]
  wire  _GEN_1240 = _GEN_2364 & way2[0] ? valid_103_1 : _GEN_1239; // @[cache.scala 154:{26,26}]
  wire  _GEN_1241 = _GEN_2367 & _GEN_2059 ? valid_104_0 : _GEN_1240; // @[cache.scala 154:{26,26}]
  wire  _GEN_1242 = _GEN_2367 & way2[0] ? valid_104_1 : _GEN_1241; // @[cache.scala 154:{26,26}]
  wire  _GEN_1243 = _GEN_2370 & _GEN_2059 ? valid_105_0 : _GEN_1242; // @[cache.scala 154:{26,26}]
  wire  _GEN_1244 = _GEN_2370 & way2[0] ? valid_105_1 : _GEN_1243; // @[cache.scala 154:{26,26}]
  wire  _GEN_1245 = _GEN_2373 & _GEN_2059 ? valid_106_0 : _GEN_1244; // @[cache.scala 154:{26,26}]
  wire  _GEN_1246 = _GEN_2373 & way2[0] ? valid_106_1 : _GEN_1245; // @[cache.scala 154:{26,26}]
  wire  _GEN_1247 = _GEN_2376 & _GEN_2059 ? valid_107_0 : _GEN_1246; // @[cache.scala 154:{26,26}]
  wire  _GEN_1248 = _GEN_2376 & way2[0] ? valid_107_1 : _GEN_1247; // @[cache.scala 154:{26,26}]
  wire  _GEN_1249 = _GEN_2379 & _GEN_2059 ? valid_108_0 : _GEN_1248; // @[cache.scala 154:{26,26}]
  wire  _GEN_1250 = _GEN_2379 & way2[0] ? valid_108_1 : _GEN_1249; // @[cache.scala 154:{26,26}]
  wire  _GEN_1251 = _GEN_2382 & _GEN_2059 ? valid_109_0 : _GEN_1250; // @[cache.scala 154:{26,26}]
  wire  _GEN_1252 = _GEN_2382 & way2[0] ? valid_109_1 : _GEN_1251; // @[cache.scala 154:{26,26}]
  wire  _GEN_1253 = _GEN_2385 & _GEN_2059 ? valid_110_0 : _GEN_1252; // @[cache.scala 154:{26,26}]
  wire  _GEN_1254 = _GEN_2385 & way2[0] ? valid_110_1 : _GEN_1253; // @[cache.scala 154:{26,26}]
  wire  _GEN_1255 = _GEN_2388 & _GEN_2059 ? valid_111_0 : _GEN_1254; // @[cache.scala 154:{26,26}]
  wire  _GEN_1256 = _GEN_2388 & way2[0] ? valid_111_1 : _GEN_1255; // @[cache.scala 154:{26,26}]
  wire  _GEN_1257 = _GEN_2391 & _GEN_2059 ? valid_112_0 : _GEN_1256; // @[cache.scala 154:{26,26}]
  wire  _GEN_1258 = _GEN_2391 & way2[0] ? valid_112_1 : _GEN_1257; // @[cache.scala 154:{26,26}]
  wire  _GEN_1259 = _GEN_2394 & _GEN_2059 ? valid_113_0 : _GEN_1258; // @[cache.scala 154:{26,26}]
  wire  _GEN_1260 = _GEN_2394 & way2[0] ? valid_113_1 : _GEN_1259; // @[cache.scala 154:{26,26}]
  wire  _GEN_1261 = _GEN_2397 & _GEN_2059 ? valid_114_0 : _GEN_1260; // @[cache.scala 154:{26,26}]
  wire  _GEN_1262 = _GEN_2397 & way2[0] ? valid_114_1 : _GEN_1261; // @[cache.scala 154:{26,26}]
  wire  _GEN_1263 = _GEN_2400 & _GEN_2059 ? valid_115_0 : _GEN_1262; // @[cache.scala 154:{26,26}]
  wire  _GEN_1264 = _GEN_2400 & way2[0] ? valid_115_1 : _GEN_1263; // @[cache.scala 154:{26,26}]
  wire  _GEN_1265 = _GEN_2403 & _GEN_2059 ? valid_116_0 : _GEN_1264; // @[cache.scala 154:{26,26}]
  wire  _GEN_1266 = _GEN_2403 & way2[0] ? valid_116_1 : _GEN_1265; // @[cache.scala 154:{26,26}]
  wire  _GEN_1267 = _GEN_2406 & _GEN_2059 ? valid_117_0 : _GEN_1266; // @[cache.scala 154:{26,26}]
  wire  _GEN_1268 = _GEN_2406 & way2[0] ? valid_117_1 : _GEN_1267; // @[cache.scala 154:{26,26}]
  wire  _GEN_1269 = _GEN_2409 & _GEN_2059 ? valid_118_0 : _GEN_1268; // @[cache.scala 154:{26,26}]
  wire  _GEN_1270 = _GEN_2409 & way2[0] ? valid_118_1 : _GEN_1269; // @[cache.scala 154:{26,26}]
  wire  _GEN_1271 = _GEN_2412 & _GEN_2059 ? valid_119_0 : _GEN_1270; // @[cache.scala 154:{26,26}]
  wire  _GEN_1272 = _GEN_2412 & way2[0] ? valid_119_1 : _GEN_1271; // @[cache.scala 154:{26,26}]
  wire  _GEN_1273 = _GEN_2415 & _GEN_2059 ? valid_120_0 : _GEN_1272; // @[cache.scala 154:{26,26}]
  wire  _GEN_1274 = _GEN_2415 & way2[0] ? valid_120_1 : _GEN_1273; // @[cache.scala 154:{26,26}]
  wire  _GEN_1275 = _GEN_2418 & _GEN_2059 ? valid_121_0 : _GEN_1274; // @[cache.scala 154:{26,26}]
  wire  _GEN_1276 = _GEN_2418 & way2[0] ? valid_121_1 : _GEN_1275; // @[cache.scala 154:{26,26}]
  wire  _GEN_1277 = _GEN_2421 & _GEN_2059 ? valid_122_0 : _GEN_1276; // @[cache.scala 154:{26,26}]
  wire  _GEN_1278 = _GEN_2421 & way2[0] ? valid_122_1 : _GEN_1277; // @[cache.scala 154:{26,26}]
  wire  _GEN_1279 = _GEN_2424 & _GEN_2059 ? valid_123_0 : _GEN_1278; // @[cache.scala 154:{26,26}]
  wire  _GEN_1280 = _GEN_2424 & way2[0] ? valid_123_1 : _GEN_1279; // @[cache.scala 154:{26,26}]
  wire  _GEN_1281 = _GEN_2427 & _GEN_2059 ? valid_124_0 : _GEN_1280; // @[cache.scala 154:{26,26}]
  wire  _GEN_1282 = _GEN_2427 & way2[0] ? valid_124_1 : _GEN_1281; // @[cache.scala 154:{26,26}]
  wire  _GEN_1283 = _GEN_2430 & _GEN_2059 ? valid_125_0 : _GEN_1282; // @[cache.scala 154:{26,26}]
  wire  _GEN_1284 = _GEN_2430 & way2[0] ? valid_125_1 : _GEN_1283; // @[cache.scala 154:{26,26}]
  wire  _GEN_1285 = _GEN_2433 & _GEN_2059 ? valid_126_0 : _GEN_1284; // @[cache.scala 154:{26,26}]
  wire  _GEN_1286 = _GEN_2433 & way2[0] ? valid_126_1 : _GEN_1285; // @[cache.scala 154:{26,26}]
  wire  _GEN_1287 = _GEN_2436 & _GEN_2059 ? valid_127_0 : _GEN_1286; // @[cache.scala 154:{26,26}]
  wire  _GEN_1288 = _GEN_2436 & way2[0] ? valid_127_1 : _GEN_1287; // @[cache.scala 154:{26,26}]
  wire  _d_way_T_2 = _io_in_r_bits_data_T & wmode; // @[cache.scala 157:33]
  wire [7:0] _d_way_T_4 = _io_in_r_bits_data_T_3 ? way2 : 8'h0; // @[cache.scala 158:16]
  wire [7:0] d_way = _io_in_r_bits_data_T & wmode ? hit_way : _d_way_T_4; // @[cache.scala 157:16]
  wire  _GEN_1546 = _GEN_2057 & d_way[0] ? dirty_0_1 : dirty_0_0; // @[cache.scala 160:{28,28}]
  wire  _GEN_3973 = ~d_way[0]; // @[cache.scala 160:{28,28}]
  wire  _GEN_1547 = _GEN_2058 & ~d_way[0] ? dirty_1_0 : _GEN_1546; // @[cache.scala 160:{28,28}]
  wire  _GEN_1548 = _GEN_2058 & d_way[0] ? dirty_1_1 : _GEN_1547; // @[cache.scala 160:{28,28}]
  wire  _GEN_1549 = _GEN_2061 & ~d_way[0] ? dirty_2_0 : _GEN_1548; // @[cache.scala 160:{28,28}]
  wire  _GEN_1550 = _GEN_2061 & d_way[0] ? dirty_2_1 : _GEN_1549; // @[cache.scala 160:{28,28}]
  wire  _GEN_1551 = _GEN_2064 & ~d_way[0] ? dirty_3_0 : _GEN_1550; // @[cache.scala 160:{28,28}]
  wire  _GEN_1552 = _GEN_2064 & d_way[0] ? dirty_3_1 : _GEN_1551; // @[cache.scala 160:{28,28}]
  wire  _GEN_1553 = _GEN_2067 & ~d_way[0] ? dirty_4_0 : _GEN_1552; // @[cache.scala 160:{28,28}]
  wire  _GEN_1554 = _GEN_2067 & d_way[0] ? dirty_4_1 : _GEN_1553; // @[cache.scala 160:{28,28}]
  wire  _GEN_1555 = _GEN_2070 & ~d_way[0] ? dirty_5_0 : _GEN_1554; // @[cache.scala 160:{28,28}]
  wire  _GEN_1556 = _GEN_2070 & d_way[0] ? dirty_5_1 : _GEN_1555; // @[cache.scala 160:{28,28}]
  wire  _GEN_1557 = _GEN_2073 & ~d_way[0] ? dirty_6_0 : _GEN_1556; // @[cache.scala 160:{28,28}]
  wire  _GEN_1558 = _GEN_2073 & d_way[0] ? dirty_6_1 : _GEN_1557; // @[cache.scala 160:{28,28}]
  wire  _GEN_1559 = _GEN_2076 & ~d_way[0] ? dirty_7_0 : _GEN_1558; // @[cache.scala 160:{28,28}]
  wire  _GEN_1560 = _GEN_2076 & d_way[0] ? dirty_7_1 : _GEN_1559; // @[cache.scala 160:{28,28}]
  wire  _GEN_1561 = _GEN_2079 & ~d_way[0] ? dirty_8_0 : _GEN_1560; // @[cache.scala 160:{28,28}]
  wire  _GEN_1562 = _GEN_2079 & d_way[0] ? dirty_8_1 : _GEN_1561; // @[cache.scala 160:{28,28}]
  wire  _GEN_1563 = _GEN_2082 & ~d_way[0] ? dirty_9_0 : _GEN_1562; // @[cache.scala 160:{28,28}]
  wire  _GEN_1564 = _GEN_2082 & d_way[0] ? dirty_9_1 : _GEN_1563; // @[cache.scala 160:{28,28}]
  wire  _GEN_1565 = _GEN_2085 & ~d_way[0] ? dirty_10_0 : _GEN_1564; // @[cache.scala 160:{28,28}]
  wire  _GEN_1566 = _GEN_2085 & d_way[0] ? dirty_10_1 : _GEN_1565; // @[cache.scala 160:{28,28}]
  wire  _GEN_1567 = _GEN_2088 & ~d_way[0] ? dirty_11_0 : _GEN_1566; // @[cache.scala 160:{28,28}]
  wire  _GEN_1568 = _GEN_2088 & d_way[0] ? dirty_11_1 : _GEN_1567; // @[cache.scala 160:{28,28}]
  wire  _GEN_1569 = _GEN_2091 & ~d_way[0] ? dirty_12_0 : _GEN_1568; // @[cache.scala 160:{28,28}]
  wire  _GEN_1570 = _GEN_2091 & d_way[0] ? dirty_12_1 : _GEN_1569; // @[cache.scala 160:{28,28}]
  wire  _GEN_1571 = _GEN_2094 & ~d_way[0] ? dirty_13_0 : _GEN_1570; // @[cache.scala 160:{28,28}]
  wire  _GEN_1572 = _GEN_2094 & d_way[0] ? dirty_13_1 : _GEN_1571; // @[cache.scala 160:{28,28}]
  wire  _GEN_1573 = _GEN_2097 & ~d_way[0] ? dirty_14_0 : _GEN_1572; // @[cache.scala 160:{28,28}]
  wire  _GEN_1574 = _GEN_2097 & d_way[0] ? dirty_14_1 : _GEN_1573; // @[cache.scala 160:{28,28}]
  wire  _GEN_1575 = _GEN_2100 & ~d_way[0] ? dirty_15_0 : _GEN_1574; // @[cache.scala 160:{28,28}]
  wire  _GEN_1576 = _GEN_2100 & d_way[0] ? dirty_15_1 : _GEN_1575; // @[cache.scala 160:{28,28}]
  wire  _GEN_1577 = _GEN_2103 & ~d_way[0] ? dirty_16_0 : _GEN_1576; // @[cache.scala 160:{28,28}]
  wire  _GEN_1578 = _GEN_2103 & d_way[0] ? dirty_16_1 : _GEN_1577; // @[cache.scala 160:{28,28}]
  wire  _GEN_1579 = _GEN_2106 & ~d_way[0] ? dirty_17_0 : _GEN_1578; // @[cache.scala 160:{28,28}]
  wire  _GEN_1580 = _GEN_2106 & d_way[0] ? dirty_17_1 : _GEN_1579; // @[cache.scala 160:{28,28}]
  wire  _GEN_1581 = _GEN_2109 & ~d_way[0] ? dirty_18_0 : _GEN_1580; // @[cache.scala 160:{28,28}]
  wire  _GEN_1582 = _GEN_2109 & d_way[0] ? dirty_18_1 : _GEN_1581; // @[cache.scala 160:{28,28}]
  wire  _GEN_1583 = _GEN_2112 & ~d_way[0] ? dirty_19_0 : _GEN_1582; // @[cache.scala 160:{28,28}]
  wire  _GEN_1584 = _GEN_2112 & d_way[0] ? dirty_19_1 : _GEN_1583; // @[cache.scala 160:{28,28}]
  wire  _GEN_1585 = _GEN_2115 & ~d_way[0] ? dirty_20_0 : _GEN_1584; // @[cache.scala 160:{28,28}]
  wire  _GEN_1586 = _GEN_2115 & d_way[0] ? dirty_20_1 : _GEN_1585; // @[cache.scala 160:{28,28}]
  wire  _GEN_1587 = _GEN_2118 & ~d_way[0] ? dirty_21_0 : _GEN_1586; // @[cache.scala 160:{28,28}]
  wire  _GEN_1588 = _GEN_2118 & d_way[0] ? dirty_21_1 : _GEN_1587; // @[cache.scala 160:{28,28}]
  wire  _GEN_1589 = _GEN_2121 & ~d_way[0] ? dirty_22_0 : _GEN_1588; // @[cache.scala 160:{28,28}]
  wire  _GEN_1590 = _GEN_2121 & d_way[0] ? dirty_22_1 : _GEN_1589; // @[cache.scala 160:{28,28}]
  wire  _GEN_1591 = _GEN_2124 & ~d_way[0] ? dirty_23_0 : _GEN_1590; // @[cache.scala 160:{28,28}]
  wire  _GEN_1592 = _GEN_2124 & d_way[0] ? dirty_23_1 : _GEN_1591; // @[cache.scala 160:{28,28}]
  wire  _GEN_1593 = _GEN_2127 & ~d_way[0] ? dirty_24_0 : _GEN_1592; // @[cache.scala 160:{28,28}]
  wire  _GEN_1594 = _GEN_2127 & d_way[0] ? dirty_24_1 : _GEN_1593; // @[cache.scala 160:{28,28}]
  wire  _GEN_1595 = _GEN_2130 & ~d_way[0] ? dirty_25_0 : _GEN_1594; // @[cache.scala 160:{28,28}]
  wire  _GEN_1596 = _GEN_2130 & d_way[0] ? dirty_25_1 : _GEN_1595; // @[cache.scala 160:{28,28}]
  wire  _GEN_1597 = _GEN_2133 & ~d_way[0] ? dirty_26_0 : _GEN_1596; // @[cache.scala 160:{28,28}]
  wire  _GEN_1598 = _GEN_2133 & d_way[0] ? dirty_26_1 : _GEN_1597; // @[cache.scala 160:{28,28}]
  wire  _GEN_1599 = _GEN_2136 & ~d_way[0] ? dirty_27_0 : _GEN_1598; // @[cache.scala 160:{28,28}]
  wire  _GEN_1600 = _GEN_2136 & d_way[0] ? dirty_27_1 : _GEN_1599; // @[cache.scala 160:{28,28}]
  wire  _GEN_1601 = _GEN_2139 & ~d_way[0] ? dirty_28_0 : _GEN_1600; // @[cache.scala 160:{28,28}]
  wire  _GEN_1602 = _GEN_2139 & d_way[0] ? dirty_28_1 : _GEN_1601; // @[cache.scala 160:{28,28}]
  wire  _GEN_1603 = _GEN_2142 & ~d_way[0] ? dirty_29_0 : _GEN_1602; // @[cache.scala 160:{28,28}]
  wire  _GEN_1604 = _GEN_2142 & d_way[0] ? dirty_29_1 : _GEN_1603; // @[cache.scala 160:{28,28}]
  wire  _GEN_1605 = _GEN_2145 & ~d_way[0] ? dirty_30_0 : _GEN_1604; // @[cache.scala 160:{28,28}]
  wire  _GEN_1606 = _GEN_2145 & d_way[0] ? dirty_30_1 : _GEN_1605; // @[cache.scala 160:{28,28}]
  wire  _GEN_1607 = _GEN_2148 & ~d_way[0] ? dirty_31_0 : _GEN_1606; // @[cache.scala 160:{28,28}]
  wire  _GEN_1608 = _GEN_2148 & d_way[0] ? dirty_31_1 : _GEN_1607; // @[cache.scala 160:{28,28}]
  wire  _GEN_1609 = _GEN_2151 & ~d_way[0] ? dirty_32_0 : _GEN_1608; // @[cache.scala 160:{28,28}]
  wire  _GEN_1610 = _GEN_2151 & d_way[0] ? dirty_32_1 : _GEN_1609; // @[cache.scala 160:{28,28}]
  wire  _GEN_1611 = _GEN_2154 & ~d_way[0] ? dirty_33_0 : _GEN_1610; // @[cache.scala 160:{28,28}]
  wire  _GEN_1612 = _GEN_2154 & d_way[0] ? dirty_33_1 : _GEN_1611; // @[cache.scala 160:{28,28}]
  wire  _GEN_1613 = _GEN_2157 & ~d_way[0] ? dirty_34_0 : _GEN_1612; // @[cache.scala 160:{28,28}]
  wire  _GEN_1614 = _GEN_2157 & d_way[0] ? dirty_34_1 : _GEN_1613; // @[cache.scala 160:{28,28}]
  wire  _GEN_1615 = _GEN_2160 & ~d_way[0] ? dirty_35_0 : _GEN_1614; // @[cache.scala 160:{28,28}]
  wire  _GEN_1616 = _GEN_2160 & d_way[0] ? dirty_35_1 : _GEN_1615; // @[cache.scala 160:{28,28}]
  wire  _GEN_1617 = _GEN_2163 & ~d_way[0] ? dirty_36_0 : _GEN_1616; // @[cache.scala 160:{28,28}]
  wire  _GEN_1618 = _GEN_2163 & d_way[0] ? dirty_36_1 : _GEN_1617; // @[cache.scala 160:{28,28}]
  wire  _GEN_1619 = _GEN_2166 & ~d_way[0] ? dirty_37_0 : _GEN_1618; // @[cache.scala 160:{28,28}]
  wire  _GEN_1620 = _GEN_2166 & d_way[0] ? dirty_37_1 : _GEN_1619; // @[cache.scala 160:{28,28}]
  wire  _GEN_1621 = _GEN_2169 & ~d_way[0] ? dirty_38_0 : _GEN_1620; // @[cache.scala 160:{28,28}]
  wire  _GEN_1622 = _GEN_2169 & d_way[0] ? dirty_38_1 : _GEN_1621; // @[cache.scala 160:{28,28}]
  wire  _GEN_1623 = _GEN_2172 & ~d_way[0] ? dirty_39_0 : _GEN_1622; // @[cache.scala 160:{28,28}]
  wire  _GEN_1624 = _GEN_2172 & d_way[0] ? dirty_39_1 : _GEN_1623; // @[cache.scala 160:{28,28}]
  wire  _GEN_1625 = _GEN_2175 & ~d_way[0] ? dirty_40_0 : _GEN_1624; // @[cache.scala 160:{28,28}]
  wire  _GEN_1626 = _GEN_2175 & d_way[0] ? dirty_40_1 : _GEN_1625; // @[cache.scala 160:{28,28}]
  wire  _GEN_1627 = _GEN_2178 & ~d_way[0] ? dirty_41_0 : _GEN_1626; // @[cache.scala 160:{28,28}]
  wire  _GEN_1628 = _GEN_2178 & d_way[0] ? dirty_41_1 : _GEN_1627; // @[cache.scala 160:{28,28}]
  wire  _GEN_1629 = _GEN_2181 & ~d_way[0] ? dirty_42_0 : _GEN_1628; // @[cache.scala 160:{28,28}]
  wire  _GEN_1630 = _GEN_2181 & d_way[0] ? dirty_42_1 : _GEN_1629; // @[cache.scala 160:{28,28}]
  wire  _GEN_1631 = _GEN_2184 & ~d_way[0] ? dirty_43_0 : _GEN_1630; // @[cache.scala 160:{28,28}]
  wire  _GEN_1632 = _GEN_2184 & d_way[0] ? dirty_43_1 : _GEN_1631; // @[cache.scala 160:{28,28}]
  wire  _GEN_1633 = _GEN_2187 & ~d_way[0] ? dirty_44_0 : _GEN_1632; // @[cache.scala 160:{28,28}]
  wire  _GEN_1634 = _GEN_2187 & d_way[0] ? dirty_44_1 : _GEN_1633; // @[cache.scala 160:{28,28}]
  wire  _GEN_1635 = _GEN_2190 & ~d_way[0] ? dirty_45_0 : _GEN_1634; // @[cache.scala 160:{28,28}]
  wire  _GEN_1636 = _GEN_2190 & d_way[0] ? dirty_45_1 : _GEN_1635; // @[cache.scala 160:{28,28}]
  wire  _GEN_1637 = _GEN_2193 & ~d_way[0] ? dirty_46_0 : _GEN_1636; // @[cache.scala 160:{28,28}]
  wire  _GEN_1638 = _GEN_2193 & d_way[0] ? dirty_46_1 : _GEN_1637; // @[cache.scala 160:{28,28}]
  wire  _GEN_1639 = _GEN_2196 & ~d_way[0] ? dirty_47_0 : _GEN_1638; // @[cache.scala 160:{28,28}]
  wire  _GEN_1640 = _GEN_2196 & d_way[0] ? dirty_47_1 : _GEN_1639; // @[cache.scala 160:{28,28}]
  wire  _GEN_1641 = _GEN_2199 & ~d_way[0] ? dirty_48_0 : _GEN_1640; // @[cache.scala 160:{28,28}]
  wire  _GEN_1642 = _GEN_2199 & d_way[0] ? dirty_48_1 : _GEN_1641; // @[cache.scala 160:{28,28}]
  wire  _GEN_1643 = _GEN_2202 & ~d_way[0] ? dirty_49_0 : _GEN_1642; // @[cache.scala 160:{28,28}]
  wire  _GEN_1644 = _GEN_2202 & d_way[0] ? dirty_49_1 : _GEN_1643; // @[cache.scala 160:{28,28}]
  wire  _GEN_1645 = _GEN_2205 & ~d_way[0] ? dirty_50_0 : _GEN_1644; // @[cache.scala 160:{28,28}]
  wire  _GEN_1646 = _GEN_2205 & d_way[0] ? dirty_50_1 : _GEN_1645; // @[cache.scala 160:{28,28}]
  wire  _GEN_1647 = _GEN_2208 & ~d_way[0] ? dirty_51_0 : _GEN_1646; // @[cache.scala 160:{28,28}]
  wire  _GEN_1648 = _GEN_2208 & d_way[0] ? dirty_51_1 : _GEN_1647; // @[cache.scala 160:{28,28}]
  wire  _GEN_1649 = _GEN_2211 & ~d_way[0] ? dirty_52_0 : _GEN_1648; // @[cache.scala 160:{28,28}]
  wire  _GEN_1650 = _GEN_2211 & d_way[0] ? dirty_52_1 : _GEN_1649; // @[cache.scala 160:{28,28}]
  wire  _GEN_1651 = _GEN_2214 & ~d_way[0] ? dirty_53_0 : _GEN_1650; // @[cache.scala 160:{28,28}]
  wire  _GEN_1652 = _GEN_2214 & d_way[0] ? dirty_53_1 : _GEN_1651; // @[cache.scala 160:{28,28}]
  wire  _GEN_1653 = _GEN_2217 & ~d_way[0] ? dirty_54_0 : _GEN_1652; // @[cache.scala 160:{28,28}]
  wire  _GEN_1654 = _GEN_2217 & d_way[0] ? dirty_54_1 : _GEN_1653; // @[cache.scala 160:{28,28}]
  wire  _GEN_1655 = _GEN_2220 & ~d_way[0] ? dirty_55_0 : _GEN_1654; // @[cache.scala 160:{28,28}]
  wire  _GEN_1656 = _GEN_2220 & d_way[0] ? dirty_55_1 : _GEN_1655; // @[cache.scala 160:{28,28}]
  wire  _GEN_1657 = _GEN_2223 & ~d_way[0] ? dirty_56_0 : _GEN_1656; // @[cache.scala 160:{28,28}]
  wire  _GEN_1658 = _GEN_2223 & d_way[0] ? dirty_56_1 : _GEN_1657; // @[cache.scala 160:{28,28}]
  wire  _GEN_1659 = _GEN_2226 & ~d_way[0] ? dirty_57_0 : _GEN_1658; // @[cache.scala 160:{28,28}]
  wire  _GEN_1660 = _GEN_2226 & d_way[0] ? dirty_57_1 : _GEN_1659; // @[cache.scala 160:{28,28}]
  wire  _GEN_1661 = _GEN_2229 & ~d_way[0] ? dirty_58_0 : _GEN_1660; // @[cache.scala 160:{28,28}]
  wire  _GEN_1662 = _GEN_2229 & d_way[0] ? dirty_58_1 : _GEN_1661; // @[cache.scala 160:{28,28}]
  wire  _GEN_1663 = _GEN_2232 & ~d_way[0] ? dirty_59_0 : _GEN_1662; // @[cache.scala 160:{28,28}]
  wire  _GEN_1664 = _GEN_2232 & d_way[0] ? dirty_59_1 : _GEN_1663; // @[cache.scala 160:{28,28}]
  wire  _GEN_1665 = _GEN_2235 & ~d_way[0] ? dirty_60_0 : _GEN_1664; // @[cache.scala 160:{28,28}]
  wire  _GEN_1666 = _GEN_2235 & d_way[0] ? dirty_60_1 : _GEN_1665; // @[cache.scala 160:{28,28}]
  wire  _GEN_1667 = _GEN_2238 & ~d_way[0] ? dirty_61_0 : _GEN_1666; // @[cache.scala 160:{28,28}]
  wire  _GEN_1668 = _GEN_2238 & d_way[0] ? dirty_61_1 : _GEN_1667; // @[cache.scala 160:{28,28}]
  wire  _GEN_1669 = _GEN_2241 & ~d_way[0] ? dirty_62_0 : _GEN_1668; // @[cache.scala 160:{28,28}]
  wire  _GEN_1670 = _GEN_2241 & d_way[0] ? dirty_62_1 : _GEN_1669; // @[cache.scala 160:{28,28}]
  wire  _GEN_1671 = _GEN_2244 & ~d_way[0] ? dirty_63_0 : _GEN_1670; // @[cache.scala 160:{28,28}]
  wire  _GEN_1672 = _GEN_2244 & d_way[0] ? dirty_63_1 : _GEN_1671; // @[cache.scala 160:{28,28}]
  wire  _GEN_1673 = _GEN_2247 & ~d_way[0] ? dirty_64_0 : _GEN_1672; // @[cache.scala 160:{28,28}]
  wire  _GEN_1674 = _GEN_2247 & d_way[0] ? dirty_64_1 : _GEN_1673; // @[cache.scala 160:{28,28}]
  wire  _GEN_1675 = _GEN_2250 & ~d_way[0] ? dirty_65_0 : _GEN_1674; // @[cache.scala 160:{28,28}]
  wire  _GEN_1676 = _GEN_2250 & d_way[0] ? dirty_65_1 : _GEN_1675; // @[cache.scala 160:{28,28}]
  wire  _GEN_1677 = _GEN_2253 & ~d_way[0] ? dirty_66_0 : _GEN_1676; // @[cache.scala 160:{28,28}]
  wire  _GEN_1678 = _GEN_2253 & d_way[0] ? dirty_66_1 : _GEN_1677; // @[cache.scala 160:{28,28}]
  wire  _GEN_1679 = _GEN_2256 & ~d_way[0] ? dirty_67_0 : _GEN_1678; // @[cache.scala 160:{28,28}]
  wire  _GEN_1680 = _GEN_2256 & d_way[0] ? dirty_67_1 : _GEN_1679; // @[cache.scala 160:{28,28}]
  wire  _GEN_1681 = _GEN_2259 & ~d_way[0] ? dirty_68_0 : _GEN_1680; // @[cache.scala 160:{28,28}]
  wire  _GEN_1682 = _GEN_2259 & d_way[0] ? dirty_68_1 : _GEN_1681; // @[cache.scala 160:{28,28}]
  wire  _GEN_1683 = _GEN_2262 & ~d_way[0] ? dirty_69_0 : _GEN_1682; // @[cache.scala 160:{28,28}]
  wire  _GEN_1684 = _GEN_2262 & d_way[0] ? dirty_69_1 : _GEN_1683; // @[cache.scala 160:{28,28}]
  wire  _GEN_1685 = _GEN_2265 & ~d_way[0] ? dirty_70_0 : _GEN_1684; // @[cache.scala 160:{28,28}]
  wire  _GEN_1686 = _GEN_2265 & d_way[0] ? dirty_70_1 : _GEN_1685; // @[cache.scala 160:{28,28}]
  wire  _GEN_1687 = _GEN_2268 & ~d_way[0] ? dirty_71_0 : _GEN_1686; // @[cache.scala 160:{28,28}]
  wire  _GEN_1688 = _GEN_2268 & d_way[0] ? dirty_71_1 : _GEN_1687; // @[cache.scala 160:{28,28}]
  wire  _GEN_1689 = _GEN_2271 & ~d_way[0] ? dirty_72_0 : _GEN_1688; // @[cache.scala 160:{28,28}]
  wire  _GEN_1690 = _GEN_2271 & d_way[0] ? dirty_72_1 : _GEN_1689; // @[cache.scala 160:{28,28}]
  wire  _GEN_1691 = _GEN_2274 & ~d_way[0] ? dirty_73_0 : _GEN_1690; // @[cache.scala 160:{28,28}]
  wire  _GEN_1692 = _GEN_2274 & d_way[0] ? dirty_73_1 : _GEN_1691; // @[cache.scala 160:{28,28}]
  wire  _GEN_1693 = _GEN_2277 & ~d_way[0] ? dirty_74_0 : _GEN_1692; // @[cache.scala 160:{28,28}]
  wire  _GEN_1694 = _GEN_2277 & d_way[0] ? dirty_74_1 : _GEN_1693; // @[cache.scala 160:{28,28}]
  wire  _GEN_1695 = _GEN_2280 & ~d_way[0] ? dirty_75_0 : _GEN_1694; // @[cache.scala 160:{28,28}]
  wire  _GEN_1696 = _GEN_2280 & d_way[0] ? dirty_75_1 : _GEN_1695; // @[cache.scala 160:{28,28}]
  wire  _GEN_1697 = _GEN_2283 & ~d_way[0] ? dirty_76_0 : _GEN_1696; // @[cache.scala 160:{28,28}]
  wire  _GEN_1698 = _GEN_2283 & d_way[0] ? dirty_76_1 : _GEN_1697; // @[cache.scala 160:{28,28}]
  wire  _GEN_1699 = _GEN_2286 & ~d_way[0] ? dirty_77_0 : _GEN_1698; // @[cache.scala 160:{28,28}]
  wire  _GEN_1700 = _GEN_2286 & d_way[0] ? dirty_77_1 : _GEN_1699; // @[cache.scala 160:{28,28}]
  wire  _GEN_1701 = _GEN_2289 & ~d_way[0] ? dirty_78_0 : _GEN_1700; // @[cache.scala 160:{28,28}]
  wire  _GEN_1702 = _GEN_2289 & d_way[0] ? dirty_78_1 : _GEN_1701; // @[cache.scala 160:{28,28}]
  wire  _GEN_1703 = _GEN_2292 & ~d_way[0] ? dirty_79_0 : _GEN_1702; // @[cache.scala 160:{28,28}]
  wire  _GEN_1704 = _GEN_2292 & d_way[0] ? dirty_79_1 : _GEN_1703; // @[cache.scala 160:{28,28}]
  wire  _GEN_1705 = _GEN_2295 & ~d_way[0] ? dirty_80_0 : _GEN_1704; // @[cache.scala 160:{28,28}]
  wire  _GEN_1706 = _GEN_2295 & d_way[0] ? dirty_80_1 : _GEN_1705; // @[cache.scala 160:{28,28}]
  wire  _GEN_1707 = _GEN_2298 & ~d_way[0] ? dirty_81_0 : _GEN_1706; // @[cache.scala 160:{28,28}]
  wire  _GEN_1708 = _GEN_2298 & d_way[0] ? dirty_81_1 : _GEN_1707; // @[cache.scala 160:{28,28}]
  wire  _GEN_1709 = _GEN_2301 & ~d_way[0] ? dirty_82_0 : _GEN_1708; // @[cache.scala 160:{28,28}]
  wire  _GEN_1710 = _GEN_2301 & d_way[0] ? dirty_82_1 : _GEN_1709; // @[cache.scala 160:{28,28}]
  wire  _GEN_1711 = _GEN_2304 & ~d_way[0] ? dirty_83_0 : _GEN_1710; // @[cache.scala 160:{28,28}]
  wire  _GEN_1712 = _GEN_2304 & d_way[0] ? dirty_83_1 : _GEN_1711; // @[cache.scala 160:{28,28}]
  wire  _GEN_1713 = _GEN_2307 & ~d_way[0] ? dirty_84_0 : _GEN_1712; // @[cache.scala 160:{28,28}]
  wire  _GEN_1714 = _GEN_2307 & d_way[0] ? dirty_84_1 : _GEN_1713; // @[cache.scala 160:{28,28}]
  wire  _GEN_1715 = _GEN_2310 & ~d_way[0] ? dirty_85_0 : _GEN_1714; // @[cache.scala 160:{28,28}]
  wire  _GEN_1716 = _GEN_2310 & d_way[0] ? dirty_85_1 : _GEN_1715; // @[cache.scala 160:{28,28}]
  wire  _GEN_1717 = _GEN_2313 & ~d_way[0] ? dirty_86_0 : _GEN_1716; // @[cache.scala 160:{28,28}]
  wire  _GEN_1718 = _GEN_2313 & d_way[0] ? dirty_86_1 : _GEN_1717; // @[cache.scala 160:{28,28}]
  wire  _GEN_1719 = _GEN_2316 & ~d_way[0] ? dirty_87_0 : _GEN_1718; // @[cache.scala 160:{28,28}]
  wire  _GEN_1720 = _GEN_2316 & d_way[0] ? dirty_87_1 : _GEN_1719; // @[cache.scala 160:{28,28}]
  wire  _GEN_1721 = _GEN_2319 & ~d_way[0] ? dirty_88_0 : _GEN_1720; // @[cache.scala 160:{28,28}]
  wire  _GEN_1722 = _GEN_2319 & d_way[0] ? dirty_88_1 : _GEN_1721; // @[cache.scala 160:{28,28}]
  wire  _GEN_1723 = _GEN_2322 & ~d_way[0] ? dirty_89_0 : _GEN_1722; // @[cache.scala 160:{28,28}]
  wire  _GEN_1724 = _GEN_2322 & d_way[0] ? dirty_89_1 : _GEN_1723; // @[cache.scala 160:{28,28}]
  wire  _GEN_1725 = _GEN_2325 & ~d_way[0] ? dirty_90_0 : _GEN_1724; // @[cache.scala 160:{28,28}]
  wire  _GEN_1726 = _GEN_2325 & d_way[0] ? dirty_90_1 : _GEN_1725; // @[cache.scala 160:{28,28}]
  wire  _GEN_1727 = _GEN_2328 & ~d_way[0] ? dirty_91_0 : _GEN_1726; // @[cache.scala 160:{28,28}]
  wire  _GEN_1728 = _GEN_2328 & d_way[0] ? dirty_91_1 : _GEN_1727; // @[cache.scala 160:{28,28}]
  wire  _GEN_1729 = _GEN_2331 & ~d_way[0] ? dirty_92_0 : _GEN_1728; // @[cache.scala 160:{28,28}]
  wire  _GEN_1730 = _GEN_2331 & d_way[0] ? dirty_92_1 : _GEN_1729; // @[cache.scala 160:{28,28}]
  wire  _GEN_1731 = _GEN_2334 & ~d_way[0] ? dirty_93_0 : _GEN_1730; // @[cache.scala 160:{28,28}]
  wire  _GEN_1732 = _GEN_2334 & d_way[0] ? dirty_93_1 : _GEN_1731; // @[cache.scala 160:{28,28}]
  wire  _GEN_1733 = _GEN_2337 & ~d_way[0] ? dirty_94_0 : _GEN_1732; // @[cache.scala 160:{28,28}]
  wire  _GEN_1734 = _GEN_2337 & d_way[0] ? dirty_94_1 : _GEN_1733; // @[cache.scala 160:{28,28}]
  wire  _GEN_1735 = _GEN_2340 & ~d_way[0] ? dirty_95_0 : _GEN_1734; // @[cache.scala 160:{28,28}]
  wire  _GEN_1736 = _GEN_2340 & d_way[0] ? dirty_95_1 : _GEN_1735; // @[cache.scala 160:{28,28}]
  wire  _GEN_1737 = _GEN_2343 & ~d_way[0] ? dirty_96_0 : _GEN_1736; // @[cache.scala 160:{28,28}]
  wire  _GEN_1738 = _GEN_2343 & d_way[0] ? dirty_96_1 : _GEN_1737; // @[cache.scala 160:{28,28}]
  wire  _GEN_1739 = _GEN_2346 & ~d_way[0] ? dirty_97_0 : _GEN_1738; // @[cache.scala 160:{28,28}]
  wire  _GEN_1740 = _GEN_2346 & d_way[0] ? dirty_97_1 : _GEN_1739; // @[cache.scala 160:{28,28}]
  wire  _GEN_1741 = _GEN_2349 & ~d_way[0] ? dirty_98_0 : _GEN_1740; // @[cache.scala 160:{28,28}]
  wire  _GEN_1742 = _GEN_2349 & d_way[0] ? dirty_98_1 : _GEN_1741; // @[cache.scala 160:{28,28}]
  wire  _GEN_1743 = _GEN_2352 & ~d_way[0] ? dirty_99_0 : _GEN_1742; // @[cache.scala 160:{28,28}]
  wire  _GEN_1744 = _GEN_2352 & d_way[0] ? dirty_99_1 : _GEN_1743; // @[cache.scala 160:{28,28}]
  wire  _GEN_1745 = _GEN_2355 & ~d_way[0] ? dirty_100_0 : _GEN_1744; // @[cache.scala 160:{28,28}]
  wire  _GEN_1746 = _GEN_2355 & d_way[0] ? dirty_100_1 : _GEN_1745; // @[cache.scala 160:{28,28}]
  wire  _GEN_1747 = _GEN_2358 & ~d_way[0] ? dirty_101_0 : _GEN_1746; // @[cache.scala 160:{28,28}]
  wire  _GEN_1748 = _GEN_2358 & d_way[0] ? dirty_101_1 : _GEN_1747; // @[cache.scala 160:{28,28}]
  wire  _GEN_1749 = _GEN_2361 & ~d_way[0] ? dirty_102_0 : _GEN_1748; // @[cache.scala 160:{28,28}]
  wire  _GEN_1750 = _GEN_2361 & d_way[0] ? dirty_102_1 : _GEN_1749; // @[cache.scala 160:{28,28}]
  wire  _GEN_1751 = _GEN_2364 & ~d_way[0] ? dirty_103_0 : _GEN_1750; // @[cache.scala 160:{28,28}]
  wire  _GEN_1752 = _GEN_2364 & d_way[0] ? dirty_103_1 : _GEN_1751; // @[cache.scala 160:{28,28}]
  wire  _GEN_1753 = _GEN_2367 & ~d_way[0] ? dirty_104_0 : _GEN_1752; // @[cache.scala 160:{28,28}]
  wire  _GEN_1754 = _GEN_2367 & d_way[0] ? dirty_104_1 : _GEN_1753; // @[cache.scala 160:{28,28}]
  wire  _GEN_1755 = _GEN_2370 & ~d_way[0] ? dirty_105_0 : _GEN_1754; // @[cache.scala 160:{28,28}]
  wire  _GEN_1756 = _GEN_2370 & d_way[0] ? dirty_105_1 : _GEN_1755; // @[cache.scala 160:{28,28}]
  wire  _GEN_1757 = _GEN_2373 & ~d_way[0] ? dirty_106_0 : _GEN_1756; // @[cache.scala 160:{28,28}]
  wire  _GEN_1758 = _GEN_2373 & d_way[0] ? dirty_106_1 : _GEN_1757; // @[cache.scala 160:{28,28}]
  wire  _GEN_1759 = _GEN_2376 & ~d_way[0] ? dirty_107_0 : _GEN_1758; // @[cache.scala 160:{28,28}]
  wire  _GEN_1760 = _GEN_2376 & d_way[0] ? dirty_107_1 : _GEN_1759; // @[cache.scala 160:{28,28}]
  wire  _GEN_1761 = _GEN_2379 & ~d_way[0] ? dirty_108_0 : _GEN_1760; // @[cache.scala 160:{28,28}]
  wire  _GEN_1762 = _GEN_2379 & d_way[0] ? dirty_108_1 : _GEN_1761; // @[cache.scala 160:{28,28}]
  wire  _GEN_1763 = _GEN_2382 & ~d_way[0] ? dirty_109_0 : _GEN_1762; // @[cache.scala 160:{28,28}]
  wire  _GEN_1764 = _GEN_2382 & d_way[0] ? dirty_109_1 : _GEN_1763; // @[cache.scala 160:{28,28}]
  wire  _GEN_1765 = _GEN_2385 & ~d_way[0] ? dirty_110_0 : _GEN_1764; // @[cache.scala 160:{28,28}]
  wire  _GEN_1766 = _GEN_2385 & d_way[0] ? dirty_110_1 : _GEN_1765; // @[cache.scala 160:{28,28}]
  wire  _GEN_1767 = _GEN_2388 & ~d_way[0] ? dirty_111_0 : _GEN_1766; // @[cache.scala 160:{28,28}]
  wire  _GEN_1768 = _GEN_2388 & d_way[0] ? dirty_111_1 : _GEN_1767; // @[cache.scala 160:{28,28}]
  wire  _GEN_1769 = _GEN_2391 & ~d_way[0] ? dirty_112_0 : _GEN_1768; // @[cache.scala 160:{28,28}]
  wire  _GEN_1770 = _GEN_2391 & d_way[0] ? dirty_112_1 : _GEN_1769; // @[cache.scala 160:{28,28}]
  wire  _GEN_1771 = _GEN_2394 & ~d_way[0] ? dirty_113_0 : _GEN_1770; // @[cache.scala 160:{28,28}]
  wire  _GEN_1772 = _GEN_2394 & d_way[0] ? dirty_113_1 : _GEN_1771; // @[cache.scala 160:{28,28}]
  wire  _GEN_1773 = _GEN_2397 & ~d_way[0] ? dirty_114_0 : _GEN_1772; // @[cache.scala 160:{28,28}]
  wire  _GEN_1774 = _GEN_2397 & d_way[0] ? dirty_114_1 : _GEN_1773; // @[cache.scala 160:{28,28}]
  wire  _GEN_1775 = _GEN_2400 & ~d_way[0] ? dirty_115_0 : _GEN_1774; // @[cache.scala 160:{28,28}]
  wire  _GEN_1776 = _GEN_2400 & d_way[0] ? dirty_115_1 : _GEN_1775; // @[cache.scala 160:{28,28}]
  wire  _GEN_1777 = _GEN_2403 & ~d_way[0] ? dirty_116_0 : _GEN_1776; // @[cache.scala 160:{28,28}]
  wire  _GEN_1778 = _GEN_2403 & d_way[0] ? dirty_116_1 : _GEN_1777; // @[cache.scala 160:{28,28}]
  wire  _GEN_1779 = _GEN_2406 & ~d_way[0] ? dirty_117_0 : _GEN_1778; // @[cache.scala 160:{28,28}]
  wire  _GEN_1780 = _GEN_2406 & d_way[0] ? dirty_117_1 : _GEN_1779; // @[cache.scala 160:{28,28}]
  wire  _GEN_1781 = _GEN_2409 & ~d_way[0] ? dirty_118_0 : _GEN_1780; // @[cache.scala 160:{28,28}]
  wire  _GEN_1782 = _GEN_2409 & d_way[0] ? dirty_118_1 : _GEN_1781; // @[cache.scala 160:{28,28}]
  wire  _GEN_1783 = _GEN_2412 & ~d_way[0] ? dirty_119_0 : _GEN_1782; // @[cache.scala 160:{28,28}]
  wire  _GEN_1784 = _GEN_2412 & d_way[0] ? dirty_119_1 : _GEN_1783; // @[cache.scala 160:{28,28}]
  wire  _GEN_1785 = _GEN_2415 & ~d_way[0] ? dirty_120_0 : _GEN_1784; // @[cache.scala 160:{28,28}]
  wire  _GEN_1786 = _GEN_2415 & d_way[0] ? dirty_120_1 : _GEN_1785; // @[cache.scala 160:{28,28}]
  wire  _GEN_1787 = _GEN_2418 & ~d_way[0] ? dirty_121_0 : _GEN_1786; // @[cache.scala 160:{28,28}]
  wire  _GEN_1788 = _GEN_2418 & d_way[0] ? dirty_121_1 : _GEN_1787; // @[cache.scala 160:{28,28}]
  wire  _GEN_1789 = _GEN_2421 & ~d_way[0] ? dirty_122_0 : _GEN_1788; // @[cache.scala 160:{28,28}]
  wire  _GEN_1790 = _GEN_2421 & d_way[0] ? dirty_122_1 : _GEN_1789; // @[cache.scala 160:{28,28}]
  wire  _GEN_1791 = _GEN_2424 & ~d_way[0] ? dirty_123_0 : _GEN_1790; // @[cache.scala 160:{28,28}]
  wire  _GEN_1792 = _GEN_2424 & d_way[0] ? dirty_123_1 : _GEN_1791; // @[cache.scala 160:{28,28}]
  wire  _GEN_1793 = _GEN_2427 & ~d_way[0] ? dirty_124_0 : _GEN_1792; // @[cache.scala 160:{28,28}]
  wire  _GEN_1794 = _GEN_2427 & d_way[0] ? dirty_124_1 : _GEN_1793; // @[cache.scala 160:{28,28}]
  wire  _GEN_1795 = _GEN_2430 & ~d_way[0] ? dirty_125_0 : _GEN_1794; // @[cache.scala 160:{28,28}]
  wire  _GEN_1796 = _GEN_2430 & d_way[0] ? dirty_125_1 : _GEN_1795; // @[cache.scala 160:{28,28}]
  wire  _GEN_1797 = _GEN_2433 & ~d_way[0] ? dirty_126_0 : _GEN_1796; // @[cache.scala 160:{28,28}]
  wire  _GEN_1798 = _GEN_2433 & d_way[0] ? dirty_126_1 : _GEN_1797; // @[cache.scala 160:{28,28}]
  wire  _GEN_1799 = _GEN_2436 & ~d_way[0] ? dirty_127_0 : _GEN_1798; // @[cache.scala 160:{28,28}]
  wire  _GEN_1800 = _GEN_2436 & d_way[0] ? dirty_127_1 : _GEN_1799; // @[cache.scala 160:{28,28}]
  wire  _dirty_T_5 = _io_in_r_bits_data_T_3 ? 1'h0 : _GEN_1800; // @[cache.scala 160:28]
  wire [63:0] _wstrb_map_T_8 = wstrb == 128'hff ? 64'hffffffffffffffff : 64'h0; // @[cache.scala 167:20]
  wire [63:0] _wstrb_map_T_9 = wstrb == 128'hf ? 64'hffffffff : _wstrb_map_T_8; // @[cache.scala 166:20]
  wire [63:0] _wstrb_map_T_10 = wstrb == 128'h3 ? 64'hffff : _wstrb_map_T_9; // @[cache.scala 165:20]
  wire [63:0] _wstrb_map_T_11 = wstrb == 128'h1 ? 64'hff : _wstrb_map_T_10; // @[cache.scala 164:20]
  wire [190:0] _GEN_0 = {{127'd0}, _wstrb_map_T_11}; // @[cache.scala 167:68]
  wire [190:0] _wstrb_map_T_12 = _GEN_0 << offset; // @[cache.scala 167:68]
  wire [254:0] _GEN_1 = {{127'd0}, wdata}; // @[cache.scala 170:22]
  wire [254:0] _wdata_map_T = _GEN_1 << offset; // @[cache.scala 170:22]
  wire  _io_ram_bits_CEN_T = state == 4'h2; // @[cache.scala 174:28]
  wire  _io_ram_bits_CEN_T_3 = state_w != 4'h0 & state_w != 4'h9; // @[cache.scala 174:61]
  wire [127:0] wstrb_map = _wstrb_map_T_12[127:0]; // @[cache.scala 163:23 164:13]
  wire [7:0] _io_ram_bits_A_T_10 = _io_ram_bits_CEN_T_3 | _io_in_r_bits_data_T_3 ? idxw : 8'h0; // @[cache.scala 178:22]
  wire [127:0] _io_ram_bits_D_T_4 = ~wstrb_map; // @[cache.scala 181:43]
  wire [127:0] _io_ram_bits_D_T_5 = buf_ & _io_ram_bits_D_T_4; // @[cache.scala 181:41]
  wire [127:0] wdata_map = _wdata_map_T[127:0]; // @[cache.scala 169:23 170:13]
  wire [127:0] _io_ram_bits_D_T_6 = wdata_map & wstrb_map; // @[cache.scala 181:66]
  wire [127:0] _io_ram_bits_D_T_7 = _io_ram_bits_D_T_5 | _io_ram_bits_D_T_6; // @[cache.scala 181:55]
  wire [127:0] _io_ram_bits_D_T_8 = wmode ? _io_ram_bits_D_T_7 : buf_; // @[cache.scala 181:22]
  reg [31:0] cnt; // @[cache.scala 193:18]
  reg [31:0] hit; // @[cache.scala 194:18]
  wire [31:0] _cnt_T_2 = cnt + 32'h1; // @[cache.scala 195:33]
  wire [31:0] _hit_T_2 = hit + 32'h1; // @[cache.scala 196:31]
  LFSR_8 lfsr8 ( // @[cache.scala 61:21]
    .clock(lfsr8_clock),
    .reset(lfsr8_reset),
    .io_out(lfsr8_io_out)
  );
  assign cache_tag_tag_read_MPORT_en = cache_tag_tag_read_MPORT_en_pipe_0;
  assign cache_tag_tag_read_MPORT_addr = cache_tag_tag_read_MPORT_addr_pipe_0;
  assign cache_tag_tag_read_MPORT_data = cache_tag[cache_tag_tag_read_MPORT_addr]; // @[cache.scala 24:30]
  assign cache_tag_MPORT_data = _tag_way_T ? _tagg_T_2 : _tagg_T_4;
  assign cache_tag_MPORT_addr = addr[10:4];
  assign cache_tag_MPORT_mask = 1'h1;
  assign cache_tag_MPORT_en = state == 4'h5;
  assign io_in_ar_ready = state == 4'h0; // @[cache.scala 84:28]
  assign io_in_r_valid = (_io_in_r_bits_data_T | _io_in_r_bits_data_T_3) & rmode; // @[cache.scala 85:64]
  assign io_in_r_bits_data = _io_in_r_bits_data_T_6[63:0]; // @[cache.scala 81:21]
  assign io_in_aw_ready = state == 4'h0; // @[cache.scala 89:28]
  assign io_in_w_ready = 1'h1; // @[cache.scala 90:17]
  assign io_in_b_valid = (_io_in_r_bits_data_T_3 | _io_in_r_bits_data_T) & wmode; // @[cache.scala 88:60]
  assign io_mem_ar_valid = state_r == 4'h0 & _state_r_T; // @[cache.scala 132:41]
  assign io_mem_ar_bits_addr = _io_mem_ar_bits_addr_T_2[31:0]; // @[cache.scala 131:23]
  assign io_mem_r_ready = 1'h1; // @[cache.scala 136:18]
  assign io_mem_aw_valid = state_w == 4'h0 & _GEN_515 & _state_r_T; // @[cache.scala 119:70]
  assign io_mem_aw_bits_addr = {_io_mem_aw_bits_addr_T_1, 4'h0}; // @[cache.scala 116:55]
  assign io_mem_w_valid = _io_mem_w_bits_data_T | state_w == 4'h6; // @[cache.scala 128:41]
  assign io_mem_w_bits_data = state_w == 4'h7 ? io_ram_bits_Q[127:64] : io_ram_bits_Q[63:0]; // @[cache.scala 125:28]
  assign io_mem_w_bits_last = state_w == 4'h7; // @[cache.scala 127:33]
  assign io_mem_b_ready = 1'h1; // @[cache.scala 129:18]
  assign io_ram_bits_CEN = state == 4'h2 | state_w != 4'h0 & state_w != 4'h9 | _io_in_r_bits_data_T_3 | _d_way_T_2; // @[cache.scala 174:106]
  assign io_ram_bits_WEN = _io_in_r_bits_data_T_3 | _d_way_T_2; // @[cache.scala 175:42]
  assign io_ram_bits_BWEN = _d_way_T_2 ? wstrb_map : 128'hffffffffffffffffffffffffffffffff; // @[cache.scala 176:25]
  assign io_ram_bits_A = _io_ram_bits_CEN_T | _d_way_T_2 ? idxh : _io_ram_bits_A_T_10; // @[cache.scala 177:22]
  assign io_ram_bits_D = _d_way_T_2 ? wdata_map : _io_ram_bits_D_T_8; // @[cache.scala 180:22]
  assign io_hitrate = {cnt,hit}; // @[Cat.scala 33:92]
  assign lfsr8_clock = clock;
  assign lfsr8_reset = reset;
  always @(posedge clock) begin
    if (cache_tag_MPORT_en & cache_tag_MPORT_mask) begin
      cache_tag[cache_tag_MPORT_addr] <= cache_tag_MPORT_data; // @[cache.scala 24:30]
    end
    cache_tag_tag_read_MPORT_en_pipe_0 <= state != 4'h5;
    if (state != 4'h5) begin
      cache_tag_tag_read_MPORT_addr_pipe_0 <= addr[10:4];
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_0_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2057 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_0_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_0_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2057 & way2[0]) begin // @[cache.scala 154:20]
      valid_0_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_1_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2058 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_1_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_1_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2058 & way2[0]) begin // @[cache.scala 154:20]
      valid_1_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_2_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2061 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_2_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_2_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2061 & way2[0]) begin // @[cache.scala 154:20]
      valid_2_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_3_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2064 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_3_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_3_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2064 & way2[0]) begin // @[cache.scala 154:20]
      valid_3_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_4_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2067 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_4_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_4_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2067 & way2[0]) begin // @[cache.scala 154:20]
      valid_4_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_5_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2070 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_5_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_5_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2070 & way2[0]) begin // @[cache.scala 154:20]
      valid_5_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_6_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2073 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_6_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_6_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2073 & way2[0]) begin // @[cache.scala 154:20]
      valid_6_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_7_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2076 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_7_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_7_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2076 & way2[0]) begin // @[cache.scala 154:20]
      valid_7_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_8_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2079 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_8_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_8_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2079 & way2[0]) begin // @[cache.scala 154:20]
      valid_8_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_9_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2082 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_9_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_9_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2082 & way2[0]) begin // @[cache.scala 154:20]
      valid_9_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_10_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2085 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_10_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_10_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2085 & way2[0]) begin // @[cache.scala 154:20]
      valid_10_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_11_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2088 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_11_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_11_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2088 & way2[0]) begin // @[cache.scala 154:20]
      valid_11_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_12_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2091 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_12_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_12_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2091 & way2[0]) begin // @[cache.scala 154:20]
      valid_12_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_13_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2094 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_13_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_13_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2094 & way2[0]) begin // @[cache.scala 154:20]
      valid_13_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_14_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2097 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_14_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_14_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2097 & way2[0]) begin // @[cache.scala 154:20]
      valid_14_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_15_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2100 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_15_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_15_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2100 & way2[0]) begin // @[cache.scala 154:20]
      valid_15_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_16_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2103 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_16_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_16_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2103 & way2[0]) begin // @[cache.scala 154:20]
      valid_16_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_17_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2106 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_17_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_17_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2106 & way2[0]) begin // @[cache.scala 154:20]
      valid_17_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_18_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2109 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_18_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_18_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2109 & way2[0]) begin // @[cache.scala 154:20]
      valid_18_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_19_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2112 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_19_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_19_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2112 & way2[0]) begin // @[cache.scala 154:20]
      valid_19_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_20_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2115 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_20_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_20_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2115 & way2[0]) begin // @[cache.scala 154:20]
      valid_20_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_21_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2118 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_21_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_21_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2118 & way2[0]) begin // @[cache.scala 154:20]
      valid_21_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_22_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2121 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_22_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_22_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2121 & way2[0]) begin // @[cache.scala 154:20]
      valid_22_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_23_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2124 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_23_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_23_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2124 & way2[0]) begin // @[cache.scala 154:20]
      valid_23_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_24_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2127 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_24_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_24_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2127 & way2[0]) begin // @[cache.scala 154:20]
      valid_24_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_25_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2130 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_25_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_25_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2130 & way2[0]) begin // @[cache.scala 154:20]
      valid_25_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_26_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2133 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_26_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_26_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2133 & way2[0]) begin // @[cache.scala 154:20]
      valid_26_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_27_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2136 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_27_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_27_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2136 & way2[0]) begin // @[cache.scala 154:20]
      valid_27_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_28_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2139 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_28_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_28_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2139 & way2[0]) begin // @[cache.scala 154:20]
      valid_28_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_29_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2142 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_29_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_29_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2142 & way2[0]) begin // @[cache.scala 154:20]
      valid_29_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_30_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2145 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_30_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_30_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2145 & way2[0]) begin // @[cache.scala 154:20]
      valid_30_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_31_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2148 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_31_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_31_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2148 & way2[0]) begin // @[cache.scala 154:20]
      valid_31_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_32_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2151 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_32_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_32_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2151 & way2[0]) begin // @[cache.scala 154:20]
      valid_32_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_33_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2154 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_33_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_33_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2154 & way2[0]) begin // @[cache.scala 154:20]
      valid_33_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_34_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2157 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_34_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_34_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2157 & way2[0]) begin // @[cache.scala 154:20]
      valid_34_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_35_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2160 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_35_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_35_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2160 & way2[0]) begin // @[cache.scala 154:20]
      valid_35_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_36_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2163 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_36_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_36_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2163 & way2[0]) begin // @[cache.scala 154:20]
      valid_36_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_37_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2166 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_37_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_37_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2166 & way2[0]) begin // @[cache.scala 154:20]
      valid_37_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_38_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2169 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_38_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_38_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2169 & way2[0]) begin // @[cache.scala 154:20]
      valid_38_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_39_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2172 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_39_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_39_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2172 & way2[0]) begin // @[cache.scala 154:20]
      valid_39_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_40_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2175 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_40_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_40_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2175 & way2[0]) begin // @[cache.scala 154:20]
      valid_40_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_41_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2178 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_41_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_41_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2178 & way2[0]) begin // @[cache.scala 154:20]
      valid_41_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_42_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2181 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_42_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_42_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2181 & way2[0]) begin // @[cache.scala 154:20]
      valid_42_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_43_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2184 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_43_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_43_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2184 & way2[0]) begin // @[cache.scala 154:20]
      valid_43_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_44_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2187 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_44_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_44_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2187 & way2[0]) begin // @[cache.scala 154:20]
      valid_44_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_45_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2190 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_45_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_45_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2190 & way2[0]) begin // @[cache.scala 154:20]
      valid_45_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_46_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2193 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_46_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_46_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2193 & way2[0]) begin // @[cache.scala 154:20]
      valid_46_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_47_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2196 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_47_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_47_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2196 & way2[0]) begin // @[cache.scala 154:20]
      valid_47_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_48_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2199 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_48_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_48_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2199 & way2[0]) begin // @[cache.scala 154:20]
      valid_48_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_49_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2202 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_49_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_49_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2202 & way2[0]) begin // @[cache.scala 154:20]
      valid_49_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_50_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2205 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_50_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_50_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2205 & way2[0]) begin // @[cache.scala 154:20]
      valid_50_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_51_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2208 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_51_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_51_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2208 & way2[0]) begin // @[cache.scala 154:20]
      valid_51_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_52_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2211 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_52_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_52_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2211 & way2[0]) begin // @[cache.scala 154:20]
      valid_52_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_53_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2214 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_53_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_53_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2214 & way2[0]) begin // @[cache.scala 154:20]
      valid_53_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_54_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2217 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_54_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_54_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2217 & way2[0]) begin // @[cache.scala 154:20]
      valid_54_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_55_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2220 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_55_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_55_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2220 & way2[0]) begin // @[cache.scala 154:20]
      valid_55_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_56_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2223 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_56_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_56_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2223 & way2[0]) begin // @[cache.scala 154:20]
      valid_56_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_57_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2226 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_57_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_57_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2226 & way2[0]) begin // @[cache.scala 154:20]
      valid_57_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_58_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2229 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_58_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_58_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2229 & way2[0]) begin // @[cache.scala 154:20]
      valid_58_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_59_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2232 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_59_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_59_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2232 & way2[0]) begin // @[cache.scala 154:20]
      valid_59_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_60_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2235 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_60_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_60_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2235 & way2[0]) begin // @[cache.scala 154:20]
      valid_60_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_61_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2238 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_61_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_61_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2238 & way2[0]) begin // @[cache.scala 154:20]
      valid_61_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_62_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2241 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_62_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_62_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2241 & way2[0]) begin // @[cache.scala 154:20]
      valid_62_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_63_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2244 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_63_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_63_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2244 & way2[0]) begin // @[cache.scala 154:20]
      valid_63_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_64_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2247 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_64_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_64_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2247 & way2[0]) begin // @[cache.scala 154:20]
      valid_64_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_65_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2250 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_65_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_65_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2250 & way2[0]) begin // @[cache.scala 154:20]
      valid_65_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_66_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2253 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_66_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_66_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2253 & way2[0]) begin // @[cache.scala 154:20]
      valid_66_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_67_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2256 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_67_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_67_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2256 & way2[0]) begin // @[cache.scala 154:20]
      valid_67_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_68_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2259 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_68_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_68_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2259 & way2[0]) begin // @[cache.scala 154:20]
      valid_68_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_69_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2262 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_69_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_69_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2262 & way2[0]) begin // @[cache.scala 154:20]
      valid_69_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_70_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2265 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_70_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_70_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2265 & way2[0]) begin // @[cache.scala 154:20]
      valid_70_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_71_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2268 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_71_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_71_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2268 & way2[0]) begin // @[cache.scala 154:20]
      valid_71_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_72_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2271 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_72_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_72_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2271 & way2[0]) begin // @[cache.scala 154:20]
      valid_72_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_73_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2274 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_73_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_73_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2274 & way2[0]) begin // @[cache.scala 154:20]
      valid_73_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_74_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2277 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_74_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_74_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2277 & way2[0]) begin // @[cache.scala 154:20]
      valid_74_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_75_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2280 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_75_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_75_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2280 & way2[0]) begin // @[cache.scala 154:20]
      valid_75_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_76_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2283 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_76_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_76_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2283 & way2[0]) begin // @[cache.scala 154:20]
      valid_76_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_77_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2286 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_77_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_77_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2286 & way2[0]) begin // @[cache.scala 154:20]
      valid_77_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_78_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2289 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_78_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_78_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2289 & way2[0]) begin // @[cache.scala 154:20]
      valid_78_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_79_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2292 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_79_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_79_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2292 & way2[0]) begin // @[cache.scala 154:20]
      valid_79_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_80_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2295 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_80_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_80_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2295 & way2[0]) begin // @[cache.scala 154:20]
      valid_80_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_81_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2298 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_81_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_81_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2298 & way2[0]) begin // @[cache.scala 154:20]
      valid_81_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_82_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2301 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_82_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_82_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2301 & way2[0]) begin // @[cache.scala 154:20]
      valid_82_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_83_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2304 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_83_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_83_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2304 & way2[0]) begin // @[cache.scala 154:20]
      valid_83_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_84_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2307 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_84_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_84_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2307 & way2[0]) begin // @[cache.scala 154:20]
      valid_84_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_85_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2310 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_85_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_85_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2310 & way2[0]) begin // @[cache.scala 154:20]
      valid_85_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_86_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2313 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_86_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_86_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2313 & way2[0]) begin // @[cache.scala 154:20]
      valid_86_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_87_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2316 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_87_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_87_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2316 & way2[0]) begin // @[cache.scala 154:20]
      valid_87_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_88_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2319 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_88_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_88_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2319 & way2[0]) begin // @[cache.scala 154:20]
      valid_88_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_89_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2322 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_89_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_89_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2322 & way2[0]) begin // @[cache.scala 154:20]
      valid_89_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_90_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2325 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_90_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_90_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2325 & way2[0]) begin // @[cache.scala 154:20]
      valid_90_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_91_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2328 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_91_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_91_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2328 & way2[0]) begin // @[cache.scala 154:20]
      valid_91_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_92_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2331 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_92_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_92_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2331 & way2[0]) begin // @[cache.scala 154:20]
      valid_92_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_93_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2334 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_93_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_93_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2334 & way2[0]) begin // @[cache.scala 154:20]
      valid_93_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_94_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2337 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_94_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_94_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2337 & way2[0]) begin // @[cache.scala 154:20]
      valid_94_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_95_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2340 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_95_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_95_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2340 & way2[0]) begin // @[cache.scala 154:20]
      valid_95_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_96_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2343 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_96_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_96_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2343 & way2[0]) begin // @[cache.scala 154:20]
      valid_96_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_97_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2346 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_97_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_97_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2346 & way2[0]) begin // @[cache.scala 154:20]
      valid_97_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_98_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2349 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_98_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_98_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2349 & way2[0]) begin // @[cache.scala 154:20]
      valid_98_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_99_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2352 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_99_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_99_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2352 & way2[0]) begin // @[cache.scala 154:20]
      valid_99_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_100_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2355 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_100_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_100_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2355 & way2[0]) begin // @[cache.scala 154:20]
      valid_100_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_101_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2358 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_101_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_101_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2358 & way2[0]) begin // @[cache.scala 154:20]
      valid_101_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_102_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2361 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_102_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_102_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2361 & way2[0]) begin // @[cache.scala 154:20]
      valid_102_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_103_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2364 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_103_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_103_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2364 & way2[0]) begin // @[cache.scala 154:20]
      valid_103_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_104_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2367 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_104_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_104_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2367 & way2[0]) begin // @[cache.scala 154:20]
      valid_104_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_105_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2370 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_105_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_105_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2370 & way2[0]) begin // @[cache.scala 154:20]
      valid_105_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_106_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2373 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_106_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_106_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2373 & way2[0]) begin // @[cache.scala 154:20]
      valid_106_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_107_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2376 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_107_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_107_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2376 & way2[0]) begin // @[cache.scala 154:20]
      valid_107_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_108_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2379 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_108_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_108_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2379 & way2[0]) begin // @[cache.scala 154:20]
      valid_108_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_109_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2382 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_109_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_109_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2382 & way2[0]) begin // @[cache.scala 154:20]
      valid_109_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_110_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2385 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_110_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_110_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2385 & way2[0]) begin // @[cache.scala 154:20]
      valid_110_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_111_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2388 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_111_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_111_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2388 & way2[0]) begin // @[cache.scala 154:20]
      valid_111_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_112_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2391 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_112_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_112_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2391 & way2[0]) begin // @[cache.scala 154:20]
      valid_112_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_113_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2394 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_113_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_113_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2394 & way2[0]) begin // @[cache.scala 154:20]
      valid_113_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_114_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2397 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_114_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_114_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2397 & way2[0]) begin // @[cache.scala 154:20]
      valid_114_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_115_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2400 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_115_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_115_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2400 & way2[0]) begin // @[cache.scala 154:20]
      valid_115_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_116_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2403 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_116_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_116_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2403 & way2[0]) begin // @[cache.scala 154:20]
      valid_116_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_117_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2406 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_117_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_117_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2406 & way2[0]) begin // @[cache.scala 154:20]
      valid_117_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_118_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2409 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_118_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_118_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2409 & way2[0]) begin // @[cache.scala 154:20]
      valid_118_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_119_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2412 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_119_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_119_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2412 & way2[0]) begin // @[cache.scala 154:20]
      valid_119_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_120_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2415 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_120_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_120_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2415 & way2[0]) begin // @[cache.scala 154:20]
      valid_120_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_121_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2418 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_121_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_121_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2418 & way2[0]) begin // @[cache.scala 154:20]
      valid_121_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_122_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2421 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_122_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_122_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2421 & way2[0]) begin // @[cache.scala 154:20]
      valid_122_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_123_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2424 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_123_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_123_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2424 & way2[0]) begin // @[cache.scala 154:20]
      valid_123_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_124_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2427 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_124_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_124_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2427 & way2[0]) begin // @[cache.scala 154:20]
      valid_124_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_125_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2430 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_125_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_125_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2430 & way2[0]) begin // @[cache.scala 154:20]
      valid_125_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_126_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2433 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_126_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_126_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2433 & way2[0]) begin // @[cache.scala 154:20]
      valid_126_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_127_0 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2436 & _GEN_2059) begin // @[cache.scala 154:20]
      valid_127_0 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 25:22]
      valid_127_1 <= 1'h0; // @[cache.scala 25:22]
    end else if (_GEN_2436 & way2[0]) begin // @[cache.scala 154:20]
      valid_127_1 <= _io_in_r_bits_data_T_3 | _GEN_1288; // @[cache.scala 154:20]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_0_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2057 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_0_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_0_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2057 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_0_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_1_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2058 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_1_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_1_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2058 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_1_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_2_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2061 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_2_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_2_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2061 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_2_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_3_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2064 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_3_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_3_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2064 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_3_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_4_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2067 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_4_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_4_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2067 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_4_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_5_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2070 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_5_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_5_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2070 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_5_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_6_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2073 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_6_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_6_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2073 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_6_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_7_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2076 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_7_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_7_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2076 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_7_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_8_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2079 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_8_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_8_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2079 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_8_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_9_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2082 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_9_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_9_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2082 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_9_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_10_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2085 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_10_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_10_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2085 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_10_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_11_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2088 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_11_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_11_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2088 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_11_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_12_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2091 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_12_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_12_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2091 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_12_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_13_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2094 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_13_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_13_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2094 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_13_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_14_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2097 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_14_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_14_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2097 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_14_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_15_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2100 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_15_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_15_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2100 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_15_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_16_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2103 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_16_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_16_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2103 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_16_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_17_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2106 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_17_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_17_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2106 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_17_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_18_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2109 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_18_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_18_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2109 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_18_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_19_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2112 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_19_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_19_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2112 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_19_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_20_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2115 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_20_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_20_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2115 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_20_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_21_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2118 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_21_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_21_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2118 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_21_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_22_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2121 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_22_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_22_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2121 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_22_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_23_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2124 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_23_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_23_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2124 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_23_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_24_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2127 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_24_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_24_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2127 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_24_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_25_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2130 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_25_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_25_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2130 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_25_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_26_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2133 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_26_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_26_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2133 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_26_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_27_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2136 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_27_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_27_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2136 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_27_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_28_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2139 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_28_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_28_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2139 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_28_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_29_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2142 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_29_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_29_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2142 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_29_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_30_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2145 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_30_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_30_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2145 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_30_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_31_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2148 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_31_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_31_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2148 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_31_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_32_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2151 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_32_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_32_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2151 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_32_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_33_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2154 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_33_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_33_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2154 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_33_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_34_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2157 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_34_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_34_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2157 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_34_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_35_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2160 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_35_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_35_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2160 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_35_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_36_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2163 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_36_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_36_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2163 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_36_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_37_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2166 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_37_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_37_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2166 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_37_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_38_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2169 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_38_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_38_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2169 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_38_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_39_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2172 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_39_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_39_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2172 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_39_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_40_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2175 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_40_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_40_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2175 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_40_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_41_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2178 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_41_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_41_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2178 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_41_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_42_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2181 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_42_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_42_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2181 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_42_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_43_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2184 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_43_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_43_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2184 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_43_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_44_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2187 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_44_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_44_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2187 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_44_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_45_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2190 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_45_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_45_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2190 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_45_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_46_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2193 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_46_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_46_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2193 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_46_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_47_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2196 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_47_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_47_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2196 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_47_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_48_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2199 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_48_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_48_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2199 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_48_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_49_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2202 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_49_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_49_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2202 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_49_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_50_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2205 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_50_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_50_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2205 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_50_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_51_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2208 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_51_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_51_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2208 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_51_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_52_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2211 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_52_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_52_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2211 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_52_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_53_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2214 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_53_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_53_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2214 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_53_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_54_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2217 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_54_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_54_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2217 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_54_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_55_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2220 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_55_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_55_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2220 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_55_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_56_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2223 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_56_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_56_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2223 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_56_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_57_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2226 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_57_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_57_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2226 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_57_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_58_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2229 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_58_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_58_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2229 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_58_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_59_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2232 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_59_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_59_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2232 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_59_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_60_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2235 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_60_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_60_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2235 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_60_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_61_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2238 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_61_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_61_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2238 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_61_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_62_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2241 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_62_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_62_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2241 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_62_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_63_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2244 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_63_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_63_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2244 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_63_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_64_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2247 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_64_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_64_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2247 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_64_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_65_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2250 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_65_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_65_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2250 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_65_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_66_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2253 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_66_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_66_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2253 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_66_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_67_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2256 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_67_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_67_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2256 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_67_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_68_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2259 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_68_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_68_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2259 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_68_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_69_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2262 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_69_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_69_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2262 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_69_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_70_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2265 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_70_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_70_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2265 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_70_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_71_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2268 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_71_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_71_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2268 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_71_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_72_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2271 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_72_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_72_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2271 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_72_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_73_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2274 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_73_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_73_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2274 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_73_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_74_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2277 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_74_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_74_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2277 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_74_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_75_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2280 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_75_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_75_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2280 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_75_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_76_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2283 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_76_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_76_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2283 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_76_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_77_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2286 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_77_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_77_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2286 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_77_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_78_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2289 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_78_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_78_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2289 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_78_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_79_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2292 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_79_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_79_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2292 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_79_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_80_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2295 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_80_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_80_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2295 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_80_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_81_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2298 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_81_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_81_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2298 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_81_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_82_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2301 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_82_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_82_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2301 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_82_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_83_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2304 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_83_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_83_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2304 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_83_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_84_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2307 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_84_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_84_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2307 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_84_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_85_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2310 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_85_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_85_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2310 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_85_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_86_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2313 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_86_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_86_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2313 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_86_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_87_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2316 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_87_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_87_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2316 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_87_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_88_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2319 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_88_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_88_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2319 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_88_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_89_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2322 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_89_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_89_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2322 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_89_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_90_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2325 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_90_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_90_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2325 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_90_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_91_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2328 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_91_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_91_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2328 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_91_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_92_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2331 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_92_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_92_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2331 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_92_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_93_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2334 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_93_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_93_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2334 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_93_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_94_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2337 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_94_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_94_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2337 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_94_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_95_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2340 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_95_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_95_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2340 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_95_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_96_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2343 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_96_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_96_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2343 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_96_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_97_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2346 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_97_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_97_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2346 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_97_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_98_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2349 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_98_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_98_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2349 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_98_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_99_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2352 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_99_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_99_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2352 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_99_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_100_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2355 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_100_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_100_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2355 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_100_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_101_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2358 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_101_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_101_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2358 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_101_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_102_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2361 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_102_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_102_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2361 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_102_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_103_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2364 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_103_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_103_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2364 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_103_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_104_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2367 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_104_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_104_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2367 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_104_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_105_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2370 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_105_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_105_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2370 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_105_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_106_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2373 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_106_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_106_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2373 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_106_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_107_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2376 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_107_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_107_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2376 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_107_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_108_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2379 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_108_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_108_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2379 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_108_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_109_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2382 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_109_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_109_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2382 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_109_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_110_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2385 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_110_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_110_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2385 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_110_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_111_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2388 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_111_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_111_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2388 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_111_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_112_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2391 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_112_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_112_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2391 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_112_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_113_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2394 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_113_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_113_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2394 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_113_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_114_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2397 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_114_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_114_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2397 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_114_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_115_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2400 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_115_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_115_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2400 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_115_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_116_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2403 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_116_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_116_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2403 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_116_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_117_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2406 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_117_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_117_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2406 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_117_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_118_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2409 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_118_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_118_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2409 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_118_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_119_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2412 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_119_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_119_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2412 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_119_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_120_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2415 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_120_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_120_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2415 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_120_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_121_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2418 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_121_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_121_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2418 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_121_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_122_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2421 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_122_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_122_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2421 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_122_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_123_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2424 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_123_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_123_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2424 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_123_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_124_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2427 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_124_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_124_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2427 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_124_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_125_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2430 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_125_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_125_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2430 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_125_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_126_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2433 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_126_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_126_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2433 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_126_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_127_0 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2436 & _GEN_3973) begin // @[cache.scala 159:21]
      dirty_127_0 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 26:22]
      dirty_127_1 <= 1'h0; // @[cache.scala 26:22]
    end else if (_GEN_2436 & d_way[0]) begin // @[cache.scala 159:21]
      dirty_127_1 <= _d_way_T_2 | _dirty_T_5; // @[cache.scala 159:21]
    end
    if (reset) begin // @[cache.scala 27:20]
      buf_ <= 128'h0; // @[cache.scala 27:20]
    end else if (!(_buf_T_1)) begin // @[cache.scala 143:13]
      if (rcnt == addr[3]) begin // @[cache.scala 146:8]
        buf_ <= _buf_T_5;
      end else begin
        buf_ <= _buf_T_7;
      end
    end
    if (reset) begin // @[cache.scala 29:21]
      addr <= 32'h0; // @[cache.scala 29:21]
    end else if (_rmode_T_2) begin // @[cache.scala 75:14]
      addr <= io_in_ar_bits_addr;
    end else if (_wmode_T_2) begin // @[cache.scala 76:14]
      addr <= io_in_aw_bits_addr;
    end
    if (reset) begin // @[cache.scala 30:22]
      wdata <= 128'h0; // @[cache.scala 30:22]
    end else if (state == 4'h1 & _wdata_T_1) begin // @[cache.scala 78:15]
      wdata <= {{64'd0}, io_in_w_bits_data};
    end
    if (reset) begin // @[cache.scala 31:22]
      wstrb <= 128'h0; // @[cache.scala 31:22]
    end else if (_wdata_T_2) begin // @[cache.scala 79:15]
      wstrb <= {{120'd0}, io_in_w_bits_strb};
    end
    if (reset) begin // @[cache.scala 37:21]
      way2 <= 8'h0; // @[cache.scala 37:21]
    end else if (_rmode_T) begin // @[cache.scala 62:14]
      way2 <= {{7'd0}, lfsr8_io_out[0]};
    end
    if (reset) begin // @[cache.scala 40:22]
      state <= 4'h0; // @[cache.scala 40:22]
    end else if (4'h5 == state) begin // @[Mux.scala 81:58]
      state <= 4'h0;
    end else if (4'h4 == state) begin // @[Mux.scala 81:58]
      if (state_r == 4'h9 & (_GEN_515 & state_w == 4'h9 | ~_GEN_515)) begin // @[cache.scala 72:20]
        state <= 4'h5;
      end else begin
        state <= 4'h4;
      end
    end else if (4'h3 == state) begin // @[Mux.scala 81:58]
      state <= 4'h0;
    end else begin
      state <= _state_T_21;
    end
    if (reset) begin // @[cache.scala 41:24]
      state_r <= 4'h0; // @[cache.scala 41:24]
    end else if (4'h9 == state_r) begin // @[Mux.scala 81:58]
      if (state != 4'h4) begin // @[cache.scala 102:20]
        state_r <= 4'h0;
      end else begin
        state_r <= 4'h9;
      end
    end else if (4'h7 == state_r) begin // @[Mux.scala 81:58]
      if (_state_r_T_4) begin // @[cache.scala 101:20]
        state_r <= 4'h9;
      end else begin
        state_r <= 4'h7;
      end
    end else if (4'h6 == state_r) begin // @[Mux.scala 81:58]
      state_r <= _state_r_T_5;
    end else begin
      state_r <= _state_r_T_11;
    end
    if (reset) begin // @[cache.scala 42:24]
      state_w <= 4'h0; // @[cache.scala 42:24]
    end else if (4'h9 == state_w) begin // @[Mux.scala 81:58]
      if (state != 4'h4) begin // @[cache.scala 102:20]
        state_w <= 4'h0;
      end else begin
        state_w <= 4'h9;
      end
    end else if (4'h7 == state_w) begin // @[Mux.scala 81:58]
      if (_state_w_T_6) begin // @[cache.scala 112:20]
        state_w <= 4'h9;
      end else begin
        state_w <= 4'h7;
      end
    end else if (4'h6 == state_w) begin // @[Mux.scala 81:58]
      state_w <= _state_w_T_5;
    end else begin
      state_w <= _state_w_T_13;
    end
    if (reset) begin // @[cache.scala 51:22]
      rmode <= 1'h0; // @[cache.scala 51:22]
    end else begin
      rmode <= state == 4'h0 & _rmode_T_1 | _rmode_T_4; // @[cache.scala 53:9]
    end
    if (reset) begin // @[cache.scala 52:22]
      wmode <= 1'h0; // @[cache.scala 52:22]
    end else begin
      wmode <= _rmode_T & _wmode_T_1 | _wmode_T_4; // @[cache.scala 54:9]
    end
    if (reset) begin // @[cache.scala 138:21]
      rcnt <= 1'h0; // @[cache.scala 138:21]
    end else if (_io_mem_ar_valid_T) begin // @[cache.scala 139:14]
      rcnt <= 1'h0;
    end else if (_state_r_T_4) begin // @[cache.scala 139:43]
      rcnt <= rcnt + 1'h1;
    end
    if (reset) begin // @[cache.scala 150:22]
      taggg <= 42'h0; // @[cache.scala 150:22]
    end else begin
      taggg <= tag_read; // @[cache.scala 151:9]
    end
    if (reset) begin // @[cache.scala 193:18]
      cnt <= 32'h0; // @[cache.scala 193:18]
    end else if (_wdata_T) begin // @[cache.scala 195:11]
      cnt <= _cnt_T_2;
    end
    if (reset) begin // @[cache.scala 194:18]
      hit <= 32'h0; // @[cache.scala 194:18]
    end else if (_io_in_r_bits_data_T) begin // @[cache.scala 196:11]
      hit <= _hit_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_tag[initvar] = _RAND_0[41:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cache_tag_tag_read_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cache_tag_tag_read_MPORT_addr_pipe_0 = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  valid_0_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_0_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_1_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_1_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_2_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_3_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_3_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_4_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_4_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_5_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_5_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_6_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_6_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_7_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_7_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_8_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_8_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_9_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_9_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_10_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_10_1 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_11_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_11_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_12_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_12_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_13_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_13_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_14_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_14_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_15_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_15_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_16_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_16_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_17_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_17_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_18_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_18_1 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_19_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_19_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_20_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_20_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_21_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_21_1 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_22_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_22_1 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_23_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_23_1 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_24_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_24_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_25_0 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_25_1 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_26_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_26_1 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_27_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_27_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_28_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_28_1 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_29_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_29_1 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_30_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_30_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_31_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_31_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_32_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_32_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_33_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_33_1 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_34_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_34_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_35_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_35_1 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_36_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_36_1 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_37_0 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_37_1 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_38_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_38_1 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_39_0 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_39_1 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_40_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_40_1 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_41_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_41_1 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_42_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_42_1 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_43_0 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_43_1 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_44_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_44_1 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_45_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_45_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_46_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_46_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_47_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_47_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_48_0 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_48_1 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_49_0 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_49_1 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_50_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_50_1 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_51_0 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_51_1 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_52_0 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_52_1 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_53_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_53_1 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_54_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_54_1 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_55_0 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_55_1 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_56_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_56_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_57_0 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_57_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_58_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_58_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_59_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_59_1 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_60_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_60_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_61_0 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_61_1 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_62_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_62_1 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_63_0 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_63_1 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_64_0 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_64_1 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_65_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_65_1 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_66_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_66_1 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_67_0 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_67_1 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_68_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_68_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_69_0 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_69_1 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_70_0 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_70_1 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_71_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_71_1 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_72_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_72_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_73_0 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_73_1 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_74_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_74_1 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_75_0 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_75_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_76_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_76_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_77_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_77_1 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_78_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_78_1 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_79_0 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_79_1 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_80_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_80_1 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_81_0 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_81_1 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_82_0 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_82_1 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_83_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_83_1 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_84_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_84_1 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_85_0 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_85_1 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_86_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_86_1 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_87_0 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_87_1 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_88_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_88_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_89_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_89_1 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_90_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_90_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_91_0 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_91_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_92_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_92_1 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_93_0 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_93_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_94_0 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_94_1 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_95_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_95_1 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_96_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_96_1 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_97_0 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_97_1 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_98_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_98_1 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_99_0 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_99_1 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_100_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_100_1 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_101_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_101_1 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_102_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_102_1 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_103_0 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_103_1 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_104_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_104_1 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_105_0 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_105_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_106_0 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_106_1 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_107_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_107_1 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_108_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_108_1 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_109_0 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_109_1 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_110_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_110_1 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_111_0 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_111_1 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_112_0 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_112_1 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_113_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_113_1 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_114_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_114_1 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_115_0 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_115_1 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_116_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_116_1 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_117_0 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_117_1 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_118_0 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_118_1 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_119_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_119_1 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_120_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_120_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_121_0 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_121_1 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_122_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_122_1 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_123_0 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_123_1 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_124_0 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_124_1 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_125_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_125_1 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_126_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_126_1 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_127_0 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_127_1 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  dirty_0_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dirty_0_1 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  dirty_1_0 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  dirty_1_1 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  dirty_2_0 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  dirty_2_1 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  dirty_3_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  dirty_3_1 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  dirty_4_0 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  dirty_4_1 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  dirty_5_0 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  dirty_5_1 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  dirty_6_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  dirty_6_1 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  dirty_7_0 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  dirty_7_1 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  dirty_8_0 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  dirty_8_1 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  dirty_9_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  dirty_9_1 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  dirty_10_0 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  dirty_10_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  dirty_11_0 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  dirty_11_1 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  dirty_12_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  dirty_12_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  dirty_13_0 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  dirty_13_1 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  dirty_14_0 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  dirty_14_1 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  dirty_15_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  dirty_15_1 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  dirty_16_0 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  dirty_16_1 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  dirty_17_0 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  dirty_17_1 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  dirty_18_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  dirty_18_1 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  dirty_19_0 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  dirty_19_1 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  dirty_20_0 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  dirty_20_1 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  dirty_21_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  dirty_21_1 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  dirty_22_0 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  dirty_22_1 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  dirty_23_0 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  dirty_23_1 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  dirty_24_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  dirty_24_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  dirty_25_0 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  dirty_25_1 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  dirty_26_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  dirty_26_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  dirty_27_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  dirty_27_1 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  dirty_28_0 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  dirty_28_1 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  dirty_29_0 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  dirty_29_1 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  dirty_30_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  dirty_30_1 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  dirty_31_0 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  dirty_31_1 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  dirty_32_0 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  dirty_32_1 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  dirty_33_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  dirty_33_1 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  dirty_34_0 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  dirty_34_1 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  dirty_35_0 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  dirty_35_1 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  dirty_36_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  dirty_36_1 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  dirty_37_0 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  dirty_37_1 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  dirty_38_0 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  dirty_38_1 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  dirty_39_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dirty_39_1 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  dirty_40_0 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  dirty_40_1 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  dirty_41_0 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  dirty_41_1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  dirty_42_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  dirty_42_1 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  dirty_43_0 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  dirty_43_1 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  dirty_44_0 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  dirty_44_1 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  dirty_45_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  dirty_45_1 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  dirty_46_0 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  dirty_46_1 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  dirty_47_0 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  dirty_47_1 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  dirty_48_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  dirty_48_1 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  dirty_49_0 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  dirty_49_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  dirty_50_0 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  dirty_50_1 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  dirty_51_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  dirty_51_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  dirty_52_0 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  dirty_52_1 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  dirty_53_0 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  dirty_53_1 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  dirty_54_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  dirty_54_1 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  dirty_55_0 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  dirty_55_1 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  dirty_56_0 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  dirty_56_1 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  dirty_57_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  dirty_57_1 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  dirty_58_0 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  dirty_58_1 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  dirty_59_0 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  dirty_59_1 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  dirty_60_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  dirty_60_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  dirty_61_0 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  dirty_61_1 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  dirty_62_0 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  dirty_62_1 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  dirty_63_0 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  dirty_63_1 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  dirty_64_0 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  dirty_64_1 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  dirty_65_0 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  dirty_65_1 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  dirty_66_0 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  dirty_66_1 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  dirty_67_0 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  dirty_67_1 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  dirty_68_0 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  dirty_68_1 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  dirty_69_0 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  dirty_69_1 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  dirty_70_0 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  dirty_70_1 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  dirty_71_0 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  dirty_71_1 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  dirty_72_0 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  dirty_72_1 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  dirty_73_0 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  dirty_73_1 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  dirty_74_0 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  dirty_74_1 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  dirty_75_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  dirty_75_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  dirty_76_0 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  dirty_76_1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  dirty_77_0 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  dirty_77_1 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  dirty_78_0 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  dirty_78_1 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  dirty_79_0 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  dirty_79_1 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  dirty_80_0 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  dirty_80_1 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  dirty_81_0 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  dirty_81_1 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  dirty_82_0 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  dirty_82_1 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  dirty_83_0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  dirty_83_1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  dirty_84_0 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  dirty_84_1 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  dirty_85_0 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  dirty_85_1 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  dirty_86_0 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  dirty_86_1 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  dirty_87_0 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  dirty_87_1 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  dirty_88_0 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  dirty_88_1 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  dirty_89_0 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  dirty_89_1 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  dirty_90_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  dirty_90_1 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  dirty_91_0 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  dirty_91_1 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  dirty_92_0 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  dirty_92_1 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  dirty_93_0 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  dirty_93_1 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  dirty_94_0 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  dirty_94_1 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  dirty_95_0 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  dirty_95_1 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  dirty_96_0 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  dirty_96_1 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  dirty_97_0 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  dirty_97_1 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  dirty_98_0 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  dirty_98_1 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  dirty_99_0 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  dirty_99_1 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  dirty_100_0 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  dirty_100_1 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  dirty_101_0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  dirty_101_1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  dirty_102_0 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  dirty_102_1 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  dirty_103_0 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  dirty_103_1 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  dirty_104_0 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  dirty_104_1 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  dirty_105_0 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  dirty_105_1 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  dirty_106_0 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  dirty_106_1 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  dirty_107_0 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  dirty_107_1 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  dirty_108_0 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  dirty_108_1 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  dirty_109_0 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  dirty_109_1 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  dirty_110_0 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  dirty_110_1 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  dirty_111_0 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  dirty_111_1 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  dirty_112_0 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  dirty_112_1 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  dirty_113_0 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  dirty_113_1 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  dirty_114_0 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  dirty_114_1 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  dirty_115_0 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  dirty_115_1 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  dirty_116_0 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  dirty_116_1 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  dirty_117_0 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  dirty_117_1 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  dirty_118_0 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  dirty_118_1 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  dirty_119_0 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  dirty_119_1 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  dirty_120_0 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  dirty_120_1 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  dirty_121_0 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  dirty_121_1 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  dirty_122_0 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  dirty_122_1 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  dirty_123_0 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  dirty_123_1 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  dirty_124_0 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  dirty_124_1 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  dirty_125_0 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  dirty_125_1 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  dirty_126_0 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  dirty_126_1 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  dirty_127_0 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  dirty_127_1 = _RAND_514[0:0];
  _RAND_515 = {4{`RANDOM}};
  buf_ = _RAND_515[127:0];
  _RAND_516 = {1{`RANDOM}};
  addr = _RAND_516[31:0];
  _RAND_517 = {4{`RANDOM}};
  wdata = _RAND_517[127:0];
  _RAND_518 = {4{`RANDOM}};
  wstrb = _RAND_518[127:0];
  _RAND_519 = {1{`RANDOM}};
  way2 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  state = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  state_r = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  state_w = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  rmode = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  wmode = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  rcnt = _RAND_525[0:0];
  _RAND_526 = {2{`RANDOM}};
  taggg = _RAND_526[41:0];
  _RAND_527 = {1{`RANDOM}};
  cnt = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  hit = _RAND_528[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheRAM(
  input          clock,
  input          reset,
  output [127:0] io_bits_Q,
  input          io_bits_CEN,
  input          io_bits_WEN,
  input  [127:0] io_bits_BWEN,
  input  [7:0]   io_bits_A,
  input  [127:0] io_bits_D
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] S011HD1P_X32Y2D128_BW_Q; // @[CacheRAM.scala 19:18]
  wire  S011HD1P_X32Y2D128_BW_CLK; // @[CacheRAM.scala 19:18]
  wire  S011HD1P_X32Y2D128_BW_CEN; // @[CacheRAM.scala 19:18]
  wire  S011HD1P_X32Y2D128_BW_WEN; // @[CacheRAM.scala 19:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_BWEN; // @[CacheRAM.scala 19:18]
  wire [5:0] S011HD1P_X32Y2D128_BW_A; // @[CacheRAM.scala 19:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_D; // @[CacheRAM.scala 19:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_1_Q; // @[CacheRAM.scala 20:18]
  wire  S011HD1P_X32Y2D128_BW_1_CLK; // @[CacheRAM.scala 20:18]
  wire  S011HD1P_X32Y2D128_BW_1_CEN; // @[CacheRAM.scala 20:18]
  wire  S011HD1P_X32Y2D128_BW_1_WEN; // @[CacheRAM.scala 20:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_1_BWEN; // @[CacheRAM.scala 20:18]
  wire [5:0] S011HD1P_X32Y2D128_BW_1_A; // @[CacheRAM.scala 20:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_1_D; // @[CacheRAM.scala 20:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_2_Q; // @[CacheRAM.scala 21:18]
  wire  S011HD1P_X32Y2D128_BW_2_CLK; // @[CacheRAM.scala 21:18]
  wire  S011HD1P_X32Y2D128_BW_2_CEN; // @[CacheRAM.scala 21:18]
  wire  S011HD1P_X32Y2D128_BW_2_WEN; // @[CacheRAM.scala 21:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_2_BWEN; // @[CacheRAM.scala 21:18]
  wire [5:0] S011HD1P_X32Y2D128_BW_2_A; // @[CacheRAM.scala 21:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_2_D; // @[CacheRAM.scala 21:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_3_Q; // @[CacheRAM.scala 22:18]
  wire  S011HD1P_X32Y2D128_BW_3_CLK; // @[CacheRAM.scala 22:18]
  wire  S011HD1P_X32Y2D128_BW_3_CEN; // @[CacheRAM.scala 22:18]
  wire  S011HD1P_X32Y2D128_BW_3_WEN; // @[CacheRAM.scala 22:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_3_BWEN; // @[CacheRAM.scala 22:18]
  wire [5:0] S011HD1P_X32Y2D128_BW_3_A; // @[CacheRAM.scala 22:18]
  wire [127:0] S011HD1P_X32Y2D128_BW_3_D; // @[CacheRAM.scala 22:18]
  reg [1:0] choose; // @[CacheRAM.scala 27:23]
  wire [127:0] _io_bits_Q_T_3 = choose == 2'h2 ? S011HD1P_X32Y2D128_BW_2_Q : S011HD1P_X32Y2D128_BW_3_Q; // @[CacheRAM.scala 39:17]
  wire [127:0] _io_bits_Q_T_4 = choose == 2'h1 ? S011HD1P_X32Y2D128_BW_1_Q : _io_bits_Q_T_3; // @[CacheRAM.scala 38:17]
  S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW ( // @[CacheRAM.scala 19:18]
    .Q(S011HD1P_X32Y2D128_BW_Q),
    .CLK(S011HD1P_X32Y2D128_BW_CLK),
    .CEN(S011HD1P_X32Y2D128_BW_CEN),
    .WEN(S011HD1P_X32Y2D128_BW_WEN),
    .BWEN(S011HD1P_X32Y2D128_BW_BWEN),
    .A(S011HD1P_X32Y2D128_BW_A),
    .D(S011HD1P_X32Y2D128_BW_D)
  );
  S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW_1 ( // @[CacheRAM.scala 20:18]
    .Q(S011HD1P_X32Y2D128_BW_1_Q),
    .CLK(S011HD1P_X32Y2D128_BW_1_CLK),
    .CEN(S011HD1P_X32Y2D128_BW_1_CEN),
    .WEN(S011HD1P_X32Y2D128_BW_1_WEN),
    .BWEN(S011HD1P_X32Y2D128_BW_1_BWEN),
    .A(S011HD1P_X32Y2D128_BW_1_A),
    .D(S011HD1P_X32Y2D128_BW_1_D)
  );
  S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW_2 ( // @[CacheRAM.scala 21:18]
    .Q(S011HD1P_X32Y2D128_BW_2_Q),
    .CLK(S011HD1P_X32Y2D128_BW_2_CLK),
    .CEN(S011HD1P_X32Y2D128_BW_2_CEN),
    .WEN(S011HD1P_X32Y2D128_BW_2_WEN),
    .BWEN(S011HD1P_X32Y2D128_BW_2_BWEN),
    .A(S011HD1P_X32Y2D128_BW_2_A),
    .D(S011HD1P_X32Y2D128_BW_2_D)
  );
  S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW_3 ( // @[CacheRAM.scala 22:18]
    .Q(S011HD1P_X32Y2D128_BW_3_Q),
    .CLK(S011HD1P_X32Y2D128_BW_3_CLK),
    .CEN(S011HD1P_X32Y2D128_BW_3_CEN),
    .WEN(S011HD1P_X32Y2D128_BW_3_WEN),
    .BWEN(S011HD1P_X32Y2D128_BW_3_BWEN),
    .A(S011HD1P_X32Y2D128_BW_3_A),
    .D(S011HD1P_X32Y2D128_BW_3_D)
  );
  assign io_bits_Q = choose == 2'h0 ? S011HD1P_X32Y2D128_BW_Q : _io_bits_Q_T_4; // @[CacheRAM.scala 37:17]
  assign S011HD1P_X32Y2D128_BW_CLK = clock; // @[CacheRAM.scala 40:11]
  assign S011HD1P_X32Y2D128_BW_CEN = ~(io_bits_CEN & io_bits_A[7:6] == 2'h0); // @[CacheRAM.scala 41:14]
  assign S011HD1P_X32Y2D128_BW_WEN = ~io_bits_WEN; // @[CacheRAM.scala 42:14]
  assign S011HD1P_X32Y2D128_BW_BWEN = ~io_bits_BWEN; // @[CacheRAM.scala 43:15]
  assign S011HD1P_X32Y2D128_BW_A = io_bits_A[5:0]; // @[CacheRAM.scala 44:21]
  assign S011HD1P_X32Y2D128_BW_D = io_bits_D; // @[CacheRAM.scala 45:9]
  assign S011HD1P_X32Y2D128_BW_1_CLK = clock; // @[CacheRAM.scala 47:11]
  assign S011HD1P_X32Y2D128_BW_1_CEN = ~(io_bits_CEN & io_bits_A[7:6] == 2'h1); // @[CacheRAM.scala 48:14]
  assign S011HD1P_X32Y2D128_BW_1_WEN = ~io_bits_WEN; // @[CacheRAM.scala 49:14]
  assign S011HD1P_X32Y2D128_BW_1_BWEN = ~io_bits_BWEN; // @[CacheRAM.scala 50:15]
  assign S011HD1P_X32Y2D128_BW_1_A = io_bits_A[5:0]; // @[CacheRAM.scala 51:21]
  assign S011HD1P_X32Y2D128_BW_1_D = io_bits_D; // @[CacheRAM.scala 52:9]
  assign S011HD1P_X32Y2D128_BW_2_CLK = clock; // @[CacheRAM.scala 54:11]
  assign S011HD1P_X32Y2D128_BW_2_CEN = ~(io_bits_CEN & io_bits_A[7:6] == 2'h2); // @[CacheRAM.scala 55:14]
  assign S011HD1P_X32Y2D128_BW_2_WEN = ~io_bits_WEN; // @[CacheRAM.scala 56:14]
  assign S011HD1P_X32Y2D128_BW_2_BWEN = ~io_bits_BWEN; // @[CacheRAM.scala 57:15]
  assign S011HD1P_X32Y2D128_BW_2_A = io_bits_A[5:0]; // @[CacheRAM.scala 58:21]
  assign S011HD1P_X32Y2D128_BW_2_D = io_bits_D; // @[CacheRAM.scala 59:9]
  assign S011HD1P_X32Y2D128_BW_3_CLK = clock; // @[CacheRAM.scala 61:11]
  assign S011HD1P_X32Y2D128_BW_3_CEN = ~(io_bits_CEN & io_bits_A[7:6] == 2'h3); // @[CacheRAM.scala 62:14]
  assign S011HD1P_X32Y2D128_BW_3_WEN = ~io_bits_WEN; // @[CacheRAM.scala 63:14]
  assign S011HD1P_X32Y2D128_BW_3_BWEN = ~io_bits_BWEN; // @[CacheRAM.scala 64:15]
  assign S011HD1P_X32Y2D128_BW_3_A = io_bits_A[5:0]; // @[CacheRAM.scala 65:21]
  assign S011HD1P_X32Y2D128_BW_3_D = io_bits_D; // @[CacheRAM.scala 66:9]
  always @(posedge clock) begin
    if (reset) begin // @[CacheRAM.scala 27:23]
      choose <= 2'h0; // @[CacheRAM.scala 27:23]
    end else begin
      choose <= io_bits_A[7:6]; // @[CacheRAM.scala 28:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  choose = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI4Arbiter(
  input         clock,
  input         reset,
  output        io_ifu_ar_ready,
  input         io_ifu_ar_valid,
  input  [31:0] io_ifu_ar_bits_addr,
  input  [7:0]  io_ifu_ar_bits_len,
  input         io_ifu_r_ready,
  output        io_ifu_r_valid,
  output [63:0] io_ifu_r_bits_data,
  output        io_ifu_aw_ready,
  input         io_ifu_aw_valid,
  input  [31:0] io_ifu_aw_bits_addr,
  output        io_ifu_w_ready,
  input         io_ifu_w_valid,
  input  [63:0] io_ifu_w_bits_data,
  input  [7:0]  io_ifu_w_bits_strb,
  input         io_ifu_w_bits_last,
  input         io_ifu_b_ready,
  output        io_ifu_b_valid,
  output        io_lsu_ar_ready,
  input         io_lsu_ar_valid,
  input  [31:0] io_lsu_ar_bits_addr,
  input  [7:0]  io_lsu_ar_bits_len,
  input         io_lsu_r_ready,
  output        io_lsu_r_valid,
  output [63:0] io_lsu_r_bits_data,
  output        io_lsu_aw_ready,
  input         io_lsu_aw_valid,
  input  [31:0] io_lsu_aw_bits_addr,
  output        io_lsu_w_ready,
  input         io_lsu_w_valid,
  input  [63:0] io_lsu_w_bits_data,
  input  [7:0]  io_lsu_w_bits_strb,
  input         io_lsu_w_bits_last,
  input         io_lsu_b_ready,
  output        io_lsu_b_valid,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [31:0] io_out_ar_bits_addr,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [63:0] io_out_r_bits_data,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [31:0] io_out_aw_bits_addr,
  output [2:0]  io_out_aw_bits_size,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output [7:0]  io_out_w_bits_strb,
  output        io_out_w_bits_last,
  input         io_out_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rstate; // @[Arbiter.scala 48:23]
  reg [1:0] wstate; // @[Arbiter.scala 49:23]
  wire [1:0] _rstate_T = io_lsu_ar_valid ? 2'h2 : 2'h0; // @[Arbiter.scala 53:18]
  wire [1:0] _rstate_T_1 = io_ifu_ar_valid ? 2'h1 : _rstate_T; // @[Arbiter.scala 52:18]
  wire  _rstate_T_2 = io_ifu_r_ready & io_ifu_r_valid; // @[Decoupled.scala 52:35]
  wire  _rstate_T_4 = io_lsu_r_ready & io_lsu_r_valid; // @[Decoupled.scala 52:35]
  wire [1:0] _wstate_T = io_lsu_aw_valid ? 2'h2 : 2'h0; // @[Arbiter.scala 59:18]
  wire [1:0] _wstate_T_1 = io_ifu_aw_valid ? 2'h1 : _wstate_T; // @[Arbiter.scala 58:18]
  wire  _wstate_T_2 = io_ifu_b_ready & io_ifu_b_valid; // @[Decoupled.scala 52:35]
  wire  _wstate_T_4 = io_lsu_b_ready & io_lsu_b_valid; // @[Decoupled.scala 52:35]
  reg [31:0] araddr; // @[Arbiter.scala 68:21]
  reg  arvalid; // @[Arbiter.scala 69:22]
  reg  ifu_arready; // @[Arbiter.scala 70:26]
  reg  lsu_arready; // @[Arbiter.scala 71:26]
  reg [63:0] ifu_rdata; // @[Arbiter.scala 72:24]
  reg [63:0] lsu_rdata; // @[Arbiter.scala 73:24]
  reg  ifu_rvalid; // @[Arbiter.scala 76:25]
  reg  lsu_rvalid; // @[Arbiter.scala 77:25]
  reg  rready; // @[Arbiter.scala 78:21]
  reg [31:0] awaddr; // @[Arbiter.scala 79:21]
  reg  awvalid; // @[Arbiter.scala 80:22]
  reg  ifu_awready; // @[Arbiter.scala 81:26]
  reg  lsu_awready; // @[Arbiter.scala 82:26]
  reg [63:0] wdata; // @[Arbiter.scala 83:20]
  reg [7:0] wstrb; // @[Arbiter.scala 84:20]
  reg  wvalid; // @[Arbiter.scala 85:21]
  reg  ifu_wready; // @[Arbiter.scala 86:25]
  reg  lsu_wready; // @[Arbiter.scala 87:25]
  reg  ifu_bvalid; // @[Arbiter.scala 90:25]
  reg  lsu_bvalid; // @[Arbiter.scala 91:25]
  reg [7:0] arlen; // @[Arbiter.scala 94:22]
  reg [2:0] arsize; // @[Arbiter.scala 95:23]
  reg [2:0] awsize; // @[Arbiter.scala 98:23]
  reg  wlast; // @[Arbiter.scala 100:22]
  wire [1:0] _araddr_T_1 = 2'h0 == rstate ? 2'h0 : 2'h1; // @[Mux.scala 81:58]
  wire [1:0] _arvalid_T_3 = 2'h1 == rstate ? {{1'd0}, io_ifu_ar_valid} : _araddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _arvalid_T_5 = 2'h2 == rstate ? {{1'd0}, io_lsu_ar_valid} : _arvalid_T_3; // @[Mux.scala 81:58]
  wire [1:0] _rready_T_3 = 2'h1 == rstate ? {{1'd0}, io_ifu_r_ready} : _araddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _rready_T_5 = 2'h2 == rstate ? {{1'd0}, io_lsu_r_ready} : _rready_T_3; // @[Mux.scala 81:58]
  wire [1:0] _awaddr_T_1 = 2'h0 == wstate ? 2'h0 : 2'h1; // @[Mux.scala 81:58]
  wire [1:0] _awvalid_T_3 = 2'h1 == wstate ? {{1'd0}, io_ifu_aw_valid} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _awvalid_T_5 = 2'h2 == wstate ? {{1'd0}, io_lsu_aw_valid} : _awvalid_T_3; // @[Mux.scala 81:58]
  wire [1:0] _wvalid_T_3 = 2'h1 == wstate ? {{1'd0}, io_ifu_w_valid} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _wvalid_T_5 = 2'h2 == wstate ? {{1'd0}, io_lsu_w_valid} : _wvalid_T_3; // @[Mux.scala 81:58]
  wire [1:0] _awburst_T_3 = 2'h1 == wstate ? 2'h0 : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _wlast_T_3 = 2'h1 == wstate ? {{1'd0}, io_ifu_w_bits_last} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _wlast_T_5 = 2'h2 == wstate ? {{1'd0}, io_lsu_w_bits_last} : _wlast_T_3; // @[Mux.scala 81:58]
  wire [1:0] _ifu_arready_T_3 = 2'h1 == rstate ? {{1'd0}, io_out_ar_ready} : _araddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_arready_T_5 = 2'h2 == rstate ? 2'h0 : _ifu_arready_T_3; // @[Mux.scala 81:58]
  wire [1:0] _ifu_rresp_T_3 = 2'h1 == rstate ? 2'h0 : _araddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_rvalid_T_3 = 2'h1 == rstate ? {{1'd0}, io_out_r_valid} : _araddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_rvalid_T_5 = 2'h2 == rstate ? 2'h0 : _ifu_rvalid_T_3; // @[Mux.scala 81:58]
  wire [1:0] _ifu_awready_T_3 = 2'h1 == wstate ? {{1'd0}, io_out_aw_ready} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_awready_T_5 = 2'h2 == wstate ? 2'h0 : _ifu_awready_T_3; // @[Mux.scala 81:58]
  wire [1:0] _ifu_wready_T_3 = 2'h1 == wstate ? {{1'd0}, io_out_w_ready} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_wready_T_5 = 2'h2 == wstate ? 2'h0 : _ifu_wready_T_3; // @[Mux.scala 81:58]
  wire [1:0] _ifu_bvalid_T_3 = 2'h1 == wstate ? {{1'd0}, io_out_b_valid} : _awaddr_T_1; // @[Mux.scala 81:58]
  wire [1:0] _ifu_bvalid_T_5 = 2'h2 == wstate ? 2'h0 : _ifu_bvalid_T_3; // @[Mux.scala 81:58]
  wire [1:0] _lsu_arready_T_5 = 2'h2 == rstate ? {{1'd0}, io_out_ar_ready} : _ifu_rresp_T_3; // @[Mux.scala 81:58]
  wire [1:0] _lsu_rvalid_T_5 = 2'h2 == rstate ? {{1'd0}, io_out_r_valid} : _ifu_rresp_T_3; // @[Mux.scala 81:58]
  wire [1:0] _lsu_awready_T_5 = 2'h2 == wstate ? {{1'd0}, io_out_aw_ready} : _awburst_T_3; // @[Mux.scala 81:58]
  wire [1:0] _lsu_wready_T_5 = 2'h2 == wstate ? {{1'd0}, io_out_w_ready} : _awburst_T_3; // @[Mux.scala 81:58]
  wire [1:0] _lsu_bvalid_T_5 = 2'h2 == wstate ? {{1'd0}, io_out_b_valid} : _awburst_T_3; // @[Mux.scala 81:58]
  wire [1:0] _GEN_0 = reset ? 2'h0 : _arvalid_T_5; // @[Arbiter.scala 113:10 69:{22,22}]
  wire [1:0] _GEN_1 = reset ? 2'h1 : _ifu_arready_T_5; // @[Arbiter.scala 210:14 70:{26,26}]
  wire [1:0] _GEN_2 = reset ? 2'h0 : _lsu_arready_T_5; // @[Arbiter.scala 266:14 71:{26,26}]
  wire [1:0] _GEN_3 = reset ? 2'h0 : _ifu_rvalid_T_5; // @[Arbiter.scala 228:13 76:{25,25}]
  wire [1:0] _GEN_4 = reset ? 2'h0 : _lsu_rvalid_T_5; // @[Arbiter.scala 284:13 77:{25,25}]
  wire [1:0] _GEN_5 = reset ? 2'h0 : _rready_T_5; // @[Arbiter.scala 78:{21,21} 119:9]
  wire [1:0] _GEN_6 = reset ? 2'h0 : _awvalid_T_5; // @[Arbiter.scala 131:10 80:{22,22}]
  wire [1:0] _GEN_7 = reset ? 2'h0 : _ifu_awready_T_5; // @[Arbiter.scala 234:14 81:{26,26}]
  wire [1:0] _GEN_8 = reset ? 2'h0 : _lsu_awready_T_5; // @[Arbiter.scala 290:14 82:{26,26}]
  wire [1:0] _GEN_9 = reset ? 2'h0 : _wvalid_T_5; // @[Arbiter.scala 85:{21,21} 149:9]
  wire [1:0] _GEN_10 = reset ? 2'h0 : _ifu_wready_T_5; // @[Arbiter.scala 240:13 86:{25,25}]
  wire [1:0] _GEN_11 = reset ? 2'h0 : _lsu_wready_T_5; // @[Arbiter.scala 296:13 87:{25,25}]
  wire [1:0] _GEN_12 = reset ? 2'h0 : _ifu_bvalid_T_5; // @[Arbiter.scala 252:13 90:{25,25}]
  wire [1:0] _GEN_13 = reset ? 2'h0 : _lsu_bvalid_T_5; // @[Arbiter.scala 308:13 91:{25,25}]
  wire [1:0] _GEN_15 = reset ? 2'h0 : _wlast_T_5; // @[Arbiter.scala 100:{22,22} 197:8]
  assign io_ifu_ar_ready = ifu_arready; // @[Arbiter.scala 209:18]
  assign io_ifu_r_valid = ifu_rvalid; // @[Arbiter.scala 227:17]
  assign io_ifu_r_bits_data = ifu_rdata; // @[Arbiter.scala 215:21]
  assign io_ifu_aw_ready = ifu_awready; // @[Arbiter.scala 233:18]
  assign io_ifu_w_ready = ifu_wready; // @[Arbiter.scala 239:17]
  assign io_ifu_b_valid = ifu_bvalid; // @[Arbiter.scala 251:17]
  assign io_lsu_ar_ready = lsu_arready; // @[Arbiter.scala 265:18]
  assign io_lsu_r_valid = lsu_rvalid; // @[Arbiter.scala 283:17]
  assign io_lsu_r_bits_data = lsu_rdata; // @[Arbiter.scala 271:21]
  assign io_lsu_aw_ready = lsu_awready; // @[Arbiter.scala 289:18]
  assign io_lsu_w_ready = lsu_wready; // @[Arbiter.scala 295:17]
  assign io_lsu_b_valid = lsu_bvalid; // @[Arbiter.scala 307:17]
  assign io_out_ar_valid = arvalid; // @[Arbiter.scala 112:18]
  assign io_out_ar_bits_addr = araddr; // @[Arbiter.scala 106:22]
  assign io_out_ar_bits_len = arlen; // @[Arbiter.scala 160:21]
  assign io_out_ar_bits_size = arsize; // @[Arbiter.scala 166:22]
  assign io_out_r_ready = rready; // @[Arbiter.scala 118:17]
  assign io_out_aw_valid = awvalid; // @[Arbiter.scala 130:18]
  assign io_out_aw_bits_addr = awaddr; // @[Arbiter.scala 124:22]
  assign io_out_aw_bits_size = awsize; // @[Arbiter.scala 184:22]
  assign io_out_w_valid = wvalid; // @[Arbiter.scala 148:17]
  assign io_out_w_bits_data = wdata; // @[Arbiter.scala 136:21]
  assign io_out_w_bits_strb = wstrb; // @[Arbiter.scala 142:21]
  assign io_out_w_bits_last = wlast; // @[Arbiter.scala 196:21]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 48:23]
      rstate <= 2'h0; // @[Arbiter.scala 48:23]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      if (_rstate_T_4) begin // @[Arbiter.scala 55:18]
        rstate <= 2'h0;
      end else begin
        rstate <= 2'h2;
      end
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      if (_rstate_T_2) begin // @[Arbiter.scala 54:18]
        rstate <= 2'h0;
      end else begin
        rstate <= 2'h1;
      end
    end else if (2'h0 == rstate) begin // @[Mux.scala 81:58]
      rstate <= _rstate_T_1;
    end else begin
      rstate <= 2'h1;
    end
    if (reset) begin // @[Arbiter.scala 49:23]
      wstate <= 2'h0; // @[Arbiter.scala 49:23]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      if (_wstate_T_4) begin // @[Arbiter.scala 61:18]
        wstate <= 2'h0;
      end else begin
        wstate <= 2'h2;
      end
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      if (_wstate_T_2) begin // @[Arbiter.scala 60:18]
        wstate <= 2'h0;
      end else begin
        wstate <= 2'h1;
      end
    end else if (2'h0 == wstate) begin // @[Mux.scala 81:58]
      wstate <= _wstate_T_1;
    end else begin
      wstate <= 2'h0;
    end
    if (reset) begin // @[Arbiter.scala 68:21]
      araddr <= 32'h0; // @[Arbiter.scala 68:21]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      araddr <= io_lsu_ar_bits_addr;
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      araddr <= io_ifu_ar_bits_addr;
    end else begin
      araddr <= {{30'd0}, _araddr_T_1};
    end
    arvalid <= _GEN_0[0]; // @[Arbiter.scala 113:10 69:{22,22}]
    ifu_arready <= _GEN_1[0]; // @[Arbiter.scala 210:14 70:{26,26}]
    lsu_arready <= _GEN_2[0]; // @[Arbiter.scala 266:14 71:{26,26}]
    if (reset) begin // @[Arbiter.scala 72:24]
      ifu_rdata <= 64'h0; // @[Arbiter.scala 72:24]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      ifu_rdata <= 64'h0;
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      ifu_rdata <= io_out_r_bits_data;
    end else begin
      ifu_rdata <= {{62'd0}, _araddr_T_1};
    end
    if (reset) begin // @[Arbiter.scala 73:24]
      lsu_rdata <= 64'h0; // @[Arbiter.scala 73:24]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      lsu_rdata <= io_out_r_bits_data;
    end else begin
      lsu_rdata <= {{62'd0}, _ifu_rresp_T_3};
    end
    ifu_rvalid <= _GEN_3[0]; // @[Arbiter.scala 228:13 76:{25,25}]
    lsu_rvalid <= _GEN_4[0]; // @[Arbiter.scala 284:13 77:{25,25}]
    rready <= _GEN_5[0]; // @[Arbiter.scala 78:{21,21} 119:9]
    if (reset) begin // @[Arbiter.scala 79:21]
      awaddr <= 32'h0; // @[Arbiter.scala 79:21]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      awaddr <= io_lsu_aw_bits_addr;
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      awaddr <= io_ifu_aw_bits_addr;
    end else begin
      awaddr <= {{30'd0}, _awaddr_T_1};
    end
    awvalid <= _GEN_6[0]; // @[Arbiter.scala 131:10 80:{22,22}]
    ifu_awready <= _GEN_7[0]; // @[Arbiter.scala 234:14 81:{26,26}]
    lsu_awready <= _GEN_8[0]; // @[Arbiter.scala 290:14 82:{26,26}]
    if (reset) begin // @[Arbiter.scala 83:20]
      wdata <= 64'h0; // @[Arbiter.scala 83:20]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      wdata <= io_lsu_w_bits_data;
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      wdata <= io_ifu_w_bits_data;
    end else begin
      wdata <= {{62'd0}, _awaddr_T_1};
    end
    if (reset) begin // @[Arbiter.scala 84:20]
      wstrb <= 8'h0; // @[Arbiter.scala 84:20]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      wstrb <= io_lsu_w_bits_strb;
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      wstrb <= io_ifu_w_bits_strb;
    end else begin
      wstrb <= {{6'd0}, _awaddr_T_1};
    end
    wvalid <= _GEN_9[0]; // @[Arbiter.scala 85:{21,21} 149:9]
    ifu_wready <= _GEN_10[0]; // @[Arbiter.scala 240:13 86:{25,25}]
    lsu_wready <= _GEN_11[0]; // @[Arbiter.scala 296:13 87:{25,25}]
    ifu_bvalid <= _GEN_12[0]; // @[Arbiter.scala 252:13 90:{25,25}]
    lsu_bvalid <= _GEN_13[0]; // @[Arbiter.scala 308:13 91:{25,25}]
    if (reset) begin // @[Arbiter.scala 94:22]
      arlen <= 8'h0; // @[Arbiter.scala 94:22]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      arlen <= io_lsu_ar_bits_len;
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      arlen <= io_ifu_ar_bits_len;
    end else begin
      arlen <= {{6'd0}, _araddr_T_1};
    end
    if (reset) begin // @[Arbiter.scala 95:23]
      arsize <= 3'h0; // @[Arbiter.scala 95:23]
    end else if (2'h2 == rstate) begin // @[Mux.scala 81:58]
      arsize <= 3'h3;
    end else if (2'h1 == rstate) begin // @[Mux.scala 81:58]
      arsize <= 3'h3;
    end else begin
      arsize <= {{1'd0}, _araddr_T_1};
    end
    if (reset) begin // @[Arbiter.scala 98:23]
      awsize <= 3'h0; // @[Arbiter.scala 98:23]
    end else if (2'h2 == wstate) begin // @[Mux.scala 81:58]
      awsize <= 3'h3;
    end else if (2'h1 == wstate) begin // @[Mux.scala 81:58]
      awsize <= 3'h3;
    end else begin
      awsize <= {{1'd0}, _awaddr_T_1};
    end
    wlast <= _GEN_15[0]; // @[Arbiter.scala 100:{22,22} 197:8]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(wstate != 2'h1)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:63 assert(wstate =/= a_ifu)\n"); // @[Arbiter.scala 63:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(wstate != 2'h1)) begin
          $fatal; // @[Arbiter.scala 63:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rstate = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  araddr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  arvalid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_arready = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lsu_arready = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  ifu_rdata = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  lsu_rdata = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  ifu_rvalid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lsu_rvalid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  rready = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  awaddr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  awvalid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ifu_awready = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lsu_awready = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  wstrb = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  wvalid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ifu_wready = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lsu_wready = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ifu_bvalid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lsu_bvalid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  arlen = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  arsize = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  awsize = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  wlast = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXILite2AXI4(
  output        io_in_ar_ready,
  input         io_in_ar_valid,
  input  [31:0] io_in_ar_bits_addr,
  input         io_in_r_ready,
  output        io_in_r_valid,
  output [63:0] io_in_r_bits_data,
  output        io_in_aw_ready,
  input         io_in_aw_valid,
  input  [31:0] io_in_aw_bits_addr,
  output        io_in_w_ready,
  input         io_in_w_valid,
  input  [63:0] io_in_w_bits_data,
  input  [7:0]  io_in_w_bits_strb,
  input         io_in_b_ready,
  output        io_in_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output [7:0]  io_mem_w_bits_strb,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid
);
  assign io_in_ar_ready = io_mem_ar_ready; // @[Crossbar.scala 203:18]
  assign io_in_r_valid = io_mem_r_valid; // @[Crossbar.scala 206:17]
  assign io_in_r_bits_data = io_mem_r_bits_data; // @[Crossbar.scala 204:21]
  assign io_in_aw_ready = io_mem_aw_ready; // @[Crossbar.scala 210:18]
  assign io_in_w_ready = io_mem_w_ready; // @[Crossbar.scala 214:17]
  assign io_in_b_valid = io_mem_b_valid; // @[Crossbar.scala 216:17]
  assign io_mem_ar_valid = io_in_ar_valid; // @[Crossbar.scala 202:18]
  assign io_mem_ar_bits_addr = io_in_ar_bits_addr; // @[Crossbar.scala 201:22]
  assign io_mem_r_ready = io_in_r_ready; // @[Crossbar.scala 207:17]
  assign io_mem_aw_valid = io_in_aw_valid; // @[Crossbar.scala 209:18]
  assign io_mem_aw_bits_addr = io_in_aw_bits_addr; // @[Crossbar.scala 208:22]
  assign io_mem_w_valid = io_in_w_valid; // @[Crossbar.scala 213:17]
  assign io_mem_w_bits_data = io_in_w_bits_data; // @[Crossbar.scala 211:21]
  assign io_mem_w_bits_strb = io_in_w_bits_strb; // @[Crossbar.scala 212:21]
  assign io_mem_w_bits_last = io_in_w_valid; // @[Crossbar.scala 227:22]
  assign io_mem_b_ready = io_in_b_ready; // @[Crossbar.scala 217:17]
endmodule
module Crossbar(
  input          clock,
  input          reset,
  output         io_in1_ar_ready,
  input          io_in1_ar_valid,
  input  [31:0]  io_in1_ar_bits_addr,
  output         io_in1_r_valid,
  output [63:0]  io_in1_r_bits_data,
  output         io_in2_ar_ready,
  input          io_in2_ar_valid,
  input  [31:0]  io_in2_ar_bits_addr,
  input          io_in2_r_ready,
  output         io_in2_r_valid,
  output [63:0]  io_in2_r_bits_data,
  output         io_in2_aw_ready,
  input          io_in2_aw_valid,
  input  [31:0]  io_in2_aw_bits_addr,
  output         io_in2_w_ready,
  input          io_in2_w_valid,
  input  [63:0]  io_in2_w_bits_data,
  input  [7:0]   io_in2_w_bits_strb,
  output         io_in2_b_valid,
  input          io_out_ar_ready,
  output         io_out_ar_valid,
  output [31:0]  io_out_ar_bits_addr,
  output [7:0]   io_out_ar_bits_len,
  output [2:0]   io_out_ar_bits_size,
  output         io_out_r_ready,
  input          io_out_r_valid,
  input  [63:0]  io_out_r_bits_data,
  input          io_out_aw_ready,
  output         io_out_aw_valid,
  output [31:0]  io_out_aw_bits_addr,
  output [2:0]   io_out_aw_bits_size,
  input          io_out_w_ready,
  output         io_out_w_valid,
  output [63:0]  io_out_w_bits_data,
  output [7:0]   io_out_w_bits_strb,
  output         io_out_w_bits_last,
  input          io_out_b_valid,
  output [127:0] io_hitrate
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  Cache_clock; // @[Crossbar.scala 14:22]
  wire  Cache_reset; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_ar_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_ar_valid; // @[Crossbar.scala 14:22]
  wire [31:0] Cache_io_in_ar_bits_addr; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_r_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_r_valid; // @[Crossbar.scala 14:22]
  wire [63:0] Cache_io_in_r_bits_data; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_aw_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_aw_valid; // @[Crossbar.scala 14:22]
  wire [31:0] Cache_io_in_aw_bits_addr; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_w_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_w_valid; // @[Crossbar.scala 14:22]
  wire [63:0] Cache_io_in_w_bits_data; // @[Crossbar.scala 14:22]
  wire [7:0] Cache_io_in_w_bits_strb; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_b_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_in_b_valid; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_ar_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_ar_valid; // @[Crossbar.scala 14:22]
  wire [31:0] Cache_io_mem_ar_bits_addr; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_r_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_r_valid; // @[Crossbar.scala 14:22]
  wire [63:0] Cache_io_mem_r_bits_data; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_aw_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_aw_valid; // @[Crossbar.scala 14:22]
  wire [31:0] Cache_io_mem_aw_bits_addr; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_w_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_w_valid; // @[Crossbar.scala 14:22]
  wire [63:0] Cache_io_mem_w_bits_data; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_w_bits_last; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_b_ready; // @[Crossbar.scala 14:22]
  wire  Cache_io_mem_b_valid; // @[Crossbar.scala 14:22]
  wire [127:0] Cache_io_ram_bits_Q; // @[Crossbar.scala 14:22]
  wire  Cache_io_ram_bits_CEN; // @[Crossbar.scala 14:22]
  wire  Cache_io_ram_bits_WEN; // @[Crossbar.scala 14:22]
  wire [127:0] Cache_io_ram_bits_BWEN; // @[Crossbar.scala 14:22]
  wire [7:0] Cache_io_ram_bits_A; // @[Crossbar.scala 14:22]
  wire [127:0] Cache_io_ram_bits_D; // @[Crossbar.scala 14:22]
  wire [63:0] Cache_io_hitrate; // @[Crossbar.scala 14:22]
  wire  CacheRAM_clock; // @[Crossbar.scala 15:25]
  wire  CacheRAM_reset; // @[Crossbar.scala 15:25]
  wire [127:0] CacheRAM_io_bits_Q; // @[Crossbar.scala 15:25]
  wire  CacheRAM_io_bits_CEN; // @[Crossbar.scala 15:25]
  wire  CacheRAM_io_bits_WEN; // @[Crossbar.scala 15:25]
  wire [127:0] CacheRAM_io_bits_BWEN; // @[Crossbar.scala 15:25]
  wire [7:0] CacheRAM_io_bits_A; // @[Crossbar.scala 15:25]
  wire [127:0] CacheRAM_io_bits_D; // @[Crossbar.scala 15:25]
  wire  Cache_1_clock; // @[Crossbar.scala 16:22]
  wire  Cache_1_reset; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_ar_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_ar_valid; // @[Crossbar.scala 16:22]
  wire [31:0] Cache_1_io_in_ar_bits_addr; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_r_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_r_valid; // @[Crossbar.scala 16:22]
  wire [63:0] Cache_1_io_in_r_bits_data; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_aw_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_aw_valid; // @[Crossbar.scala 16:22]
  wire [31:0] Cache_1_io_in_aw_bits_addr; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_w_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_w_valid; // @[Crossbar.scala 16:22]
  wire [63:0] Cache_1_io_in_w_bits_data; // @[Crossbar.scala 16:22]
  wire [7:0] Cache_1_io_in_w_bits_strb; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_b_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_in_b_valid; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_ar_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_ar_valid; // @[Crossbar.scala 16:22]
  wire [31:0] Cache_1_io_mem_ar_bits_addr; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_r_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_r_valid; // @[Crossbar.scala 16:22]
  wire [63:0] Cache_1_io_mem_r_bits_data; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_aw_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_aw_valid; // @[Crossbar.scala 16:22]
  wire [31:0] Cache_1_io_mem_aw_bits_addr; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_w_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_w_valid; // @[Crossbar.scala 16:22]
  wire [63:0] Cache_1_io_mem_w_bits_data; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_w_bits_last; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_b_ready; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_mem_b_valid; // @[Crossbar.scala 16:22]
  wire [127:0] Cache_1_io_ram_bits_Q; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_ram_bits_CEN; // @[Crossbar.scala 16:22]
  wire  Cache_1_io_ram_bits_WEN; // @[Crossbar.scala 16:22]
  wire [127:0] Cache_1_io_ram_bits_BWEN; // @[Crossbar.scala 16:22]
  wire [7:0] Cache_1_io_ram_bits_A; // @[Crossbar.scala 16:22]
  wire [127:0] Cache_1_io_ram_bits_D; // @[Crossbar.scala 16:22]
  wire [63:0] Cache_1_io_hitrate; // @[Crossbar.scala 16:22]
  wire  CacheRAM_1_clock; // @[Crossbar.scala 17:25]
  wire  CacheRAM_1_reset; // @[Crossbar.scala 17:25]
  wire [127:0] CacheRAM_1_io_bits_Q; // @[Crossbar.scala 17:25]
  wire  CacheRAM_1_io_bits_CEN; // @[Crossbar.scala 17:25]
  wire  CacheRAM_1_io_bits_WEN; // @[Crossbar.scala 17:25]
  wire [127:0] CacheRAM_1_io_bits_BWEN; // @[Crossbar.scala 17:25]
  wire [7:0] CacheRAM_1_io_bits_A; // @[Crossbar.scala 17:25]
  wire [127:0] CacheRAM_1_io_bits_D; // @[Crossbar.scala 17:25]
  wire  AXI4Arbiter_clock; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_reset; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_ar_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_ar_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_ifu_ar_bits_addr; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_ifu_ar_bits_len; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_r_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_r_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_ifu_r_bits_data; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_aw_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_aw_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_ifu_aw_bits_addr; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_w_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_w_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_ifu_w_bits_data; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_ifu_w_bits_strb; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_w_bits_last; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_b_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_ifu_b_valid; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_ar_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_ar_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_lsu_ar_bits_addr; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_lsu_ar_bits_len; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_r_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_r_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_lsu_r_bits_data; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_aw_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_aw_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_lsu_aw_bits_addr; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_w_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_w_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_lsu_w_bits_data; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_lsu_w_bits_strb; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_w_bits_last; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_b_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_lsu_b_valid; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_ar_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_ar_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_out_ar_bits_addr; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_out_ar_bits_len; // @[Crossbar.scala 18:23]
  wire [2:0] AXI4Arbiter_io_out_ar_bits_size; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_r_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_r_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_out_r_bits_data; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_aw_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_aw_valid; // @[Crossbar.scala 18:23]
  wire [31:0] AXI4Arbiter_io_out_aw_bits_addr; // @[Crossbar.scala 18:23]
  wire [2:0] AXI4Arbiter_io_out_aw_bits_size; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_w_ready; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_w_valid; // @[Crossbar.scala 18:23]
  wire [63:0] AXI4Arbiter_io_out_w_bits_data; // @[Crossbar.scala 18:23]
  wire [7:0] AXI4Arbiter_io_out_w_bits_strb; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_w_bits_last; // @[Crossbar.scala 18:23]
  wire  AXI4Arbiter_io_out_b_valid; // @[Crossbar.scala 18:23]
  wire  AXILite2AXI4_io_in_ar_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_ar_valid; // @[Crossbar.scala 19:22]
  wire [31:0] AXILite2AXI4_io_in_ar_bits_addr; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_r_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_r_valid; // @[Crossbar.scala 19:22]
  wire [63:0] AXILite2AXI4_io_in_r_bits_data; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_aw_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_aw_valid; // @[Crossbar.scala 19:22]
  wire [31:0] AXILite2AXI4_io_in_aw_bits_addr; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_w_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_w_valid; // @[Crossbar.scala 19:22]
  wire [63:0] AXILite2AXI4_io_in_w_bits_data; // @[Crossbar.scala 19:22]
  wire [7:0] AXILite2AXI4_io_in_w_bits_strb; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_b_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_in_b_valid; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_ar_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_ar_valid; // @[Crossbar.scala 19:22]
  wire [31:0] AXILite2AXI4_io_mem_ar_bits_addr; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_r_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_r_valid; // @[Crossbar.scala 19:22]
  wire [63:0] AXILite2AXI4_io_mem_r_bits_data; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_aw_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_aw_valid; // @[Crossbar.scala 19:22]
  wire [31:0] AXILite2AXI4_io_mem_aw_bits_addr; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_w_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_w_valid; // @[Crossbar.scala 19:22]
  wire [63:0] AXILite2AXI4_io_mem_w_bits_data; // @[Crossbar.scala 19:22]
  wire [7:0] AXILite2AXI4_io_mem_w_bits_strb; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_w_bits_last; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_b_ready; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_io_mem_b_valid; // @[Crossbar.scala 19:22]
  wire  AXILite2AXI4_1_io_in_ar_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_ar_valid; // @[Crossbar.scala 20:22]
  wire [31:0] AXILite2AXI4_1_io_in_ar_bits_addr; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_r_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_r_valid; // @[Crossbar.scala 20:22]
  wire [63:0] AXILite2AXI4_1_io_in_r_bits_data; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_aw_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_aw_valid; // @[Crossbar.scala 20:22]
  wire [31:0] AXILite2AXI4_1_io_in_aw_bits_addr; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_w_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_w_valid; // @[Crossbar.scala 20:22]
  wire [63:0] AXILite2AXI4_1_io_in_w_bits_data; // @[Crossbar.scala 20:22]
  wire [7:0] AXILite2AXI4_1_io_in_w_bits_strb; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_b_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_in_b_valid; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_ar_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_ar_valid; // @[Crossbar.scala 20:22]
  wire [31:0] AXILite2AXI4_1_io_mem_ar_bits_addr; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_r_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_r_valid; // @[Crossbar.scala 20:22]
  wire [63:0] AXILite2AXI4_1_io_mem_r_bits_data; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_aw_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_aw_valid; // @[Crossbar.scala 20:22]
  wire [31:0] AXILite2AXI4_1_io_mem_aw_bits_addr; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_w_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_w_valid; // @[Crossbar.scala 20:22]
  wire [63:0] AXILite2AXI4_1_io_mem_w_bits_data; // @[Crossbar.scala 20:22]
  wire [7:0] AXILite2AXI4_1_io_mem_w_bits_strb; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_w_bits_last; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_b_ready; // @[Crossbar.scala 20:22]
  wire  AXILite2AXI4_1_io_mem_b_valid; // @[Crossbar.scala 20:22]
  reg [1:0] istate; // @[Crossbar.scala 38:23]
  wire [1:0] _istate_T_3 = ~io_in1_ar_valid ? 2'h0 : 2'h1; // @[Crossbar.scala 40:21]
  wire  _istate_T_4 = AXI4Arbiter_io_ifu_r_ready & AXI4Arbiter_io_ifu_r_valid; // @[Decoupled.scala 52:35]
  wire  _istate_T_6 = Cache_io_in_r_ready & Cache_io_in_r_valid; // @[Decoupled.scala 52:35]
  reg [1:0] dstate; // @[Crossbar.scala 47:23]
  wire [1:0] _dstate_T_6 = ~(io_in2_aw_valid | io_in2_ar_valid) ? 2'h0 : 2'h1; // @[Crossbar.scala 49:21]
  wire  _dstate_T_7 = AXI4Arbiter_io_lsu_r_ready & AXI4Arbiter_io_lsu_r_valid; // @[Decoupled.scala 52:35]
  wire  _dstate_T_8 = AXI4Arbiter_io_lsu_b_ready & AXI4Arbiter_io_lsu_b_valid; // @[Decoupled.scala 52:35]
  wire  _dstate_T_11 = Cache_1_io_in_r_ready & Cache_1_io_in_r_valid; // @[Decoupled.scala 52:35]
  wire  _dstate_T_12 = Cache_1_io_in_b_ready & Cache_1_io_in_b_valid; // @[Decoupled.scala 52:35]
  wire  _T = istate == 2'h1; // @[Crossbar.scala 57:48]
  wire  _T_4 = dstate == 2'h1; // @[Crossbar.scala 67:48]
  wire  _T_8 = istate == 2'h2; // @[Crossbar.scala 77:49]
  wire  _T_12 = dstate == 2'h2; // @[Crossbar.scala 88:49]
  Cache Cache ( // @[Crossbar.scala 14:22]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_ar_ready(Cache_io_in_ar_ready),
    .io_in_ar_valid(Cache_io_in_ar_valid),
    .io_in_ar_bits_addr(Cache_io_in_ar_bits_addr),
    .io_in_r_ready(Cache_io_in_r_ready),
    .io_in_r_valid(Cache_io_in_r_valid),
    .io_in_r_bits_data(Cache_io_in_r_bits_data),
    .io_in_aw_ready(Cache_io_in_aw_ready),
    .io_in_aw_valid(Cache_io_in_aw_valid),
    .io_in_aw_bits_addr(Cache_io_in_aw_bits_addr),
    .io_in_w_ready(Cache_io_in_w_ready),
    .io_in_w_valid(Cache_io_in_w_valid),
    .io_in_w_bits_data(Cache_io_in_w_bits_data),
    .io_in_w_bits_strb(Cache_io_in_w_bits_strb),
    .io_in_b_ready(Cache_io_in_b_ready),
    .io_in_b_valid(Cache_io_in_b_valid),
    .io_mem_ar_ready(Cache_io_mem_ar_ready),
    .io_mem_ar_valid(Cache_io_mem_ar_valid),
    .io_mem_ar_bits_addr(Cache_io_mem_ar_bits_addr),
    .io_mem_r_ready(Cache_io_mem_r_ready),
    .io_mem_r_valid(Cache_io_mem_r_valid),
    .io_mem_r_bits_data(Cache_io_mem_r_bits_data),
    .io_mem_aw_ready(Cache_io_mem_aw_ready),
    .io_mem_aw_valid(Cache_io_mem_aw_valid),
    .io_mem_aw_bits_addr(Cache_io_mem_aw_bits_addr),
    .io_mem_w_ready(Cache_io_mem_w_ready),
    .io_mem_w_valid(Cache_io_mem_w_valid),
    .io_mem_w_bits_data(Cache_io_mem_w_bits_data),
    .io_mem_w_bits_last(Cache_io_mem_w_bits_last),
    .io_mem_b_ready(Cache_io_mem_b_ready),
    .io_mem_b_valid(Cache_io_mem_b_valid),
    .io_ram_bits_Q(Cache_io_ram_bits_Q),
    .io_ram_bits_CEN(Cache_io_ram_bits_CEN),
    .io_ram_bits_WEN(Cache_io_ram_bits_WEN),
    .io_ram_bits_BWEN(Cache_io_ram_bits_BWEN),
    .io_ram_bits_A(Cache_io_ram_bits_A),
    .io_ram_bits_D(Cache_io_ram_bits_D),
    .io_hitrate(Cache_io_hitrate)
  );
  CacheRAM CacheRAM ( // @[Crossbar.scala 15:25]
    .clock(CacheRAM_clock),
    .reset(CacheRAM_reset),
    .io_bits_Q(CacheRAM_io_bits_Q),
    .io_bits_CEN(CacheRAM_io_bits_CEN),
    .io_bits_WEN(CacheRAM_io_bits_WEN),
    .io_bits_BWEN(CacheRAM_io_bits_BWEN),
    .io_bits_A(CacheRAM_io_bits_A),
    .io_bits_D(CacheRAM_io_bits_D)
  );
  Cache Cache_1 ( // @[Crossbar.scala 16:22]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_ar_ready(Cache_1_io_in_ar_ready),
    .io_in_ar_valid(Cache_1_io_in_ar_valid),
    .io_in_ar_bits_addr(Cache_1_io_in_ar_bits_addr),
    .io_in_r_ready(Cache_1_io_in_r_ready),
    .io_in_r_valid(Cache_1_io_in_r_valid),
    .io_in_r_bits_data(Cache_1_io_in_r_bits_data),
    .io_in_aw_ready(Cache_1_io_in_aw_ready),
    .io_in_aw_valid(Cache_1_io_in_aw_valid),
    .io_in_aw_bits_addr(Cache_1_io_in_aw_bits_addr),
    .io_in_w_ready(Cache_1_io_in_w_ready),
    .io_in_w_valid(Cache_1_io_in_w_valid),
    .io_in_w_bits_data(Cache_1_io_in_w_bits_data),
    .io_in_w_bits_strb(Cache_1_io_in_w_bits_strb),
    .io_in_b_ready(Cache_1_io_in_b_ready),
    .io_in_b_valid(Cache_1_io_in_b_valid),
    .io_mem_ar_ready(Cache_1_io_mem_ar_ready),
    .io_mem_ar_valid(Cache_1_io_mem_ar_valid),
    .io_mem_ar_bits_addr(Cache_1_io_mem_ar_bits_addr),
    .io_mem_r_ready(Cache_1_io_mem_r_ready),
    .io_mem_r_valid(Cache_1_io_mem_r_valid),
    .io_mem_r_bits_data(Cache_1_io_mem_r_bits_data),
    .io_mem_aw_ready(Cache_1_io_mem_aw_ready),
    .io_mem_aw_valid(Cache_1_io_mem_aw_valid),
    .io_mem_aw_bits_addr(Cache_1_io_mem_aw_bits_addr),
    .io_mem_w_ready(Cache_1_io_mem_w_ready),
    .io_mem_w_valid(Cache_1_io_mem_w_valid),
    .io_mem_w_bits_data(Cache_1_io_mem_w_bits_data),
    .io_mem_w_bits_last(Cache_1_io_mem_w_bits_last),
    .io_mem_b_ready(Cache_1_io_mem_b_ready),
    .io_mem_b_valid(Cache_1_io_mem_b_valid),
    .io_ram_bits_Q(Cache_1_io_ram_bits_Q),
    .io_ram_bits_CEN(Cache_1_io_ram_bits_CEN),
    .io_ram_bits_WEN(Cache_1_io_ram_bits_WEN),
    .io_ram_bits_BWEN(Cache_1_io_ram_bits_BWEN),
    .io_ram_bits_A(Cache_1_io_ram_bits_A),
    .io_ram_bits_D(Cache_1_io_ram_bits_D),
    .io_hitrate(Cache_1_io_hitrate)
  );
  CacheRAM CacheRAM_1 ( // @[Crossbar.scala 17:25]
    .clock(CacheRAM_1_clock),
    .reset(CacheRAM_1_reset),
    .io_bits_Q(CacheRAM_1_io_bits_Q),
    .io_bits_CEN(CacheRAM_1_io_bits_CEN),
    .io_bits_WEN(CacheRAM_1_io_bits_WEN),
    .io_bits_BWEN(CacheRAM_1_io_bits_BWEN),
    .io_bits_A(CacheRAM_1_io_bits_A),
    .io_bits_D(CacheRAM_1_io_bits_D)
  );
  AXI4Arbiter AXI4Arbiter ( // @[Crossbar.scala 18:23]
    .clock(AXI4Arbiter_clock),
    .reset(AXI4Arbiter_reset),
    .io_ifu_ar_ready(AXI4Arbiter_io_ifu_ar_ready),
    .io_ifu_ar_valid(AXI4Arbiter_io_ifu_ar_valid),
    .io_ifu_ar_bits_addr(AXI4Arbiter_io_ifu_ar_bits_addr),
    .io_ifu_ar_bits_len(AXI4Arbiter_io_ifu_ar_bits_len),
    .io_ifu_r_ready(AXI4Arbiter_io_ifu_r_ready),
    .io_ifu_r_valid(AXI4Arbiter_io_ifu_r_valid),
    .io_ifu_r_bits_data(AXI4Arbiter_io_ifu_r_bits_data),
    .io_ifu_aw_ready(AXI4Arbiter_io_ifu_aw_ready),
    .io_ifu_aw_valid(AXI4Arbiter_io_ifu_aw_valid),
    .io_ifu_aw_bits_addr(AXI4Arbiter_io_ifu_aw_bits_addr),
    .io_ifu_w_ready(AXI4Arbiter_io_ifu_w_ready),
    .io_ifu_w_valid(AXI4Arbiter_io_ifu_w_valid),
    .io_ifu_w_bits_data(AXI4Arbiter_io_ifu_w_bits_data),
    .io_ifu_w_bits_strb(AXI4Arbiter_io_ifu_w_bits_strb),
    .io_ifu_w_bits_last(AXI4Arbiter_io_ifu_w_bits_last),
    .io_ifu_b_ready(AXI4Arbiter_io_ifu_b_ready),
    .io_ifu_b_valid(AXI4Arbiter_io_ifu_b_valid),
    .io_lsu_ar_ready(AXI4Arbiter_io_lsu_ar_ready),
    .io_lsu_ar_valid(AXI4Arbiter_io_lsu_ar_valid),
    .io_lsu_ar_bits_addr(AXI4Arbiter_io_lsu_ar_bits_addr),
    .io_lsu_ar_bits_len(AXI4Arbiter_io_lsu_ar_bits_len),
    .io_lsu_r_ready(AXI4Arbiter_io_lsu_r_ready),
    .io_lsu_r_valid(AXI4Arbiter_io_lsu_r_valid),
    .io_lsu_r_bits_data(AXI4Arbiter_io_lsu_r_bits_data),
    .io_lsu_aw_ready(AXI4Arbiter_io_lsu_aw_ready),
    .io_lsu_aw_valid(AXI4Arbiter_io_lsu_aw_valid),
    .io_lsu_aw_bits_addr(AXI4Arbiter_io_lsu_aw_bits_addr),
    .io_lsu_w_ready(AXI4Arbiter_io_lsu_w_ready),
    .io_lsu_w_valid(AXI4Arbiter_io_lsu_w_valid),
    .io_lsu_w_bits_data(AXI4Arbiter_io_lsu_w_bits_data),
    .io_lsu_w_bits_strb(AXI4Arbiter_io_lsu_w_bits_strb),
    .io_lsu_w_bits_last(AXI4Arbiter_io_lsu_w_bits_last),
    .io_lsu_b_ready(AXI4Arbiter_io_lsu_b_ready),
    .io_lsu_b_valid(AXI4Arbiter_io_lsu_b_valid),
    .io_out_ar_ready(AXI4Arbiter_io_out_ar_ready),
    .io_out_ar_valid(AXI4Arbiter_io_out_ar_valid),
    .io_out_ar_bits_addr(AXI4Arbiter_io_out_ar_bits_addr),
    .io_out_ar_bits_len(AXI4Arbiter_io_out_ar_bits_len),
    .io_out_ar_bits_size(AXI4Arbiter_io_out_ar_bits_size),
    .io_out_r_ready(AXI4Arbiter_io_out_r_ready),
    .io_out_r_valid(AXI4Arbiter_io_out_r_valid),
    .io_out_r_bits_data(AXI4Arbiter_io_out_r_bits_data),
    .io_out_aw_ready(AXI4Arbiter_io_out_aw_ready),
    .io_out_aw_valid(AXI4Arbiter_io_out_aw_valid),
    .io_out_aw_bits_addr(AXI4Arbiter_io_out_aw_bits_addr),
    .io_out_aw_bits_size(AXI4Arbiter_io_out_aw_bits_size),
    .io_out_w_ready(AXI4Arbiter_io_out_w_ready),
    .io_out_w_valid(AXI4Arbiter_io_out_w_valid),
    .io_out_w_bits_data(AXI4Arbiter_io_out_w_bits_data),
    .io_out_w_bits_strb(AXI4Arbiter_io_out_w_bits_strb),
    .io_out_w_bits_last(AXI4Arbiter_io_out_w_bits_last),
    .io_out_b_valid(AXI4Arbiter_io_out_b_valid)
  );
  AXILite2AXI4 AXILite2AXI4 ( // @[Crossbar.scala 19:22]
    .io_in_ar_ready(AXILite2AXI4_io_in_ar_ready),
    .io_in_ar_valid(AXILite2AXI4_io_in_ar_valid),
    .io_in_ar_bits_addr(AXILite2AXI4_io_in_ar_bits_addr),
    .io_in_r_ready(AXILite2AXI4_io_in_r_ready),
    .io_in_r_valid(AXILite2AXI4_io_in_r_valid),
    .io_in_r_bits_data(AXILite2AXI4_io_in_r_bits_data),
    .io_in_aw_ready(AXILite2AXI4_io_in_aw_ready),
    .io_in_aw_valid(AXILite2AXI4_io_in_aw_valid),
    .io_in_aw_bits_addr(AXILite2AXI4_io_in_aw_bits_addr),
    .io_in_w_ready(AXILite2AXI4_io_in_w_ready),
    .io_in_w_valid(AXILite2AXI4_io_in_w_valid),
    .io_in_w_bits_data(AXILite2AXI4_io_in_w_bits_data),
    .io_in_w_bits_strb(AXILite2AXI4_io_in_w_bits_strb),
    .io_in_b_ready(AXILite2AXI4_io_in_b_ready),
    .io_in_b_valid(AXILite2AXI4_io_in_b_valid),
    .io_mem_ar_ready(AXILite2AXI4_io_mem_ar_ready),
    .io_mem_ar_valid(AXILite2AXI4_io_mem_ar_valid),
    .io_mem_ar_bits_addr(AXILite2AXI4_io_mem_ar_bits_addr),
    .io_mem_r_ready(AXILite2AXI4_io_mem_r_ready),
    .io_mem_r_valid(AXILite2AXI4_io_mem_r_valid),
    .io_mem_r_bits_data(AXILite2AXI4_io_mem_r_bits_data),
    .io_mem_aw_ready(AXILite2AXI4_io_mem_aw_ready),
    .io_mem_aw_valid(AXILite2AXI4_io_mem_aw_valid),
    .io_mem_aw_bits_addr(AXILite2AXI4_io_mem_aw_bits_addr),
    .io_mem_w_ready(AXILite2AXI4_io_mem_w_ready),
    .io_mem_w_valid(AXILite2AXI4_io_mem_w_valid),
    .io_mem_w_bits_data(AXILite2AXI4_io_mem_w_bits_data),
    .io_mem_w_bits_strb(AXILite2AXI4_io_mem_w_bits_strb),
    .io_mem_w_bits_last(AXILite2AXI4_io_mem_w_bits_last),
    .io_mem_b_ready(AXILite2AXI4_io_mem_b_ready),
    .io_mem_b_valid(AXILite2AXI4_io_mem_b_valid)
  );
  AXILite2AXI4 AXILite2AXI4_1 ( // @[Crossbar.scala 20:22]
    .io_in_ar_ready(AXILite2AXI4_1_io_in_ar_ready),
    .io_in_ar_valid(AXILite2AXI4_1_io_in_ar_valid),
    .io_in_ar_bits_addr(AXILite2AXI4_1_io_in_ar_bits_addr),
    .io_in_r_ready(AXILite2AXI4_1_io_in_r_ready),
    .io_in_r_valid(AXILite2AXI4_1_io_in_r_valid),
    .io_in_r_bits_data(AXILite2AXI4_1_io_in_r_bits_data),
    .io_in_aw_ready(AXILite2AXI4_1_io_in_aw_ready),
    .io_in_aw_valid(AXILite2AXI4_1_io_in_aw_valid),
    .io_in_aw_bits_addr(AXILite2AXI4_1_io_in_aw_bits_addr),
    .io_in_w_ready(AXILite2AXI4_1_io_in_w_ready),
    .io_in_w_valid(AXILite2AXI4_1_io_in_w_valid),
    .io_in_w_bits_data(AXILite2AXI4_1_io_in_w_bits_data),
    .io_in_w_bits_strb(AXILite2AXI4_1_io_in_w_bits_strb),
    .io_in_b_ready(AXILite2AXI4_1_io_in_b_ready),
    .io_in_b_valid(AXILite2AXI4_1_io_in_b_valid),
    .io_mem_ar_ready(AXILite2AXI4_1_io_mem_ar_ready),
    .io_mem_ar_valid(AXILite2AXI4_1_io_mem_ar_valid),
    .io_mem_ar_bits_addr(AXILite2AXI4_1_io_mem_ar_bits_addr),
    .io_mem_r_ready(AXILite2AXI4_1_io_mem_r_ready),
    .io_mem_r_valid(AXILite2AXI4_1_io_mem_r_valid),
    .io_mem_r_bits_data(AXILite2AXI4_1_io_mem_r_bits_data),
    .io_mem_aw_ready(AXILite2AXI4_1_io_mem_aw_ready),
    .io_mem_aw_valid(AXILite2AXI4_1_io_mem_aw_valid),
    .io_mem_aw_bits_addr(AXILite2AXI4_1_io_mem_aw_bits_addr),
    .io_mem_w_ready(AXILite2AXI4_1_io_mem_w_ready),
    .io_mem_w_valid(AXILite2AXI4_1_io_mem_w_valid),
    .io_mem_w_bits_data(AXILite2AXI4_1_io_mem_w_bits_data),
    .io_mem_w_bits_strb(AXILite2AXI4_1_io_mem_w_bits_strb),
    .io_mem_w_bits_last(AXILite2AXI4_1_io_mem_w_bits_last),
    .io_mem_b_ready(AXILite2AXI4_1_io_mem_b_ready),
    .io_mem_b_valid(AXILite2AXI4_1_io_mem_b_valid)
  );
  assign io_in1_ar_ready = _T_8 ? Cache_io_in_ar_ready : AXILite2AXI4_1_io_in_ar_ready; // @[Crossbar.scala 98:23]
  assign io_in1_r_valid = _T_8 ? Cache_io_in_r_valid : AXILite2AXI4_1_io_in_r_valid; // @[Crossbar.scala 99:22]
  assign io_in1_r_bits_data = _T_8 ? Cache_io_in_r_bits_data : AXILite2AXI4_1_io_in_r_bits_data; // @[Crossbar.scala 103:26]
  assign io_in2_ar_ready = _T_12 ? Cache_1_io_in_ar_ready : AXILite2AXI4_io_in_ar_ready; // @[Crossbar.scala 108:23]
  assign io_in2_r_valid = _T_12 ? Cache_1_io_in_r_valid : AXILite2AXI4_io_in_r_valid; // @[Crossbar.scala 109:22]
  assign io_in2_r_bits_data = _T_12 ? Cache_1_io_in_r_bits_data : AXILite2AXI4_io_in_r_bits_data; // @[Crossbar.scala 113:26]
  assign io_in2_aw_ready = _T_12 ? Cache_1_io_in_aw_ready : AXILite2AXI4_io_in_aw_ready; // @[Crossbar.scala 110:23]
  assign io_in2_w_ready = _T_12 | AXILite2AXI4_io_in_w_ready; // @[Crossbar.scala 111:22]
  assign io_in2_b_valid = _T_12 ? Cache_1_io_in_b_valid : AXILite2AXI4_io_in_b_valid; // @[Crossbar.scala 112:22]
  assign io_out_ar_valid = AXI4Arbiter_io_out_ar_valid; // @[Crossbar.scala 35:11]
  assign io_out_ar_bits_addr = AXI4Arbiter_io_out_ar_bits_addr; // @[Crossbar.scala 35:11]
  assign io_out_ar_bits_len = AXI4Arbiter_io_out_ar_bits_len; // @[Crossbar.scala 35:11]
  assign io_out_ar_bits_size = AXI4Arbiter_io_out_ar_bits_size; // @[Crossbar.scala 35:11]
  assign io_out_r_ready = AXI4Arbiter_io_out_r_ready; // @[Crossbar.scala 35:11]
  assign io_out_aw_valid = AXI4Arbiter_io_out_aw_valid; // @[Crossbar.scala 35:11]
  assign io_out_aw_bits_addr = AXI4Arbiter_io_out_aw_bits_addr; // @[Crossbar.scala 35:11]
  assign io_out_aw_bits_size = AXI4Arbiter_io_out_aw_bits_size; // @[Crossbar.scala 35:11]
  assign io_out_w_valid = AXI4Arbiter_io_out_w_valid; // @[Crossbar.scala 35:11]
  assign io_out_w_bits_data = AXI4Arbiter_io_out_w_bits_data; // @[Crossbar.scala 35:11]
  assign io_out_w_bits_strb = AXI4Arbiter_io_out_w_bits_strb; // @[Crossbar.scala 35:11]
  assign io_out_w_bits_last = AXI4Arbiter_io_out_w_bits_last; // @[Crossbar.scala 35:11]
  assign io_hitrate = {Cache_io_hitrate,Cache_1_io_hitrate}; // @[Cat.scala 33:92]
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_ar_valid = io_in1_ar_valid & istate == 2'h2; // @[Crossbar.scala 77:39]
  assign Cache_io_in_ar_bits_addr = io_in1_ar_bits_addr; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_r_ready = 1'h1; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_aw_valid = 1'h0; // @[Crossbar.scala 80:39]
  assign Cache_io_in_aw_bits_addr = 32'h0; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_w_valid = 1'h0; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_w_bits_data = 64'h0; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_w_bits_strb = 8'h0; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_in_b_ready = 1'h0; // @[Crossbar.scala 22:18 27:11]
  assign Cache_io_mem_ar_ready = AXI4Arbiter_io_ifu_ar_ready & _T_8; // @[Crossbar.scala 174:47]
  assign Cache_io_mem_r_valid = AXI4Arbiter_io_ifu_r_valid; // @[Crossbar.scala 175:23]
  assign Cache_io_mem_r_bits_data = AXI4Arbiter_io_ifu_r_bits_data; // @[Crossbar.scala 179:27]
  assign Cache_io_mem_aw_ready = AXI4Arbiter_io_ifu_aw_ready & _T_8; // @[Crossbar.scala 176:47]
  assign Cache_io_mem_w_ready = AXI4Arbiter_io_ifu_w_ready; // @[Crossbar.scala 177:23]
  assign Cache_io_mem_b_valid = AXI4Arbiter_io_ifu_b_valid; // @[Crossbar.scala 178:23]
  assign Cache_io_ram_bits_Q = CacheRAM_io_bits_Q; // @[Crossbar.scala 28:15]
  assign CacheRAM_clock = clock;
  assign CacheRAM_reset = reset;
  assign CacheRAM_io_bits_CEN = Cache_io_ram_bits_CEN; // @[Crossbar.scala 28:15]
  assign CacheRAM_io_bits_WEN = Cache_io_ram_bits_WEN; // @[Crossbar.scala 28:15]
  assign CacheRAM_io_bits_BWEN = Cache_io_ram_bits_BWEN; // @[Crossbar.scala 28:15]
  assign CacheRAM_io_bits_A = Cache_io_ram_bits_A; // @[Crossbar.scala 28:15]
  assign CacheRAM_io_bits_D = Cache_io_ram_bits_D; // @[Crossbar.scala 28:15]
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_ar_valid = io_in2_ar_valid & dstate == 2'h2; // @[Crossbar.scala 88:39]
  assign Cache_1_io_in_ar_bits_addr = io_in2_ar_bits_addr; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_r_ready = io_in2_r_ready; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_aw_valid = io_in2_aw_valid & _T_12; // @[Crossbar.scala 91:39]
  assign Cache_1_io_in_aw_bits_addr = io_in2_aw_bits_addr; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_w_valid = io_in2_w_valid; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_w_bits_data = io_in2_w_bits_data; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_w_bits_strb = io_in2_w_bits_strb; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_in_b_ready = 1'h1; // @[Crossbar.scala 23:18 32:11]
  assign Cache_1_io_mem_ar_ready = AXI4Arbiter_io_lsu_ar_ready & _T_12; // @[Crossbar.scala 185:47]
  assign Cache_1_io_mem_r_valid = AXI4Arbiter_io_lsu_r_valid; // @[Crossbar.scala 186:23]
  assign Cache_1_io_mem_r_bits_data = AXI4Arbiter_io_lsu_r_bits_data; // @[Crossbar.scala 190:27]
  assign Cache_1_io_mem_aw_ready = AXI4Arbiter_io_lsu_aw_ready & _T_12; // @[Crossbar.scala 187:47]
  assign Cache_1_io_mem_w_ready = AXI4Arbiter_io_lsu_w_ready; // @[Crossbar.scala 188:23]
  assign Cache_1_io_mem_b_valid = AXI4Arbiter_io_lsu_b_valid; // @[Crossbar.scala 189:23]
  assign Cache_1_io_ram_bits_Q = CacheRAM_1_io_bits_Q; // @[Crossbar.scala 33:15]
  assign CacheRAM_1_clock = clock;
  assign CacheRAM_1_reset = reset;
  assign CacheRAM_1_io_bits_CEN = Cache_1_io_ram_bits_CEN; // @[Crossbar.scala 33:15]
  assign CacheRAM_1_io_bits_WEN = Cache_1_io_ram_bits_WEN; // @[Crossbar.scala 33:15]
  assign CacheRAM_1_io_bits_BWEN = Cache_1_io_ram_bits_BWEN; // @[Crossbar.scala 33:15]
  assign CacheRAM_1_io_bits_A = Cache_1_io_ram_bits_A; // @[Crossbar.scala 33:15]
  assign CacheRAM_1_io_bits_D = Cache_1_io_ram_bits_D; // @[Crossbar.scala 33:15]
  assign AXI4Arbiter_clock = clock;
  assign AXI4Arbiter_reset = reset;
  assign AXI4Arbiter_io_ifu_ar_valid = _T ? AXILite2AXI4_1_io_mem_ar_valid : Cache_io_mem_ar_valid; // @[Crossbar.scala 117:30]
  assign AXI4Arbiter_io_ifu_ar_bits_addr = _T ? AXILite2AXI4_1_io_mem_ar_bits_addr : Cache_io_mem_ar_bits_addr; // @[Crossbar.scala 118:34]
  assign AXI4Arbiter_io_ifu_ar_bits_len = _T ? 8'h0 : 8'h1; // @[Crossbar.scala 119:33]
  assign AXI4Arbiter_io_ifu_r_ready = _T ? AXILite2AXI4_1_io_mem_r_ready : 1'h1; // @[Crossbar.scala 122:29]
  assign AXI4Arbiter_io_ifu_aw_valid = _T ? AXILite2AXI4_1_io_mem_aw_valid : Cache_io_mem_aw_valid; // @[Crossbar.scala 123:30]
  assign AXI4Arbiter_io_ifu_aw_bits_addr = _T ? AXILite2AXI4_1_io_mem_aw_bits_addr : Cache_io_mem_aw_bits_addr; // @[Crossbar.scala 124:34]
  assign AXI4Arbiter_io_ifu_w_valid = _T ? AXILite2AXI4_1_io_mem_w_valid : Cache_io_mem_w_valid; // @[Crossbar.scala 128:29]
  assign AXI4Arbiter_io_ifu_w_bits_data = _T ? AXILite2AXI4_1_io_mem_w_bits_data : Cache_io_mem_w_bits_data; // @[Crossbar.scala 129:33]
  assign AXI4Arbiter_io_ifu_w_bits_strb = _T ? AXILite2AXI4_1_io_mem_w_bits_strb : 8'hff; // @[Crossbar.scala 130:33]
  assign AXI4Arbiter_io_ifu_w_bits_last = _T ? AXILite2AXI4_1_io_mem_w_bits_last : Cache_io_mem_w_bits_last; // @[Crossbar.scala 131:33]
  assign AXI4Arbiter_io_ifu_b_ready = _T ? AXILite2AXI4_1_io_mem_b_ready : 1'h1; // @[Crossbar.scala 132:29]
  assign AXI4Arbiter_io_lsu_ar_valid = _T_4 ? AXILite2AXI4_io_mem_ar_valid : Cache_1_io_mem_ar_valid; // @[Crossbar.scala 136:30]
  assign AXI4Arbiter_io_lsu_ar_bits_addr = _T_4 ? AXILite2AXI4_io_mem_ar_bits_addr : Cache_1_io_mem_ar_bits_addr; // @[Crossbar.scala 137:34]
  assign AXI4Arbiter_io_lsu_ar_bits_len = _T_4 ? 8'h0 : 8'h1; // @[Crossbar.scala 138:33]
  assign AXI4Arbiter_io_lsu_r_ready = _T_4 ? AXILite2AXI4_io_mem_r_ready : 1'h1; // @[Crossbar.scala 141:29]
  assign AXI4Arbiter_io_lsu_aw_valid = _T_4 ? AXILite2AXI4_io_mem_aw_valid : Cache_1_io_mem_aw_valid; // @[Crossbar.scala 142:30]
  assign AXI4Arbiter_io_lsu_aw_bits_addr = _T_4 ? AXILite2AXI4_io_mem_aw_bits_addr : Cache_1_io_mem_aw_bits_addr; // @[Crossbar.scala 143:34]
  assign AXI4Arbiter_io_lsu_w_valid = _T_4 ? AXILite2AXI4_io_mem_w_valid : Cache_1_io_mem_w_valid; // @[Crossbar.scala 147:29]
  assign AXI4Arbiter_io_lsu_w_bits_data = _T_4 ? AXILite2AXI4_io_mem_w_bits_data : Cache_1_io_mem_w_bits_data; // @[Crossbar.scala 148:33]
  assign AXI4Arbiter_io_lsu_w_bits_strb = _T_4 ? AXILite2AXI4_io_mem_w_bits_strb : 8'hff; // @[Crossbar.scala 149:33]
  assign AXI4Arbiter_io_lsu_w_bits_last = _T_4 ? AXILite2AXI4_io_mem_w_bits_last : Cache_1_io_mem_w_bits_last; // @[Crossbar.scala 150:33]
  assign AXI4Arbiter_io_lsu_b_ready = _T_4 ? AXILite2AXI4_io_mem_b_ready : 1'h1; // @[Crossbar.scala 151:29]
  assign AXI4Arbiter_io_out_ar_ready = io_out_ar_ready; // @[Crossbar.scala 35:11]
  assign AXI4Arbiter_io_out_r_valid = io_out_r_valid; // @[Crossbar.scala 35:11]
  assign AXI4Arbiter_io_out_r_bits_data = io_out_r_bits_data; // @[Crossbar.scala 35:11]
  assign AXI4Arbiter_io_out_aw_ready = io_out_aw_ready; // @[Crossbar.scala 35:11]
  assign AXI4Arbiter_io_out_w_ready = io_out_w_ready; // @[Crossbar.scala 35:11]
  assign AXI4Arbiter_io_out_b_valid = io_out_b_valid; // @[Crossbar.scala 35:11]
  assign AXILite2AXI4_io_in_ar_valid = io_in2_ar_valid & dstate == 2'h1; // @[Crossbar.scala 67:39]
  assign AXILite2AXI4_io_in_ar_bits_addr = io_in2_ar_bits_addr; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_r_ready = io_in2_r_ready; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_aw_valid = io_in2_aw_valid & _T_4; // @[Crossbar.scala 70:39]
  assign AXILite2AXI4_io_in_aw_bits_addr = io_in2_aw_bits_addr; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_w_valid = io_in2_w_valid; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_w_bits_data = io_in2_w_bits_data; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_w_bits_strb = io_in2_w_bits_strb; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_in_b_ready = 1'h1; // @[Crossbar.scala 23:18 32:11]
  assign AXILite2AXI4_io_mem_ar_ready = AXI4Arbiter_io_lsu_ar_ready & _T_4; // @[Crossbar.scala 164:47]
  assign AXILite2AXI4_io_mem_r_valid = AXI4Arbiter_io_lsu_r_valid; // @[Crossbar.scala 165:23]
  assign AXILite2AXI4_io_mem_r_bits_data = AXI4Arbiter_io_lsu_r_bits_data; // @[Crossbar.scala 169:27]
  assign AXILite2AXI4_io_mem_aw_ready = AXI4Arbiter_io_lsu_aw_ready & _T_4; // @[Crossbar.scala 166:47]
  assign AXILite2AXI4_io_mem_w_ready = AXI4Arbiter_io_lsu_w_ready; // @[Crossbar.scala 167:23]
  assign AXILite2AXI4_io_mem_b_valid = AXI4Arbiter_io_lsu_b_valid; // @[Crossbar.scala 168:23]
  assign AXILite2AXI4_1_io_in_ar_valid = io_in1_ar_valid & istate == 2'h1; // @[Crossbar.scala 57:39]
  assign AXILite2AXI4_1_io_in_ar_bits_addr = io_in1_ar_bits_addr; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_r_ready = 1'h1; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_aw_valid = 1'h0; // @[Crossbar.scala 60:39]
  assign AXILite2AXI4_1_io_in_aw_bits_addr = 32'h0; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_w_valid = 1'h0; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_w_bits_data = 64'h0; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_w_bits_strb = 8'h0; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_in_b_ready = 1'h0; // @[Crossbar.scala 22:18 27:11]
  assign AXILite2AXI4_1_io_mem_ar_ready = AXI4Arbiter_io_ifu_ar_ready & _T; // @[Crossbar.scala 153:47]
  assign AXILite2AXI4_1_io_mem_r_valid = AXI4Arbiter_io_ifu_r_valid; // @[Crossbar.scala 154:23]
  assign AXILite2AXI4_1_io_mem_r_bits_data = AXI4Arbiter_io_ifu_r_bits_data; // @[Crossbar.scala 158:27]
  assign AXILite2AXI4_1_io_mem_aw_ready = AXI4Arbiter_io_ifu_aw_ready & _T; // @[Crossbar.scala 155:47]
  assign AXILite2AXI4_1_io_mem_w_ready = AXI4Arbiter_io_ifu_w_ready; // @[Crossbar.scala 156:23]
  assign AXILite2AXI4_1_io_mem_b_valid = AXI4Arbiter_io_ifu_b_valid; // @[Crossbar.scala 157:23]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 38:23]
      istate <= 2'h0; // @[Crossbar.scala 38:23]
    end else if (2'h2 == istate) begin // @[Mux.scala 81:58]
      if (_istate_T_6) begin // @[Crossbar.scala 44:21]
        istate <= 2'h0;
      end else begin
        istate <= 2'h2;
      end
    end else if (2'h1 == istate) begin // @[Mux.scala 81:58]
      if (_istate_T_4) begin // @[Crossbar.scala 43:21]
        istate <= 2'h0;
      end else begin
        istate <= 2'h1;
      end
    end else if (2'h0 == istate) begin // @[Mux.scala 81:58]
      istate <= _istate_T_3;
    end else begin
      istate <= 2'h0;
    end
    if (reset) begin // @[Crossbar.scala 47:23]
      dstate <= 2'h0; // @[Crossbar.scala 47:23]
    end else if (2'h2 == dstate) begin // @[Mux.scala 81:58]
      if (_dstate_T_11 | _dstate_T_12) begin // @[Crossbar.scala 53:21]
        dstate <= 2'h0;
      end else begin
        dstate <= 2'h2;
      end
    end else if (2'h1 == dstate) begin // @[Mux.scala 81:58]
      if (_dstate_T_7 | _dstate_T_8) begin // @[Crossbar.scala 52:21]
        dstate <= 2'h0;
      end else begin
        dstate <= 2'h1;
      end
    end else if (2'h0 == dstate) begin // @[Mux.scala 81:58]
      dstate <= _dstate_T_6;
    end else begin
      dstate <= 2'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  istate = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  dstate = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module top(
  input         clock,
  input         reset,
  output [63:0] io_pc,
  output        io_valid,
  output [63:0] io_hitrate_i,
  output [63:0] io_hitrate_d
);
  wire  sram_clock; // @[top.scala 12:20]
  wire  sram_reset; // @[top.scala 12:20]
  wire  sram_io_ar_ready; // @[top.scala 12:20]
  wire  sram_io_ar_valid; // @[top.scala 12:20]
  wire [31:0] sram_io_ar_bits_addr; // @[top.scala 12:20]
  wire [7:0] sram_io_ar_bits_len; // @[top.scala 12:20]
  wire [2:0] sram_io_ar_bits_size; // @[top.scala 12:20]
  wire  sram_io_r_ready; // @[top.scala 12:20]
  wire  sram_io_r_valid; // @[top.scala 12:20]
  wire [63:0] sram_io_r_bits_data; // @[top.scala 12:20]
  wire  sram_io_aw_ready; // @[top.scala 12:20]
  wire  sram_io_aw_valid; // @[top.scala 12:20]
  wire [31:0] sram_io_aw_bits_addr; // @[top.scala 12:20]
  wire [2:0] sram_io_aw_bits_size; // @[top.scala 12:20]
  wire  sram_io_w_ready; // @[top.scala 12:20]
  wire  sram_io_w_valid; // @[top.scala 12:20]
  wire [63:0] sram_io_w_bits_data; // @[top.scala 12:20]
  wire [7:0] sram_io_w_bits_strb; // @[top.scala 12:20]
  wire  sram_io_w_bits_last; // @[top.scala 12:20]
  wire  sram_io_b_valid; // @[top.scala 12:20]
  wire  ifu_clock; // @[top.scala 13:19]
  wire  ifu_reset; // @[top.scala 13:19]
  wire [63:0] ifu_io_pc_dnpc; // @[top.scala 13:19]
  wire  ifu_io_clearJump; // @[top.scala 13:19]
  wire  ifu_io_lm_ar_ready; // @[top.scala 13:19]
  wire  ifu_io_lm_ar_valid; // @[top.scala 13:19]
  wire [31:0] ifu_io_lm_ar_bits_addr; // @[top.scala 13:19]
  wire  ifu_io_lm_r_ready; // @[top.scala 13:19]
  wire  ifu_io_lm_r_valid; // @[top.scala 13:19]
  wire [63:0] ifu_io_lm_r_bits_data; // @[top.scala 13:19]
  wire  ifu_io_out_ready; // @[top.scala 13:19]
  wire  ifu_io_out_valid; // @[top.scala 13:19]
  wire [31:0] ifu_io_out_bits_pc; // @[top.scala 13:19]
  wire [31:0] ifu_io_out_bits_inst; // @[top.scala 13:19]
  wire  ifu_io_out_bits_isJump; // @[top.scala 13:19]
  wire  idu_clock; // @[top.scala 14:19]
  wire  idu_reset; // @[top.scala 14:19]
  wire  idu_io_in_ready; // @[top.scala 14:19]
  wire  idu_io_in_valid; // @[top.scala 14:19]
  wire [31:0] idu_io_in_bits_pc; // @[top.scala 14:19]
  wire [31:0] idu_io_in_bits_inst; // @[top.scala 14:19]
  wire  idu_io_in_bits_isJump; // @[top.scala 14:19]
  wire  idu_io_out_ready; // @[top.scala 14:19]
  wire  idu_io_out_valid; // @[top.scala 14:19]
  wire [31:0] idu_io_out_bits_pc; // @[top.scala 14:19]
  wire [31:0] idu_io_out_bits_inst; // @[top.scala 14:19]
  wire [4:0] idu_io_out_bits_rs1; // @[top.scala 14:19]
  wire [4:0] idu_io_out_bits_rs2; // @[top.scala 14:19]
  wire [4:0] idu_io_out_bits_rd; // @[top.scala 14:19]
  wire [63:0] idu_io_out_bits_imm; // @[top.scala 14:19]
  wire [79:0] idu_io_out_bits_op; // @[top.scala 14:19]
  wire [5:0] idu_io_out_bits_typ; // @[top.scala 14:19]
  wire  idu_io_out_bits_isJump; // @[top.scala 14:19]
  wire [4:0] idu_io_out_bits_clearidx; // @[top.scala 14:19]
  wire [4:0] idu_io_sb_lookidx1; // @[top.scala 14:19]
  wire [4:0] idu_io_sb_lookidx2; // @[top.scala 14:19]
  wire [4:0] idu_io_sb_setidx; // @[top.scala 14:19]
  wire  idu_io_sb_isBusy; // @[top.scala 14:19]
  wire  exu_clock; // @[top.scala 15:19]
  wire  exu_reset; // @[top.scala 15:19]
  wire  exu_io_in_ready; // @[top.scala 15:19]
  wire  exu_io_in_valid; // @[top.scala 15:19]
  wire [31:0] exu_io_in_bits_pc; // @[top.scala 15:19]
  wire [31:0] exu_io_in_bits_inst; // @[top.scala 15:19]
  wire [4:0] exu_io_in_bits_rs1; // @[top.scala 15:19]
  wire [4:0] exu_io_in_bits_rs2; // @[top.scala 15:19]
  wire [4:0] exu_io_in_bits_rd; // @[top.scala 15:19]
  wire [63:0] exu_io_in_bits_imm; // @[top.scala 15:19]
  wire [79:0] exu_io_in_bits_op; // @[top.scala 15:19]
  wire [5:0] exu_io_in_bits_typ; // @[top.scala 15:19]
  wire  exu_io_in_bits_isJump; // @[top.scala 15:19]
  wire [4:0] exu_io_in_bits_clearidx; // @[top.scala 15:19]
  wire  exu_io_out_ready; // @[top.scala 15:19]
  wire  exu_io_out_valid; // @[top.scala 15:19]
  wire [31:0] exu_io_out_bits_pc; // @[top.scala 15:19]
  wire [63:0] exu_io_out_bits_pc_dnpc; // @[top.scala 15:19]
  wire [4:0] exu_io_out_bits_gpr_idx_w; // @[top.scala 15:19]
  wire  exu_io_out_bits_gpr_en_w; // @[top.scala 15:19]
  wire [63:0] exu_io_out_bits_gpr_val_w; // @[top.scala 15:19]
  wire  exu_io_out_bits_csr_en_w; // @[top.scala 15:19]
  wire [11:0] exu_io_out_bits_csr_idx_w; // @[top.scala 15:19]
  wire [63:0] exu_io_out_bits_csr_val_w; // @[top.scala 15:19]
  wire [63:0] exu_io_out_bits_csr_no; // @[top.scala 15:19]
  wire [63:0] exu_io_out_bits_csr_epc; // @[top.scala 15:19]
  wire  exu_io_out_bits_isJump; // @[top.scala 15:19]
  wire [4:0] exu_io_out_bits_clearidx; // @[top.scala 15:19]
  wire [4:0] exu_io_gpr_idx_r1; // @[top.scala 15:19]
  wire [4:0] exu_io_gpr_idx_r2; // @[top.scala 15:19]
  wire  exu_io_gpr_en_r1; // @[top.scala 15:19]
  wire  exu_io_gpr_en_r2; // @[top.scala 15:19]
  wire [63:0] exu_io_gpr_val_r1; // @[top.scala 15:19]
  wire [63:0] exu_io_gpr_val_r2; // @[top.scala 15:19]
  wire [11:0] exu_io_csr_idx_r; // @[top.scala 15:19]
  wire  exu_io_csr_en_r; // @[top.scala 15:19]
  wire [63:0] exu_io_csr_val_r; // @[top.scala 15:19]
  wire  exu_io_lm_ar_ready; // @[top.scala 15:19]
  wire  exu_io_lm_ar_valid; // @[top.scala 15:19]
  wire [31:0] exu_io_lm_ar_bits_addr; // @[top.scala 15:19]
  wire  exu_io_lm_r_ready; // @[top.scala 15:19]
  wire  exu_io_lm_r_valid; // @[top.scala 15:19]
  wire [63:0] exu_io_lm_r_bits_data; // @[top.scala 15:19]
  wire  exu_io_lm_aw_ready; // @[top.scala 15:19]
  wire  exu_io_lm_aw_valid; // @[top.scala 15:19]
  wire [31:0] exu_io_lm_aw_bits_addr; // @[top.scala 15:19]
  wire  exu_io_lm_w_ready; // @[top.scala 15:19]
  wire  exu_io_lm_w_valid; // @[top.scala 15:19]
  wire [63:0] exu_io_lm_w_bits_data; // @[top.scala 15:19]
  wire [7:0] exu_io_lm_w_bits_strb; // @[top.scala 15:19]
  wire  exu_io_lm_b_valid; // @[top.scala 15:19]
  wire  wbu_clock; // @[top.scala 16:19]
  wire  wbu_reset; // @[top.scala 16:19]
  wire  wbu_io_in_ready; // @[top.scala 16:19]
  wire  wbu_io_in_valid; // @[top.scala 16:19]
  wire [31:0] wbu_io_in_bits_pc; // @[top.scala 16:19]
  wire [63:0] wbu_io_in_bits_pc_dnpc; // @[top.scala 16:19]
  wire [4:0] wbu_io_in_bits_gpr_idx_w; // @[top.scala 16:19]
  wire  wbu_io_in_bits_gpr_en_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_in_bits_gpr_val_w; // @[top.scala 16:19]
  wire  wbu_io_in_bits_csr_en_w; // @[top.scala 16:19]
  wire [11:0] wbu_io_in_bits_csr_idx_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_in_bits_csr_val_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_in_bits_csr_no; // @[top.scala 16:19]
  wire [63:0] wbu_io_in_bits_csr_epc; // @[top.scala 16:19]
  wire  wbu_io_in_bits_isJump; // @[top.scala 16:19]
  wire [4:0] wbu_io_in_bits_clearidx; // @[top.scala 16:19]
  wire [4:0] wbu_io_gpr_idx_w; // @[top.scala 16:19]
  wire  wbu_io_gpr_en_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_gpr_val_w; // @[top.scala 16:19]
  wire  wbu_io_csr_en_w; // @[top.scala 16:19]
  wire [11:0] wbu_io_csr_idx_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_csr_val_w; // @[top.scala 16:19]
  wire [63:0] wbu_io_csr_no; // @[top.scala 16:19]
  wire [63:0] wbu_io_csr_epc; // @[top.scala 16:19]
  wire [63:0] wbu_io_pc_dnpc; // @[top.scala 16:19]
  wire  wbu_io_valid; // @[top.scala 16:19]
  wire  wbu_io_isJump; // @[top.scala 16:19]
  wire [4:0] wbu_io_sb_clearidx; // @[top.scala 16:19]
  wire  gpr_clock; // @[top.scala 17:19]
  wire  gpr_reset; // @[top.scala 17:19]
  wire [4:0] gpr_io_r_idx_r1; // @[top.scala 17:19]
  wire [4:0] gpr_io_r_idx_r2; // @[top.scala 17:19]
  wire  gpr_io_r_en_r1; // @[top.scala 17:19]
  wire  gpr_io_r_en_r2; // @[top.scala 17:19]
  wire [63:0] gpr_io_r_val_r1; // @[top.scala 17:19]
  wire [63:0] gpr_io_r_val_r2; // @[top.scala 17:19]
  wire [4:0] gpr_io_w_idx_w; // @[top.scala 17:19]
  wire  gpr_io_w_en_w; // @[top.scala 17:19]
  wire [63:0] gpr_io_w_val_w; // @[top.scala 17:19]
  wire  csr_clock; // @[top.scala 18:19]
  wire  csr_reset; // @[top.scala 18:19]
  wire [11:0] csr_io_r_idx_r; // @[top.scala 18:19]
  wire  csr_io_r_en_r; // @[top.scala 18:19]
  wire [63:0] csr_io_r_val_r; // @[top.scala 18:19]
  wire  csr_io_w_en_w; // @[top.scala 18:19]
  wire [11:0] csr_io_w_idx_w; // @[top.scala 18:19]
  wire [63:0] csr_io_w_val_w; // @[top.scala 18:19]
  wire [63:0] csr_io_w_no; // @[top.scala 18:19]
  wire [63:0] csr_io_w_epc; // @[top.scala 18:19]
  wire  scoreboard_clock; // @[top.scala 19:26]
  wire  scoreboard_reset; // @[top.scala 19:26]
  wire [4:0] scoreboard_io_ID_lookidx1; // @[top.scala 19:26]
  wire [4:0] scoreboard_io_ID_lookidx2; // @[top.scala 19:26]
  wire [4:0] scoreboard_io_ID_setidx; // @[top.scala 19:26]
  wire  scoreboard_io_ID_isBusy; // @[top.scala 19:26]
  wire [4:0] scoreboard_io_WB_clearidx; // @[top.scala 19:26]
  wire  crossbar_clock; // @[top.scala 36:24]
  wire  crossbar_reset; // @[top.scala 36:24]
  wire  crossbar_io_in1_ar_ready; // @[top.scala 36:24]
  wire  crossbar_io_in1_ar_valid; // @[top.scala 36:24]
  wire [31:0] crossbar_io_in1_ar_bits_addr; // @[top.scala 36:24]
  wire  crossbar_io_in1_r_valid; // @[top.scala 36:24]
  wire [63:0] crossbar_io_in1_r_bits_data; // @[top.scala 36:24]
  wire  crossbar_io_in2_ar_ready; // @[top.scala 36:24]
  wire  crossbar_io_in2_ar_valid; // @[top.scala 36:24]
  wire [31:0] crossbar_io_in2_ar_bits_addr; // @[top.scala 36:24]
  wire  crossbar_io_in2_r_ready; // @[top.scala 36:24]
  wire  crossbar_io_in2_r_valid; // @[top.scala 36:24]
  wire [63:0] crossbar_io_in2_r_bits_data; // @[top.scala 36:24]
  wire  crossbar_io_in2_aw_ready; // @[top.scala 36:24]
  wire  crossbar_io_in2_aw_valid; // @[top.scala 36:24]
  wire [31:0] crossbar_io_in2_aw_bits_addr; // @[top.scala 36:24]
  wire  crossbar_io_in2_w_ready; // @[top.scala 36:24]
  wire  crossbar_io_in2_w_valid; // @[top.scala 36:24]
  wire [63:0] crossbar_io_in2_w_bits_data; // @[top.scala 36:24]
  wire [7:0] crossbar_io_in2_w_bits_strb; // @[top.scala 36:24]
  wire  crossbar_io_in2_b_valid; // @[top.scala 36:24]
  wire  crossbar_io_out_ar_ready; // @[top.scala 36:24]
  wire  crossbar_io_out_ar_valid; // @[top.scala 36:24]
  wire [31:0] crossbar_io_out_ar_bits_addr; // @[top.scala 36:24]
  wire [7:0] crossbar_io_out_ar_bits_len; // @[top.scala 36:24]
  wire [2:0] crossbar_io_out_ar_bits_size; // @[top.scala 36:24]
  wire  crossbar_io_out_r_ready; // @[top.scala 36:24]
  wire  crossbar_io_out_r_valid; // @[top.scala 36:24]
  wire [63:0] crossbar_io_out_r_bits_data; // @[top.scala 36:24]
  wire  crossbar_io_out_aw_ready; // @[top.scala 36:24]
  wire  crossbar_io_out_aw_valid; // @[top.scala 36:24]
  wire [31:0] crossbar_io_out_aw_bits_addr; // @[top.scala 36:24]
  wire [2:0] crossbar_io_out_aw_bits_size; // @[top.scala 36:24]
  wire  crossbar_io_out_w_ready; // @[top.scala 36:24]
  wire  crossbar_io_out_w_valid; // @[top.scala 36:24]
  wire [63:0] crossbar_io_out_w_bits_data; // @[top.scala 36:24]
  wire [7:0] crossbar_io_out_w_bits_strb; // @[top.scala 36:24]
  wire  crossbar_io_out_w_bits_last; // @[top.scala 36:24]
  wire  crossbar_io_out_b_valid; // @[top.scala 36:24]
  wire [127:0] crossbar_io_hitrate; // @[top.scala 36:24]
  AXI4SRAM sram ( // @[top.scala 12:20]
    .clock(sram_clock),
    .reset(sram_reset),
    .io_ar_ready(sram_io_ar_ready),
    .io_ar_valid(sram_io_ar_valid),
    .io_ar_bits_addr(sram_io_ar_bits_addr),
    .io_ar_bits_len(sram_io_ar_bits_len),
    .io_ar_bits_size(sram_io_ar_bits_size),
    .io_r_ready(sram_io_r_ready),
    .io_r_valid(sram_io_r_valid),
    .io_r_bits_data(sram_io_r_bits_data),
    .io_aw_ready(sram_io_aw_ready),
    .io_aw_valid(sram_io_aw_valid),
    .io_aw_bits_addr(sram_io_aw_bits_addr),
    .io_aw_bits_size(sram_io_aw_bits_size),
    .io_w_ready(sram_io_w_ready),
    .io_w_valid(sram_io_w_valid),
    .io_w_bits_data(sram_io_w_bits_data),
    .io_w_bits_strb(sram_io_w_bits_strb),
    .io_w_bits_last(sram_io_w_bits_last),
    .io_b_valid(sram_io_b_valid)
  );
  IFU ifu ( // @[top.scala 13:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_pc_dnpc(ifu_io_pc_dnpc),
    .io_clearJump(ifu_io_clearJump),
    .io_lm_ar_ready(ifu_io_lm_ar_ready),
    .io_lm_ar_valid(ifu_io_lm_ar_valid),
    .io_lm_ar_bits_addr(ifu_io_lm_ar_bits_addr),
    .io_lm_r_ready(ifu_io_lm_r_ready),
    .io_lm_r_valid(ifu_io_lm_r_valid),
    .io_lm_r_bits_data(ifu_io_lm_r_bits_data),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_inst(ifu_io_out_bits_inst),
    .io_out_bits_isJump(ifu_io_out_bits_isJump)
  );
  IDU idu ( // @[top.scala 14:19]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_ready(idu_io_in_ready),
    .io_in_valid(idu_io_in_valid),
    .io_in_bits_pc(idu_io_in_bits_pc),
    .io_in_bits_inst(idu_io_in_bits_inst),
    .io_in_bits_isJump(idu_io_in_bits_isJump),
    .io_out_ready(idu_io_out_ready),
    .io_out_valid(idu_io_out_valid),
    .io_out_bits_pc(idu_io_out_bits_pc),
    .io_out_bits_inst(idu_io_out_bits_inst),
    .io_out_bits_rs1(idu_io_out_bits_rs1),
    .io_out_bits_rs2(idu_io_out_bits_rs2),
    .io_out_bits_rd(idu_io_out_bits_rd),
    .io_out_bits_imm(idu_io_out_bits_imm),
    .io_out_bits_op(idu_io_out_bits_op),
    .io_out_bits_typ(idu_io_out_bits_typ),
    .io_out_bits_isJump(idu_io_out_bits_isJump),
    .io_out_bits_clearidx(idu_io_out_bits_clearidx),
    .io_sb_lookidx1(idu_io_sb_lookidx1),
    .io_sb_lookidx2(idu_io_sb_lookidx2),
    .io_sb_setidx(idu_io_sb_setidx),
    .io_sb_isBusy(idu_io_sb_isBusy)
  );
  EXU exu ( // @[top.scala 15:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_in_ready(exu_io_in_ready),
    .io_in_valid(exu_io_in_valid),
    .io_in_bits_pc(exu_io_in_bits_pc),
    .io_in_bits_inst(exu_io_in_bits_inst),
    .io_in_bits_rs1(exu_io_in_bits_rs1),
    .io_in_bits_rs2(exu_io_in_bits_rs2),
    .io_in_bits_rd(exu_io_in_bits_rd),
    .io_in_bits_imm(exu_io_in_bits_imm),
    .io_in_bits_op(exu_io_in_bits_op),
    .io_in_bits_typ(exu_io_in_bits_typ),
    .io_in_bits_isJump(exu_io_in_bits_isJump),
    .io_in_bits_clearidx(exu_io_in_bits_clearidx),
    .io_out_ready(exu_io_out_ready),
    .io_out_valid(exu_io_out_valid),
    .io_out_bits_pc(exu_io_out_bits_pc),
    .io_out_bits_pc_dnpc(exu_io_out_bits_pc_dnpc),
    .io_out_bits_gpr_idx_w(exu_io_out_bits_gpr_idx_w),
    .io_out_bits_gpr_en_w(exu_io_out_bits_gpr_en_w),
    .io_out_bits_gpr_val_w(exu_io_out_bits_gpr_val_w),
    .io_out_bits_csr_en_w(exu_io_out_bits_csr_en_w),
    .io_out_bits_csr_idx_w(exu_io_out_bits_csr_idx_w),
    .io_out_bits_csr_val_w(exu_io_out_bits_csr_val_w),
    .io_out_bits_csr_no(exu_io_out_bits_csr_no),
    .io_out_bits_csr_epc(exu_io_out_bits_csr_epc),
    .io_out_bits_isJump(exu_io_out_bits_isJump),
    .io_out_bits_clearidx(exu_io_out_bits_clearidx),
    .io_gpr_idx_r1(exu_io_gpr_idx_r1),
    .io_gpr_idx_r2(exu_io_gpr_idx_r2),
    .io_gpr_en_r1(exu_io_gpr_en_r1),
    .io_gpr_en_r2(exu_io_gpr_en_r2),
    .io_gpr_val_r1(exu_io_gpr_val_r1),
    .io_gpr_val_r2(exu_io_gpr_val_r2),
    .io_csr_idx_r(exu_io_csr_idx_r),
    .io_csr_en_r(exu_io_csr_en_r),
    .io_csr_val_r(exu_io_csr_val_r),
    .io_lm_ar_ready(exu_io_lm_ar_ready),
    .io_lm_ar_valid(exu_io_lm_ar_valid),
    .io_lm_ar_bits_addr(exu_io_lm_ar_bits_addr),
    .io_lm_r_ready(exu_io_lm_r_ready),
    .io_lm_r_valid(exu_io_lm_r_valid),
    .io_lm_r_bits_data(exu_io_lm_r_bits_data),
    .io_lm_aw_ready(exu_io_lm_aw_ready),
    .io_lm_aw_valid(exu_io_lm_aw_valid),
    .io_lm_aw_bits_addr(exu_io_lm_aw_bits_addr),
    .io_lm_w_ready(exu_io_lm_w_ready),
    .io_lm_w_valid(exu_io_lm_w_valid),
    .io_lm_w_bits_data(exu_io_lm_w_bits_data),
    .io_lm_w_bits_strb(exu_io_lm_w_bits_strb),
    .io_lm_b_valid(exu_io_lm_b_valid)
  );
  WBU wbu ( // @[top.scala 16:19]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io_in_ready(wbu_io_in_ready),
    .io_in_valid(wbu_io_in_valid),
    .io_in_bits_pc(wbu_io_in_bits_pc),
    .io_in_bits_pc_dnpc(wbu_io_in_bits_pc_dnpc),
    .io_in_bits_gpr_idx_w(wbu_io_in_bits_gpr_idx_w),
    .io_in_bits_gpr_en_w(wbu_io_in_bits_gpr_en_w),
    .io_in_bits_gpr_val_w(wbu_io_in_bits_gpr_val_w),
    .io_in_bits_csr_en_w(wbu_io_in_bits_csr_en_w),
    .io_in_bits_csr_idx_w(wbu_io_in_bits_csr_idx_w),
    .io_in_bits_csr_val_w(wbu_io_in_bits_csr_val_w),
    .io_in_bits_csr_no(wbu_io_in_bits_csr_no),
    .io_in_bits_csr_epc(wbu_io_in_bits_csr_epc),
    .io_in_bits_isJump(wbu_io_in_bits_isJump),
    .io_in_bits_clearidx(wbu_io_in_bits_clearidx),
    .io_gpr_idx_w(wbu_io_gpr_idx_w),
    .io_gpr_en_w(wbu_io_gpr_en_w),
    .io_gpr_val_w(wbu_io_gpr_val_w),
    .io_csr_en_w(wbu_io_csr_en_w),
    .io_csr_idx_w(wbu_io_csr_idx_w),
    .io_csr_val_w(wbu_io_csr_val_w),
    .io_csr_no(wbu_io_csr_no),
    .io_csr_epc(wbu_io_csr_epc),
    .io_pc_dnpc(wbu_io_pc_dnpc),
    .io_valid(wbu_io_valid),
    .io_isJump(wbu_io_isJump),
    .io_sb_clearidx(wbu_io_sb_clearidx)
  );
  GPR gpr ( // @[top.scala 17:19]
    .clock(gpr_clock),
    .reset(gpr_reset),
    .io_r_idx_r1(gpr_io_r_idx_r1),
    .io_r_idx_r2(gpr_io_r_idx_r2),
    .io_r_en_r1(gpr_io_r_en_r1),
    .io_r_en_r2(gpr_io_r_en_r2),
    .io_r_val_r1(gpr_io_r_val_r1),
    .io_r_val_r2(gpr_io_r_val_r2),
    .io_w_idx_w(gpr_io_w_idx_w),
    .io_w_en_w(gpr_io_w_en_w),
    .io_w_val_w(gpr_io_w_val_w)
  );
  CSR csr ( // @[top.scala 18:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_r_idx_r(csr_io_r_idx_r),
    .io_r_en_r(csr_io_r_en_r),
    .io_r_val_r(csr_io_r_val_r),
    .io_w_en_w(csr_io_w_en_w),
    .io_w_idx_w(csr_io_w_idx_w),
    .io_w_val_w(csr_io_w_val_w),
    .io_w_no(csr_io_w_no),
    .io_w_epc(csr_io_w_epc)
  );
  ScoreBoard scoreboard ( // @[top.scala 19:26]
    .clock(scoreboard_clock),
    .reset(scoreboard_reset),
    .io_ID_lookidx1(scoreboard_io_ID_lookidx1),
    .io_ID_lookidx2(scoreboard_io_ID_lookidx2),
    .io_ID_setidx(scoreboard_io_ID_setidx),
    .io_ID_isBusy(scoreboard_io_ID_isBusy),
    .io_WB_clearidx(scoreboard_io_WB_clearidx)
  );
  Crossbar crossbar ( // @[top.scala 36:24]
    .clock(crossbar_clock),
    .reset(crossbar_reset),
    .io_in1_ar_ready(crossbar_io_in1_ar_ready),
    .io_in1_ar_valid(crossbar_io_in1_ar_valid),
    .io_in1_ar_bits_addr(crossbar_io_in1_ar_bits_addr),
    .io_in1_r_valid(crossbar_io_in1_r_valid),
    .io_in1_r_bits_data(crossbar_io_in1_r_bits_data),
    .io_in2_ar_ready(crossbar_io_in2_ar_ready),
    .io_in2_ar_valid(crossbar_io_in2_ar_valid),
    .io_in2_ar_bits_addr(crossbar_io_in2_ar_bits_addr),
    .io_in2_r_ready(crossbar_io_in2_r_ready),
    .io_in2_r_valid(crossbar_io_in2_r_valid),
    .io_in2_r_bits_data(crossbar_io_in2_r_bits_data),
    .io_in2_aw_ready(crossbar_io_in2_aw_ready),
    .io_in2_aw_valid(crossbar_io_in2_aw_valid),
    .io_in2_aw_bits_addr(crossbar_io_in2_aw_bits_addr),
    .io_in2_w_ready(crossbar_io_in2_w_ready),
    .io_in2_w_valid(crossbar_io_in2_w_valid),
    .io_in2_w_bits_data(crossbar_io_in2_w_bits_data),
    .io_in2_w_bits_strb(crossbar_io_in2_w_bits_strb),
    .io_in2_b_valid(crossbar_io_in2_b_valid),
    .io_out_ar_ready(crossbar_io_out_ar_ready),
    .io_out_ar_valid(crossbar_io_out_ar_valid),
    .io_out_ar_bits_addr(crossbar_io_out_ar_bits_addr),
    .io_out_ar_bits_len(crossbar_io_out_ar_bits_len),
    .io_out_ar_bits_size(crossbar_io_out_ar_bits_size),
    .io_out_r_ready(crossbar_io_out_r_ready),
    .io_out_r_valid(crossbar_io_out_r_valid),
    .io_out_r_bits_data(crossbar_io_out_r_bits_data),
    .io_out_aw_ready(crossbar_io_out_aw_ready),
    .io_out_aw_valid(crossbar_io_out_aw_valid),
    .io_out_aw_bits_addr(crossbar_io_out_aw_bits_addr),
    .io_out_aw_bits_size(crossbar_io_out_aw_bits_size),
    .io_out_w_ready(crossbar_io_out_w_ready),
    .io_out_w_valid(crossbar_io_out_w_valid),
    .io_out_w_bits_data(crossbar_io_out_w_bits_data),
    .io_out_w_bits_strb(crossbar_io_out_w_bits_strb),
    .io_out_w_bits_last(crossbar_io_out_w_bits_last),
    .io_out_b_valid(crossbar_io_out_b_valid),
    .io_hitrate(crossbar_io_hitrate)
  );
  assign io_pc = wbu_io_pc_dnpc; // @[top.scala 34:10]
  assign io_valid = wbu_io_valid; // @[top.scala 33:13]
  assign io_hitrate_i = crossbar_io_hitrate[127:64]; // @[top.scala 42:38]
  assign io_hitrate_d = crossbar_io_hitrate[63:0]; // @[top.scala 43:38]
  assign sram_clock = clock;
  assign sram_reset = reset;
  assign sram_io_ar_valid = crossbar_io_out_ar_valid; // @[top.scala 39:20]
  assign sram_io_ar_bits_addr = crossbar_io_out_ar_bits_addr; // @[top.scala 39:20]
  assign sram_io_ar_bits_len = crossbar_io_out_ar_bits_len; // @[top.scala 39:20]
  assign sram_io_ar_bits_size = crossbar_io_out_ar_bits_size; // @[top.scala 39:20]
  assign sram_io_r_ready = crossbar_io_out_r_ready; // @[top.scala 39:20]
  assign sram_io_aw_valid = crossbar_io_out_aw_valid; // @[top.scala 39:20]
  assign sram_io_aw_bits_addr = crossbar_io_out_aw_bits_addr; // @[top.scala 39:20]
  assign sram_io_aw_bits_size = crossbar_io_out_aw_bits_size; // @[top.scala 39:20]
  assign sram_io_w_valid = crossbar_io_out_w_valid; // @[top.scala 39:20]
  assign sram_io_w_bits_data = crossbar_io_out_w_bits_data; // @[top.scala 39:20]
  assign sram_io_w_bits_strb = crossbar_io_out_w_bits_strb; // @[top.scala 39:20]
  assign sram_io_w_bits_last = crossbar_io_out_w_bits_last; // @[top.scala 39:20]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_pc_dnpc = wbu_io_pc_dnpc; // @[top.scala 23:19]
  assign ifu_io_clearJump = wbu_io_isJump; // @[top.scala 24:21]
  assign ifu_io_lm_ar_ready = crossbar_io_in1_ar_ready; // @[top.scala 37:20]
  assign ifu_io_lm_r_valid = crossbar_io_in1_r_valid; // @[top.scala 37:20]
  assign ifu_io_lm_r_bits_data = crossbar_io_in1_r_bits_data; // @[top.scala 37:20]
  assign ifu_io_out_ready = idu_io_in_ready; // @[top.scala 25:14]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_valid = ifu_io_out_valid; // @[top.scala 25:14]
  assign idu_io_in_bits_pc = ifu_io_out_bits_pc; // @[top.scala 25:14]
  assign idu_io_in_bits_inst = ifu_io_out_bits_inst; // @[top.scala 25:14]
  assign idu_io_in_bits_isJump = ifu_io_out_bits_isJump; // @[top.scala 25:14]
  assign idu_io_out_ready = exu_io_in_ready; // @[top.scala 26:14]
  assign idu_io_sb_isBusy = scoreboard_io_ID_isBusy; // @[top.scala 21:21]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_in_valid = idu_io_out_valid; // @[top.scala 26:14]
  assign exu_io_in_bits_pc = idu_io_out_bits_pc; // @[top.scala 26:14]
  assign exu_io_in_bits_inst = idu_io_out_bits_inst; // @[top.scala 26:14]
  assign exu_io_in_bits_rs1 = idu_io_out_bits_rs1; // @[top.scala 26:14]
  assign exu_io_in_bits_rs2 = idu_io_out_bits_rs2; // @[top.scala 26:14]
  assign exu_io_in_bits_rd = idu_io_out_bits_rd; // @[top.scala 26:14]
  assign exu_io_in_bits_imm = idu_io_out_bits_imm; // @[top.scala 26:14]
  assign exu_io_in_bits_op = idu_io_out_bits_op; // @[top.scala 26:14]
  assign exu_io_in_bits_typ = idu_io_out_bits_typ; // @[top.scala 26:14]
  assign exu_io_in_bits_isJump = idu_io_out_bits_isJump; // @[top.scala 26:14]
  assign exu_io_in_bits_clearidx = idu_io_out_bits_clearidx; // @[top.scala 26:14]
  assign exu_io_out_ready = wbu_io_in_ready; // @[top.scala 29:14]
  assign exu_io_gpr_val_r1 = gpr_io_r_val_r1; // @[top.scala 27:15]
  assign exu_io_gpr_val_r2 = gpr_io_r_val_r2; // @[top.scala 27:15]
  assign exu_io_csr_val_r = csr_io_r_val_r; // @[top.scala 28:15]
  assign exu_io_lm_ar_ready = crossbar_io_in2_ar_ready; // @[top.scala 38:20]
  assign exu_io_lm_r_valid = crossbar_io_in2_r_valid; // @[top.scala 38:20]
  assign exu_io_lm_r_bits_data = crossbar_io_in2_r_bits_data; // @[top.scala 38:20]
  assign exu_io_lm_aw_ready = crossbar_io_in2_aw_ready; // @[top.scala 38:20]
  assign exu_io_lm_w_ready = crossbar_io_in2_w_ready; // @[top.scala 38:20]
  assign exu_io_lm_b_valid = crossbar_io_in2_b_valid; // @[top.scala 38:20]
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io_in_valid = exu_io_out_valid; // @[top.scala 29:14]
  assign wbu_io_in_bits_pc = exu_io_out_bits_pc; // @[top.scala 29:14]
  assign wbu_io_in_bits_pc_dnpc = exu_io_out_bits_pc_dnpc; // @[top.scala 29:14]
  assign wbu_io_in_bits_gpr_idx_w = exu_io_out_bits_gpr_idx_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_gpr_en_w = exu_io_out_bits_gpr_en_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_gpr_val_w = exu_io_out_bits_gpr_val_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_csr_en_w = exu_io_out_bits_csr_en_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_csr_idx_w = exu_io_out_bits_csr_idx_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_csr_val_w = exu_io_out_bits_csr_val_w; // @[top.scala 29:14]
  assign wbu_io_in_bits_csr_no = exu_io_out_bits_csr_no; // @[top.scala 29:14]
  assign wbu_io_in_bits_csr_epc = exu_io_out_bits_csr_epc; // @[top.scala 29:14]
  assign wbu_io_in_bits_isJump = exu_io_out_bits_isJump; // @[top.scala 29:14]
  assign wbu_io_in_bits_clearidx = exu_io_out_bits_clearidx; // @[top.scala 29:14]
  assign gpr_clock = clock;
  assign gpr_reset = reset;
  assign gpr_io_r_idx_r1 = exu_io_gpr_idx_r1; // @[top.scala 27:15]
  assign gpr_io_r_idx_r2 = exu_io_gpr_idx_r2; // @[top.scala 27:15]
  assign gpr_io_r_en_r1 = exu_io_gpr_en_r1; // @[top.scala 27:15]
  assign gpr_io_r_en_r2 = exu_io_gpr_en_r2; // @[top.scala 27:15]
  assign gpr_io_w_idx_w = wbu_io_gpr_idx_w; // @[top.scala 30:15]
  assign gpr_io_w_en_w = wbu_io_gpr_en_w; // @[top.scala 30:15]
  assign gpr_io_w_val_w = wbu_io_gpr_val_w; // @[top.scala 30:15]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_r_idx_r = exu_io_csr_idx_r; // @[top.scala 28:15]
  assign csr_io_r_en_r = exu_io_csr_en_r; // @[top.scala 28:15]
  assign csr_io_w_en_w = wbu_io_csr_en_w; // @[top.scala 31:15]
  assign csr_io_w_idx_w = wbu_io_csr_idx_w; // @[top.scala 31:15]
  assign csr_io_w_val_w = wbu_io_csr_val_w; // @[top.scala 31:15]
  assign csr_io_w_no = wbu_io_csr_no; // @[top.scala 31:15]
  assign csr_io_w_epc = wbu_io_csr_epc; // @[top.scala 31:15]
  assign scoreboard_clock = clock;
  assign scoreboard_reset = reset;
  assign scoreboard_io_ID_lookidx1 = idu_io_sb_lookidx1; // @[top.scala 21:21]
  assign scoreboard_io_ID_lookidx2 = idu_io_sb_lookidx2; // @[top.scala 21:21]
  assign scoreboard_io_ID_setidx = idu_io_sb_setidx; // @[top.scala 21:21]
  assign scoreboard_io_WB_clearidx = wbu_io_sb_clearidx; // @[top.scala 22:21]
  assign crossbar_clock = clock;
  assign crossbar_reset = reset;
  assign crossbar_io_in1_ar_valid = ifu_io_lm_ar_valid; // @[top.scala 37:20]
  assign crossbar_io_in1_ar_bits_addr = ifu_io_lm_ar_bits_addr; // @[top.scala 37:20]
  assign crossbar_io_in2_ar_valid = exu_io_lm_ar_valid; // @[top.scala 38:20]
  assign crossbar_io_in2_ar_bits_addr = exu_io_lm_ar_bits_addr; // @[top.scala 38:20]
  assign crossbar_io_in2_r_ready = exu_io_lm_r_ready; // @[top.scala 38:20]
  assign crossbar_io_in2_aw_valid = exu_io_lm_aw_valid; // @[top.scala 38:20]
  assign crossbar_io_in2_aw_bits_addr = exu_io_lm_aw_bits_addr; // @[top.scala 38:20]
  assign crossbar_io_in2_w_valid = exu_io_lm_w_valid; // @[top.scala 38:20]
  assign crossbar_io_in2_w_bits_data = exu_io_lm_w_bits_data; // @[top.scala 38:20]
  assign crossbar_io_in2_w_bits_strb = exu_io_lm_w_bits_strb; // @[top.scala 38:20]
  assign crossbar_io_out_ar_ready = sram_io_ar_ready; // @[top.scala 39:20]
  assign crossbar_io_out_r_valid = sram_io_r_valid; // @[top.scala 39:20]
  assign crossbar_io_out_r_bits_data = sram_io_r_bits_data; // @[top.scala 39:20]
  assign crossbar_io_out_aw_ready = sram_io_aw_ready; // @[top.scala 39:20]
  assign crossbar_io_out_w_ready = sram_io_w_ready; // @[top.scala 39:20]
  assign crossbar_io_out_b_valid = sram_io_b_valid; // @[top.scala 39:20]
endmodule
