module toptest;
initial
begin
	$dumpfile("top.vcd");
	$dumpvars(0,toptest);
end
endmodule
