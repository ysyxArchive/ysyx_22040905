module gen_sel(
  input  [2:0] io_src,
  output [3:0] io_out
);
  wire  y_sub = io_src[0]; // @[WallaceTest.scala 55:21]
  wire  y = io_src[1]; // @[WallaceTest.scala 56:16]
  wire  y_add = io_src[2]; // @[WallaceTest.scala 57:20]
  wire  _sel_negative_T = ~y_sub; // @[WallaceTest.scala 59:36]
  wire  _sel_negative_T_2 = ~y; // @[WallaceTest.scala 59:45]
  wire  _sel_negative_T_4 = y & ~y_sub | ~y & y_sub; // @[WallaceTest.scala 59:43]
  wire  sel_negative = y_add & (y & ~y_sub | ~y & y_sub); // @[WallaceTest.scala 59:29]
  wire  _sel_positive_T = ~y_add; // @[WallaceTest.scala 60:23]
  wire  sel_positive = ~y_add & _sel_negative_T_4; // @[WallaceTest.scala 60:30]
  wire  sel_double_negative = y_add & _sel_negative_T_2 & _sel_negative_T; // @[WallaceTest.scala 61:41]
  wire  sel_double_positive = _sel_positive_T & y & y_sub; // @[WallaceTest.scala 62:41]
  wire [1:0] io_out_lo = {sel_positive,sel_negative}; // @[Cat.scala 33:92]
  wire [1:0] io_out_hi = {sel_double_positive,sel_double_negative}; // @[Cat.scala 33:92]
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 33:92]
endmodule
module gen_p_i(
  input        io_x,
  input        io_x_sub,
  input  [3:0] io_sel,
  output       io_p
);
  wire  sel_negative = io_sel[0]; // @[WallaceTest.scala 40:26]
  wire  sel_positive = io_sel[1]; // @[WallaceTest.scala 41:26]
  wire  sel_double_negative = io_sel[2]; // @[WallaceTest.scala 42:33]
  wire  sel_double_positive = io_sel[3]; // @[WallaceTest.scala 43:33]
  wire  _io_p_T_6 = ~(sel_negative & ~io_x) & ~(sel_double_negative & ~io_x_sub); // @[WallaceTest.scala 45:37]
  wire  _io_p_T_12 = _io_p_T_6 & ~(sel_positive & io_x) & ~(sel_double_positive & io_x_sub); // @[WallaceTest.scala 46:37]
  assign io_p = ~_io_p_T_12; // @[WallaceTest.scala 45:11]
endmodule
module gen_p(
  input  [2:0]   io_src,
  input  [131:0] io_x,
  output [131:0] io_p,
  output         io_c
);
  wire [2:0] gen_sel_io_src; // @[WallaceTest.scala 75:17]
  wire [3:0] gen_sel_io_out; // @[WallaceTest.scala 75:17]
  wire  gen_p_i_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_1_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_1_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_1_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_1_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_2_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_2_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_2_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_2_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_3_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_3_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_3_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_3_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_4_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_4_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_4_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_4_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_5_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_5_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_5_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_5_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_6_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_6_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_6_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_6_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_7_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_7_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_7_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_7_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_8_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_8_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_8_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_8_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_9_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_9_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_9_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_9_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_10_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_10_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_10_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_10_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_11_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_11_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_11_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_11_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_12_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_12_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_12_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_12_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_13_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_13_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_13_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_13_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_14_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_14_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_14_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_14_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_15_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_15_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_15_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_15_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_16_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_16_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_16_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_16_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_17_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_17_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_17_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_17_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_18_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_18_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_18_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_18_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_19_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_19_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_19_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_19_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_20_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_20_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_20_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_20_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_21_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_21_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_21_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_21_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_22_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_22_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_22_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_22_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_23_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_23_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_23_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_23_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_24_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_24_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_24_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_24_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_25_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_25_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_25_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_25_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_26_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_26_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_26_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_26_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_27_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_27_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_27_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_27_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_28_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_28_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_28_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_28_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_29_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_29_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_29_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_29_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_30_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_30_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_30_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_30_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_31_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_31_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_31_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_31_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_32_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_32_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_32_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_32_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_33_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_33_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_33_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_33_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_34_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_34_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_34_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_34_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_35_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_35_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_35_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_35_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_36_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_36_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_36_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_36_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_37_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_37_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_37_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_37_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_38_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_38_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_38_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_38_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_39_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_39_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_39_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_39_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_40_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_40_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_40_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_40_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_41_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_41_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_41_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_41_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_42_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_42_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_42_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_42_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_43_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_43_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_43_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_43_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_44_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_44_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_44_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_44_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_45_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_45_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_45_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_45_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_46_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_46_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_46_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_46_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_47_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_47_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_47_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_47_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_48_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_48_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_48_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_48_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_49_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_49_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_49_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_49_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_50_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_50_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_50_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_50_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_51_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_51_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_51_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_51_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_52_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_52_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_52_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_52_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_53_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_53_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_53_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_53_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_54_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_54_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_54_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_54_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_55_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_55_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_55_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_55_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_56_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_56_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_56_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_56_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_57_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_57_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_57_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_57_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_58_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_58_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_58_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_58_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_59_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_59_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_59_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_59_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_60_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_60_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_60_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_60_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_61_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_61_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_61_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_61_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_62_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_62_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_62_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_62_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_63_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_63_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_63_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_63_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_64_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_64_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_64_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_64_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_65_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_65_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_65_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_65_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_66_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_66_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_66_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_66_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_67_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_67_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_67_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_67_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_68_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_68_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_68_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_68_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_69_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_69_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_69_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_69_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_70_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_70_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_70_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_70_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_71_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_71_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_71_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_71_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_72_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_72_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_72_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_72_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_73_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_73_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_73_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_73_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_74_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_74_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_74_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_74_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_75_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_75_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_75_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_75_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_76_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_76_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_76_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_76_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_77_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_77_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_77_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_77_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_78_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_78_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_78_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_78_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_79_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_79_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_79_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_79_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_80_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_80_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_80_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_80_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_81_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_81_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_81_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_81_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_82_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_82_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_82_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_82_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_83_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_83_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_83_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_83_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_84_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_84_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_84_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_84_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_85_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_85_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_85_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_85_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_86_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_86_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_86_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_86_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_87_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_87_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_87_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_87_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_88_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_88_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_88_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_88_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_89_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_89_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_89_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_89_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_90_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_90_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_90_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_90_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_91_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_91_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_91_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_91_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_92_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_92_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_92_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_92_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_93_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_93_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_93_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_93_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_94_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_94_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_94_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_94_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_95_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_95_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_95_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_95_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_96_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_96_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_96_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_96_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_97_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_97_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_97_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_97_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_98_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_98_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_98_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_98_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_99_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_99_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_99_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_99_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_100_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_100_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_100_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_100_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_101_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_101_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_101_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_101_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_102_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_102_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_102_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_102_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_103_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_103_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_103_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_103_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_104_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_104_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_104_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_104_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_105_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_105_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_105_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_105_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_106_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_106_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_106_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_106_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_107_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_107_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_107_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_107_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_108_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_108_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_108_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_108_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_109_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_109_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_109_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_109_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_110_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_110_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_110_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_110_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_111_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_111_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_111_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_111_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_112_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_112_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_112_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_112_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_113_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_113_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_113_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_113_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_114_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_114_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_114_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_114_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_115_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_115_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_115_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_115_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_116_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_116_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_116_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_116_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_117_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_117_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_117_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_117_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_118_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_118_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_118_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_118_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_119_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_119_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_119_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_119_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_120_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_120_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_120_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_120_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_121_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_121_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_121_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_121_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_122_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_122_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_122_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_122_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_123_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_123_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_123_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_123_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_124_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_124_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_124_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_124_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_125_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_125_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_125_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_125_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_126_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_126_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_126_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_126_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_127_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_127_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_127_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_127_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_128_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_128_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_128_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_128_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_129_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_129_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_129_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_129_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_130_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_130_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_130_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_130_io_p; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_131_io_x; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_131_io_x_sub; // @[WallaceTest.scala 76:29]
  wire [3:0] gen_p_i_131_io_sel; // @[WallaceTest.scala 76:29]
  wire  gen_p_i_131_io_p; // @[WallaceTest.scala 76:29]
  wire [7:0] io_p_lo_lo_lo_lo = {gen_p_i_7_io_p,gen_p_i_6_io_p,gen_p_i_5_io_p,gen_p_i_4_io_p,gen_p_i_3_io_p,
    gen_p_i_2_io_p,gen_p_i_1_io_p,gen_p_i_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_lo_hi_lo = {gen_p_i_23_io_p,gen_p_i_22_io_p,gen_p_i_21_io_p,gen_p_i_20_io_p,gen_p_i_19_io_p,
    gen_p_i_18_io_p,gen_p_i_17_io_p,gen_p_i_16_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_lo_lo_hi = {gen_p_i_32_io_p,gen_p_i_31_io_p,gen_p_i_30_io_p,gen_p_i_29_io_p,gen_p_i_28_io_p,
    gen_p_i_27_io_p,gen_p_i_26_io_p,gen_p_i_25_io_p,gen_p_i_24_io_p,io_p_lo_lo_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_lo_lo = {io_p_lo_lo_hi,gen_p_i_15_io_p,gen_p_i_14_io_p,gen_p_i_13_io_p,gen_p_i_12_io_p,
    gen_p_i_11_io_p,gen_p_i_10_io_p,gen_p_i_9_io_p,gen_p_i_8_io_p,io_p_lo_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_hi_lo_lo = {gen_p_i_40_io_p,gen_p_i_39_io_p,gen_p_i_38_io_p,gen_p_i_37_io_p,gen_p_i_36_io_p,
    gen_p_i_35_io_p,gen_p_i_34_io_p,gen_p_i_33_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_lo_hi_hi_lo = {gen_p_i_56_io_p,gen_p_i_55_io_p,gen_p_i_54_io_p,gen_p_i_53_io_p,gen_p_i_52_io_p,
    gen_p_i_51_io_p,gen_p_i_50_io_p,gen_p_i_49_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_lo_hi_hi = {gen_p_i_65_io_p,gen_p_i_64_io_p,gen_p_i_63_io_p,gen_p_i_62_io_p,gen_p_i_61_io_p,
    gen_p_i_60_io_p,gen_p_i_59_io_p,gen_p_i_58_io_p,gen_p_i_57_io_p,io_p_lo_hi_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_lo_hi = {io_p_lo_hi_hi,gen_p_i_48_io_p,gen_p_i_47_io_p,gen_p_i_46_io_p,gen_p_i_45_io_p,
    gen_p_i_44_io_p,gen_p_i_43_io_p,gen_p_i_42_io_p,gen_p_i_41_io_p,io_p_lo_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [65:0] io_p_lo = {io_p_lo_hi,io_p_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_lo_lo_lo = {gen_p_i_73_io_p,gen_p_i_72_io_p,gen_p_i_71_io_p,gen_p_i_70_io_p,gen_p_i_69_io_p,
    gen_p_i_68_io_p,gen_p_i_67_io_p,gen_p_i_66_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_lo_hi_lo = {gen_p_i_89_io_p,gen_p_i_88_io_p,gen_p_i_87_io_p,gen_p_i_86_io_p,gen_p_i_85_io_p,
    gen_p_i_84_io_p,gen_p_i_83_io_p,gen_p_i_82_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_hi_lo_hi = {gen_p_i_98_io_p,gen_p_i_97_io_p,gen_p_i_96_io_p,gen_p_i_95_io_p,gen_p_i_94_io_p,
    gen_p_i_93_io_p,gen_p_i_92_io_p,gen_p_i_91_io_p,gen_p_i_90_io_p,io_p_hi_lo_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_hi_lo = {io_p_hi_lo_hi,gen_p_i_81_io_p,gen_p_i_80_io_p,gen_p_i_79_io_p,gen_p_i_78_io_p,
    gen_p_i_77_io_p,gen_p_i_76_io_p,gen_p_i_75_io_p,gen_p_i_74_io_p,io_p_hi_lo_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_hi_lo_lo = {gen_p_i_106_io_p,gen_p_i_105_io_p,gen_p_i_104_io_p,gen_p_i_103_io_p,gen_p_i_102_io_p,
    gen_p_i_101_io_p,gen_p_i_100_io_p,gen_p_i_99_io_p}; // @[Cat.scala 33:92]
  wire [7:0] io_p_hi_hi_hi_lo = {gen_p_i_122_io_p,gen_p_i_121_io_p,gen_p_i_120_io_p,gen_p_i_119_io_p,gen_p_i_118_io_p,
    gen_p_i_117_io_p,gen_p_i_116_io_p,gen_p_i_115_io_p}; // @[Cat.scala 33:92]
  wire [16:0] io_p_hi_hi_hi = {gen_p_i_131_io_p,gen_p_i_130_io_p,gen_p_i_129_io_p,gen_p_i_128_io_p,gen_p_i_127_io_p,
    gen_p_i_126_io_p,gen_p_i_125_io_p,gen_p_i_124_io_p,gen_p_i_123_io_p,io_p_hi_hi_hi_lo}; // @[Cat.scala 33:92]
  wire [32:0] io_p_hi_hi = {io_p_hi_hi_hi,gen_p_i_114_io_p,gen_p_i_113_io_p,gen_p_i_112_io_p,gen_p_i_111_io_p,
    gen_p_i_110_io_p,gen_p_i_109_io_p,gen_p_i_108_io_p,gen_p_i_107_io_p,io_p_hi_hi_lo_lo}; // @[Cat.scala 33:92]
  wire [65:0] io_p_hi = {io_p_hi_hi,io_p_hi_lo}; // @[Cat.scala 33:92]
  gen_sel gen_sel ( // @[WallaceTest.scala 75:17]
    .io_src(gen_sel_io_src),
    .io_out(gen_sel_io_out)
  );
  gen_p_i gen_p_i ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_io_x),
    .io_x_sub(gen_p_i_io_x_sub),
    .io_sel(gen_p_i_io_sel),
    .io_p(gen_p_i_io_p)
  );
  gen_p_i gen_p_i_1 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_1_io_x),
    .io_x_sub(gen_p_i_1_io_x_sub),
    .io_sel(gen_p_i_1_io_sel),
    .io_p(gen_p_i_1_io_p)
  );
  gen_p_i gen_p_i_2 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_2_io_x),
    .io_x_sub(gen_p_i_2_io_x_sub),
    .io_sel(gen_p_i_2_io_sel),
    .io_p(gen_p_i_2_io_p)
  );
  gen_p_i gen_p_i_3 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_3_io_x),
    .io_x_sub(gen_p_i_3_io_x_sub),
    .io_sel(gen_p_i_3_io_sel),
    .io_p(gen_p_i_3_io_p)
  );
  gen_p_i gen_p_i_4 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_4_io_x),
    .io_x_sub(gen_p_i_4_io_x_sub),
    .io_sel(gen_p_i_4_io_sel),
    .io_p(gen_p_i_4_io_p)
  );
  gen_p_i gen_p_i_5 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_5_io_x),
    .io_x_sub(gen_p_i_5_io_x_sub),
    .io_sel(gen_p_i_5_io_sel),
    .io_p(gen_p_i_5_io_p)
  );
  gen_p_i gen_p_i_6 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_6_io_x),
    .io_x_sub(gen_p_i_6_io_x_sub),
    .io_sel(gen_p_i_6_io_sel),
    .io_p(gen_p_i_6_io_p)
  );
  gen_p_i gen_p_i_7 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_7_io_x),
    .io_x_sub(gen_p_i_7_io_x_sub),
    .io_sel(gen_p_i_7_io_sel),
    .io_p(gen_p_i_7_io_p)
  );
  gen_p_i gen_p_i_8 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_8_io_x),
    .io_x_sub(gen_p_i_8_io_x_sub),
    .io_sel(gen_p_i_8_io_sel),
    .io_p(gen_p_i_8_io_p)
  );
  gen_p_i gen_p_i_9 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_9_io_x),
    .io_x_sub(gen_p_i_9_io_x_sub),
    .io_sel(gen_p_i_9_io_sel),
    .io_p(gen_p_i_9_io_p)
  );
  gen_p_i gen_p_i_10 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_10_io_x),
    .io_x_sub(gen_p_i_10_io_x_sub),
    .io_sel(gen_p_i_10_io_sel),
    .io_p(gen_p_i_10_io_p)
  );
  gen_p_i gen_p_i_11 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_11_io_x),
    .io_x_sub(gen_p_i_11_io_x_sub),
    .io_sel(gen_p_i_11_io_sel),
    .io_p(gen_p_i_11_io_p)
  );
  gen_p_i gen_p_i_12 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_12_io_x),
    .io_x_sub(gen_p_i_12_io_x_sub),
    .io_sel(gen_p_i_12_io_sel),
    .io_p(gen_p_i_12_io_p)
  );
  gen_p_i gen_p_i_13 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_13_io_x),
    .io_x_sub(gen_p_i_13_io_x_sub),
    .io_sel(gen_p_i_13_io_sel),
    .io_p(gen_p_i_13_io_p)
  );
  gen_p_i gen_p_i_14 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_14_io_x),
    .io_x_sub(gen_p_i_14_io_x_sub),
    .io_sel(gen_p_i_14_io_sel),
    .io_p(gen_p_i_14_io_p)
  );
  gen_p_i gen_p_i_15 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_15_io_x),
    .io_x_sub(gen_p_i_15_io_x_sub),
    .io_sel(gen_p_i_15_io_sel),
    .io_p(gen_p_i_15_io_p)
  );
  gen_p_i gen_p_i_16 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_16_io_x),
    .io_x_sub(gen_p_i_16_io_x_sub),
    .io_sel(gen_p_i_16_io_sel),
    .io_p(gen_p_i_16_io_p)
  );
  gen_p_i gen_p_i_17 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_17_io_x),
    .io_x_sub(gen_p_i_17_io_x_sub),
    .io_sel(gen_p_i_17_io_sel),
    .io_p(gen_p_i_17_io_p)
  );
  gen_p_i gen_p_i_18 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_18_io_x),
    .io_x_sub(gen_p_i_18_io_x_sub),
    .io_sel(gen_p_i_18_io_sel),
    .io_p(gen_p_i_18_io_p)
  );
  gen_p_i gen_p_i_19 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_19_io_x),
    .io_x_sub(gen_p_i_19_io_x_sub),
    .io_sel(gen_p_i_19_io_sel),
    .io_p(gen_p_i_19_io_p)
  );
  gen_p_i gen_p_i_20 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_20_io_x),
    .io_x_sub(gen_p_i_20_io_x_sub),
    .io_sel(gen_p_i_20_io_sel),
    .io_p(gen_p_i_20_io_p)
  );
  gen_p_i gen_p_i_21 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_21_io_x),
    .io_x_sub(gen_p_i_21_io_x_sub),
    .io_sel(gen_p_i_21_io_sel),
    .io_p(gen_p_i_21_io_p)
  );
  gen_p_i gen_p_i_22 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_22_io_x),
    .io_x_sub(gen_p_i_22_io_x_sub),
    .io_sel(gen_p_i_22_io_sel),
    .io_p(gen_p_i_22_io_p)
  );
  gen_p_i gen_p_i_23 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_23_io_x),
    .io_x_sub(gen_p_i_23_io_x_sub),
    .io_sel(gen_p_i_23_io_sel),
    .io_p(gen_p_i_23_io_p)
  );
  gen_p_i gen_p_i_24 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_24_io_x),
    .io_x_sub(gen_p_i_24_io_x_sub),
    .io_sel(gen_p_i_24_io_sel),
    .io_p(gen_p_i_24_io_p)
  );
  gen_p_i gen_p_i_25 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_25_io_x),
    .io_x_sub(gen_p_i_25_io_x_sub),
    .io_sel(gen_p_i_25_io_sel),
    .io_p(gen_p_i_25_io_p)
  );
  gen_p_i gen_p_i_26 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_26_io_x),
    .io_x_sub(gen_p_i_26_io_x_sub),
    .io_sel(gen_p_i_26_io_sel),
    .io_p(gen_p_i_26_io_p)
  );
  gen_p_i gen_p_i_27 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_27_io_x),
    .io_x_sub(gen_p_i_27_io_x_sub),
    .io_sel(gen_p_i_27_io_sel),
    .io_p(gen_p_i_27_io_p)
  );
  gen_p_i gen_p_i_28 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_28_io_x),
    .io_x_sub(gen_p_i_28_io_x_sub),
    .io_sel(gen_p_i_28_io_sel),
    .io_p(gen_p_i_28_io_p)
  );
  gen_p_i gen_p_i_29 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_29_io_x),
    .io_x_sub(gen_p_i_29_io_x_sub),
    .io_sel(gen_p_i_29_io_sel),
    .io_p(gen_p_i_29_io_p)
  );
  gen_p_i gen_p_i_30 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_30_io_x),
    .io_x_sub(gen_p_i_30_io_x_sub),
    .io_sel(gen_p_i_30_io_sel),
    .io_p(gen_p_i_30_io_p)
  );
  gen_p_i gen_p_i_31 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_31_io_x),
    .io_x_sub(gen_p_i_31_io_x_sub),
    .io_sel(gen_p_i_31_io_sel),
    .io_p(gen_p_i_31_io_p)
  );
  gen_p_i gen_p_i_32 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_32_io_x),
    .io_x_sub(gen_p_i_32_io_x_sub),
    .io_sel(gen_p_i_32_io_sel),
    .io_p(gen_p_i_32_io_p)
  );
  gen_p_i gen_p_i_33 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_33_io_x),
    .io_x_sub(gen_p_i_33_io_x_sub),
    .io_sel(gen_p_i_33_io_sel),
    .io_p(gen_p_i_33_io_p)
  );
  gen_p_i gen_p_i_34 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_34_io_x),
    .io_x_sub(gen_p_i_34_io_x_sub),
    .io_sel(gen_p_i_34_io_sel),
    .io_p(gen_p_i_34_io_p)
  );
  gen_p_i gen_p_i_35 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_35_io_x),
    .io_x_sub(gen_p_i_35_io_x_sub),
    .io_sel(gen_p_i_35_io_sel),
    .io_p(gen_p_i_35_io_p)
  );
  gen_p_i gen_p_i_36 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_36_io_x),
    .io_x_sub(gen_p_i_36_io_x_sub),
    .io_sel(gen_p_i_36_io_sel),
    .io_p(gen_p_i_36_io_p)
  );
  gen_p_i gen_p_i_37 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_37_io_x),
    .io_x_sub(gen_p_i_37_io_x_sub),
    .io_sel(gen_p_i_37_io_sel),
    .io_p(gen_p_i_37_io_p)
  );
  gen_p_i gen_p_i_38 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_38_io_x),
    .io_x_sub(gen_p_i_38_io_x_sub),
    .io_sel(gen_p_i_38_io_sel),
    .io_p(gen_p_i_38_io_p)
  );
  gen_p_i gen_p_i_39 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_39_io_x),
    .io_x_sub(gen_p_i_39_io_x_sub),
    .io_sel(gen_p_i_39_io_sel),
    .io_p(gen_p_i_39_io_p)
  );
  gen_p_i gen_p_i_40 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_40_io_x),
    .io_x_sub(gen_p_i_40_io_x_sub),
    .io_sel(gen_p_i_40_io_sel),
    .io_p(gen_p_i_40_io_p)
  );
  gen_p_i gen_p_i_41 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_41_io_x),
    .io_x_sub(gen_p_i_41_io_x_sub),
    .io_sel(gen_p_i_41_io_sel),
    .io_p(gen_p_i_41_io_p)
  );
  gen_p_i gen_p_i_42 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_42_io_x),
    .io_x_sub(gen_p_i_42_io_x_sub),
    .io_sel(gen_p_i_42_io_sel),
    .io_p(gen_p_i_42_io_p)
  );
  gen_p_i gen_p_i_43 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_43_io_x),
    .io_x_sub(gen_p_i_43_io_x_sub),
    .io_sel(gen_p_i_43_io_sel),
    .io_p(gen_p_i_43_io_p)
  );
  gen_p_i gen_p_i_44 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_44_io_x),
    .io_x_sub(gen_p_i_44_io_x_sub),
    .io_sel(gen_p_i_44_io_sel),
    .io_p(gen_p_i_44_io_p)
  );
  gen_p_i gen_p_i_45 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_45_io_x),
    .io_x_sub(gen_p_i_45_io_x_sub),
    .io_sel(gen_p_i_45_io_sel),
    .io_p(gen_p_i_45_io_p)
  );
  gen_p_i gen_p_i_46 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_46_io_x),
    .io_x_sub(gen_p_i_46_io_x_sub),
    .io_sel(gen_p_i_46_io_sel),
    .io_p(gen_p_i_46_io_p)
  );
  gen_p_i gen_p_i_47 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_47_io_x),
    .io_x_sub(gen_p_i_47_io_x_sub),
    .io_sel(gen_p_i_47_io_sel),
    .io_p(gen_p_i_47_io_p)
  );
  gen_p_i gen_p_i_48 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_48_io_x),
    .io_x_sub(gen_p_i_48_io_x_sub),
    .io_sel(gen_p_i_48_io_sel),
    .io_p(gen_p_i_48_io_p)
  );
  gen_p_i gen_p_i_49 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_49_io_x),
    .io_x_sub(gen_p_i_49_io_x_sub),
    .io_sel(gen_p_i_49_io_sel),
    .io_p(gen_p_i_49_io_p)
  );
  gen_p_i gen_p_i_50 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_50_io_x),
    .io_x_sub(gen_p_i_50_io_x_sub),
    .io_sel(gen_p_i_50_io_sel),
    .io_p(gen_p_i_50_io_p)
  );
  gen_p_i gen_p_i_51 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_51_io_x),
    .io_x_sub(gen_p_i_51_io_x_sub),
    .io_sel(gen_p_i_51_io_sel),
    .io_p(gen_p_i_51_io_p)
  );
  gen_p_i gen_p_i_52 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_52_io_x),
    .io_x_sub(gen_p_i_52_io_x_sub),
    .io_sel(gen_p_i_52_io_sel),
    .io_p(gen_p_i_52_io_p)
  );
  gen_p_i gen_p_i_53 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_53_io_x),
    .io_x_sub(gen_p_i_53_io_x_sub),
    .io_sel(gen_p_i_53_io_sel),
    .io_p(gen_p_i_53_io_p)
  );
  gen_p_i gen_p_i_54 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_54_io_x),
    .io_x_sub(gen_p_i_54_io_x_sub),
    .io_sel(gen_p_i_54_io_sel),
    .io_p(gen_p_i_54_io_p)
  );
  gen_p_i gen_p_i_55 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_55_io_x),
    .io_x_sub(gen_p_i_55_io_x_sub),
    .io_sel(gen_p_i_55_io_sel),
    .io_p(gen_p_i_55_io_p)
  );
  gen_p_i gen_p_i_56 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_56_io_x),
    .io_x_sub(gen_p_i_56_io_x_sub),
    .io_sel(gen_p_i_56_io_sel),
    .io_p(gen_p_i_56_io_p)
  );
  gen_p_i gen_p_i_57 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_57_io_x),
    .io_x_sub(gen_p_i_57_io_x_sub),
    .io_sel(gen_p_i_57_io_sel),
    .io_p(gen_p_i_57_io_p)
  );
  gen_p_i gen_p_i_58 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_58_io_x),
    .io_x_sub(gen_p_i_58_io_x_sub),
    .io_sel(gen_p_i_58_io_sel),
    .io_p(gen_p_i_58_io_p)
  );
  gen_p_i gen_p_i_59 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_59_io_x),
    .io_x_sub(gen_p_i_59_io_x_sub),
    .io_sel(gen_p_i_59_io_sel),
    .io_p(gen_p_i_59_io_p)
  );
  gen_p_i gen_p_i_60 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_60_io_x),
    .io_x_sub(gen_p_i_60_io_x_sub),
    .io_sel(gen_p_i_60_io_sel),
    .io_p(gen_p_i_60_io_p)
  );
  gen_p_i gen_p_i_61 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_61_io_x),
    .io_x_sub(gen_p_i_61_io_x_sub),
    .io_sel(gen_p_i_61_io_sel),
    .io_p(gen_p_i_61_io_p)
  );
  gen_p_i gen_p_i_62 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_62_io_x),
    .io_x_sub(gen_p_i_62_io_x_sub),
    .io_sel(gen_p_i_62_io_sel),
    .io_p(gen_p_i_62_io_p)
  );
  gen_p_i gen_p_i_63 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_63_io_x),
    .io_x_sub(gen_p_i_63_io_x_sub),
    .io_sel(gen_p_i_63_io_sel),
    .io_p(gen_p_i_63_io_p)
  );
  gen_p_i gen_p_i_64 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_64_io_x),
    .io_x_sub(gen_p_i_64_io_x_sub),
    .io_sel(gen_p_i_64_io_sel),
    .io_p(gen_p_i_64_io_p)
  );
  gen_p_i gen_p_i_65 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_65_io_x),
    .io_x_sub(gen_p_i_65_io_x_sub),
    .io_sel(gen_p_i_65_io_sel),
    .io_p(gen_p_i_65_io_p)
  );
  gen_p_i gen_p_i_66 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_66_io_x),
    .io_x_sub(gen_p_i_66_io_x_sub),
    .io_sel(gen_p_i_66_io_sel),
    .io_p(gen_p_i_66_io_p)
  );
  gen_p_i gen_p_i_67 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_67_io_x),
    .io_x_sub(gen_p_i_67_io_x_sub),
    .io_sel(gen_p_i_67_io_sel),
    .io_p(gen_p_i_67_io_p)
  );
  gen_p_i gen_p_i_68 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_68_io_x),
    .io_x_sub(gen_p_i_68_io_x_sub),
    .io_sel(gen_p_i_68_io_sel),
    .io_p(gen_p_i_68_io_p)
  );
  gen_p_i gen_p_i_69 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_69_io_x),
    .io_x_sub(gen_p_i_69_io_x_sub),
    .io_sel(gen_p_i_69_io_sel),
    .io_p(gen_p_i_69_io_p)
  );
  gen_p_i gen_p_i_70 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_70_io_x),
    .io_x_sub(gen_p_i_70_io_x_sub),
    .io_sel(gen_p_i_70_io_sel),
    .io_p(gen_p_i_70_io_p)
  );
  gen_p_i gen_p_i_71 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_71_io_x),
    .io_x_sub(gen_p_i_71_io_x_sub),
    .io_sel(gen_p_i_71_io_sel),
    .io_p(gen_p_i_71_io_p)
  );
  gen_p_i gen_p_i_72 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_72_io_x),
    .io_x_sub(gen_p_i_72_io_x_sub),
    .io_sel(gen_p_i_72_io_sel),
    .io_p(gen_p_i_72_io_p)
  );
  gen_p_i gen_p_i_73 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_73_io_x),
    .io_x_sub(gen_p_i_73_io_x_sub),
    .io_sel(gen_p_i_73_io_sel),
    .io_p(gen_p_i_73_io_p)
  );
  gen_p_i gen_p_i_74 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_74_io_x),
    .io_x_sub(gen_p_i_74_io_x_sub),
    .io_sel(gen_p_i_74_io_sel),
    .io_p(gen_p_i_74_io_p)
  );
  gen_p_i gen_p_i_75 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_75_io_x),
    .io_x_sub(gen_p_i_75_io_x_sub),
    .io_sel(gen_p_i_75_io_sel),
    .io_p(gen_p_i_75_io_p)
  );
  gen_p_i gen_p_i_76 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_76_io_x),
    .io_x_sub(gen_p_i_76_io_x_sub),
    .io_sel(gen_p_i_76_io_sel),
    .io_p(gen_p_i_76_io_p)
  );
  gen_p_i gen_p_i_77 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_77_io_x),
    .io_x_sub(gen_p_i_77_io_x_sub),
    .io_sel(gen_p_i_77_io_sel),
    .io_p(gen_p_i_77_io_p)
  );
  gen_p_i gen_p_i_78 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_78_io_x),
    .io_x_sub(gen_p_i_78_io_x_sub),
    .io_sel(gen_p_i_78_io_sel),
    .io_p(gen_p_i_78_io_p)
  );
  gen_p_i gen_p_i_79 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_79_io_x),
    .io_x_sub(gen_p_i_79_io_x_sub),
    .io_sel(gen_p_i_79_io_sel),
    .io_p(gen_p_i_79_io_p)
  );
  gen_p_i gen_p_i_80 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_80_io_x),
    .io_x_sub(gen_p_i_80_io_x_sub),
    .io_sel(gen_p_i_80_io_sel),
    .io_p(gen_p_i_80_io_p)
  );
  gen_p_i gen_p_i_81 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_81_io_x),
    .io_x_sub(gen_p_i_81_io_x_sub),
    .io_sel(gen_p_i_81_io_sel),
    .io_p(gen_p_i_81_io_p)
  );
  gen_p_i gen_p_i_82 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_82_io_x),
    .io_x_sub(gen_p_i_82_io_x_sub),
    .io_sel(gen_p_i_82_io_sel),
    .io_p(gen_p_i_82_io_p)
  );
  gen_p_i gen_p_i_83 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_83_io_x),
    .io_x_sub(gen_p_i_83_io_x_sub),
    .io_sel(gen_p_i_83_io_sel),
    .io_p(gen_p_i_83_io_p)
  );
  gen_p_i gen_p_i_84 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_84_io_x),
    .io_x_sub(gen_p_i_84_io_x_sub),
    .io_sel(gen_p_i_84_io_sel),
    .io_p(gen_p_i_84_io_p)
  );
  gen_p_i gen_p_i_85 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_85_io_x),
    .io_x_sub(gen_p_i_85_io_x_sub),
    .io_sel(gen_p_i_85_io_sel),
    .io_p(gen_p_i_85_io_p)
  );
  gen_p_i gen_p_i_86 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_86_io_x),
    .io_x_sub(gen_p_i_86_io_x_sub),
    .io_sel(gen_p_i_86_io_sel),
    .io_p(gen_p_i_86_io_p)
  );
  gen_p_i gen_p_i_87 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_87_io_x),
    .io_x_sub(gen_p_i_87_io_x_sub),
    .io_sel(gen_p_i_87_io_sel),
    .io_p(gen_p_i_87_io_p)
  );
  gen_p_i gen_p_i_88 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_88_io_x),
    .io_x_sub(gen_p_i_88_io_x_sub),
    .io_sel(gen_p_i_88_io_sel),
    .io_p(gen_p_i_88_io_p)
  );
  gen_p_i gen_p_i_89 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_89_io_x),
    .io_x_sub(gen_p_i_89_io_x_sub),
    .io_sel(gen_p_i_89_io_sel),
    .io_p(gen_p_i_89_io_p)
  );
  gen_p_i gen_p_i_90 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_90_io_x),
    .io_x_sub(gen_p_i_90_io_x_sub),
    .io_sel(gen_p_i_90_io_sel),
    .io_p(gen_p_i_90_io_p)
  );
  gen_p_i gen_p_i_91 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_91_io_x),
    .io_x_sub(gen_p_i_91_io_x_sub),
    .io_sel(gen_p_i_91_io_sel),
    .io_p(gen_p_i_91_io_p)
  );
  gen_p_i gen_p_i_92 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_92_io_x),
    .io_x_sub(gen_p_i_92_io_x_sub),
    .io_sel(gen_p_i_92_io_sel),
    .io_p(gen_p_i_92_io_p)
  );
  gen_p_i gen_p_i_93 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_93_io_x),
    .io_x_sub(gen_p_i_93_io_x_sub),
    .io_sel(gen_p_i_93_io_sel),
    .io_p(gen_p_i_93_io_p)
  );
  gen_p_i gen_p_i_94 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_94_io_x),
    .io_x_sub(gen_p_i_94_io_x_sub),
    .io_sel(gen_p_i_94_io_sel),
    .io_p(gen_p_i_94_io_p)
  );
  gen_p_i gen_p_i_95 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_95_io_x),
    .io_x_sub(gen_p_i_95_io_x_sub),
    .io_sel(gen_p_i_95_io_sel),
    .io_p(gen_p_i_95_io_p)
  );
  gen_p_i gen_p_i_96 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_96_io_x),
    .io_x_sub(gen_p_i_96_io_x_sub),
    .io_sel(gen_p_i_96_io_sel),
    .io_p(gen_p_i_96_io_p)
  );
  gen_p_i gen_p_i_97 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_97_io_x),
    .io_x_sub(gen_p_i_97_io_x_sub),
    .io_sel(gen_p_i_97_io_sel),
    .io_p(gen_p_i_97_io_p)
  );
  gen_p_i gen_p_i_98 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_98_io_x),
    .io_x_sub(gen_p_i_98_io_x_sub),
    .io_sel(gen_p_i_98_io_sel),
    .io_p(gen_p_i_98_io_p)
  );
  gen_p_i gen_p_i_99 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_99_io_x),
    .io_x_sub(gen_p_i_99_io_x_sub),
    .io_sel(gen_p_i_99_io_sel),
    .io_p(gen_p_i_99_io_p)
  );
  gen_p_i gen_p_i_100 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_100_io_x),
    .io_x_sub(gen_p_i_100_io_x_sub),
    .io_sel(gen_p_i_100_io_sel),
    .io_p(gen_p_i_100_io_p)
  );
  gen_p_i gen_p_i_101 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_101_io_x),
    .io_x_sub(gen_p_i_101_io_x_sub),
    .io_sel(gen_p_i_101_io_sel),
    .io_p(gen_p_i_101_io_p)
  );
  gen_p_i gen_p_i_102 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_102_io_x),
    .io_x_sub(gen_p_i_102_io_x_sub),
    .io_sel(gen_p_i_102_io_sel),
    .io_p(gen_p_i_102_io_p)
  );
  gen_p_i gen_p_i_103 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_103_io_x),
    .io_x_sub(gen_p_i_103_io_x_sub),
    .io_sel(gen_p_i_103_io_sel),
    .io_p(gen_p_i_103_io_p)
  );
  gen_p_i gen_p_i_104 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_104_io_x),
    .io_x_sub(gen_p_i_104_io_x_sub),
    .io_sel(gen_p_i_104_io_sel),
    .io_p(gen_p_i_104_io_p)
  );
  gen_p_i gen_p_i_105 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_105_io_x),
    .io_x_sub(gen_p_i_105_io_x_sub),
    .io_sel(gen_p_i_105_io_sel),
    .io_p(gen_p_i_105_io_p)
  );
  gen_p_i gen_p_i_106 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_106_io_x),
    .io_x_sub(gen_p_i_106_io_x_sub),
    .io_sel(gen_p_i_106_io_sel),
    .io_p(gen_p_i_106_io_p)
  );
  gen_p_i gen_p_i_107 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_107_io_x),
    .io_x_sub(gen_p_i_107_io_x_sub),
    .io_sel(gen_p_i_107_io_sel),
    .io_p(gen_p_i_107_io_p)
  );
  gen_p_i gen_p_i_108 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_108_io_x),
    .io_x_sub(gen_p_i_108_io_x_sub),
    .io_sel(gen_p_i_108_io_sel),
    .io_p(gen_p_i_108_io_p)
  );
  gen_p_i gen_p_i_109 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_109_io_x),
    .io_x_sub(gen_p_i_109_io_x_sub),
    .io_sel(gen_p_i_109_io_sel),
    .io_p(gen_p_i_109_io_p)
  );
  gen_p_i gen_p_i_110 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_110_io_x),
    .io_x_sub(gen_p_i_110_io_x_sub),
    .io_sel(gen_p_i_110_io_sel),
    .io_p(gen_p_i_110_io_p)
  );
  gen_p_i gen_p_i_111 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_111_io_x),
    .io_x_sub(gen_p_i_111_io_x_sub),
    .io_sel(gen_p_i_111_io_sel),
    .io_p(gen_p_i_111_io_p)
  );
  gen_p_i gen_p_i_112 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_112_io_x),
    .io_x_sub(gen_p_i_112_io_x_sub),
    .io_sel(gen_p_i_112_io_sel),
    .io_p(gen_p_i_112_io_p)
  );
  gen_p_i gen_p_i_113 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_113_io_x),
    .io_x_sub(gen_p_i_113_io_x_sub),
    .io_sel(gen_p_i_113_io_sel),
    .io_p(gen_p_i_113_io_p)
  );
  gen_p_i gen_p_i_114 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_114_io_x),
    .io_x_sub(gen_p_i_114_io_x_sub),
    .io_sel(gen_p_i_114_io_sel),
    .io_p(gen_p_i_114_io_p)
  );
  gen_p_i gen_p_i_115 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_115_io_x),
    .io_x_sub(gen_p_i_115_io_x_sub),
    .io_sel(gen_p_i_115_io_sel),
    .io_p(gen_p_i_115_io_p)
  );
  gen_p_i gen_p_i_116 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_116_io_x),
    .io_x_sub(gen_p_i_116_io_x_sub),
    .io_sel(gen_p_i_116_io_sel),
    .io_p(gen_p_i_116_io_p)
  );
  gen_p_i gen_p_i_117 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_117_io_x),
    .io_x_sub(gen_p_i_117_io_x_sub),
    .io_sel(gen_p_i_117_io_sel),
    .io_p(gen_p_i_117_io_p)
  );
  gen_p_i gen_p_i_118 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_118_io_x),
    .io_x_sub(gen_p_i_118_io_x_sub),
    .io_sel(gen_p_i_118_io_sel),
    .io_p(gen_p_i_118_io_p)
  );
  gen_p_i gen_p_i_119 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_119_io_x),
    .io_x_sub(gen_p_i_119_io_x_sub),
    .io_sel(gen_p_i_119_io_sel),
    .io_p(gen_p_i_119_io_p)
  );
  gen_p_i gen_p_i_120 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_120_io_x),
    .io_x_sub(gen_p_i_120_io_x_sub),
    .io_sel(gen_p_i_120_io_sel),
    .io_p(gen_p_i_120_io_p)
  );
  gen_p_i gen_p_i_121 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_121_io_x),
    .io_x_sub(gen_p_i_121_io_x_sub),
    .io_sel(gen_p_i_121_io_sel),
    .io_p(gen_p_i_121_io_p)
  );
  gen_p_i gen_p_i_122 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_122_io_x),
    .io_x_sub(gen_p_i_122_io_x_sub),
    .io_sel(gen_p_i_122_io_sel),
    .io_p(gen_p_i_122_io_p)
  );
  gen_p_i gen_p_i_123 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_123_io_x),
    .io_x_sub(gen_p_i_123_io_x_sub),
    .io_sel(gen_p_i_123_io_sel),
    .io_p(gen_p_i_123_io_p)
  );
  gen_p_i gen_p_i_124 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_124_io_x),
    .io_x_sub(gen_p_i_124_io_x_sub),
    .io_sel(gen_p_i_124_io_sel),
    .io_p(gen_p_i_124_io_p)
  );
  gen_p_i gen_p_i_125 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_125_io_x),
    .io_x_sub(gen_p_i_125_io_x_sub),
    .io_sel(gen_p_i_125_io_sel),
    .io_p(gen_p_i_125_io_p)
  );
  gen_p_i gen_p_i_126 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_126_io_x),
    .io_x_sub(gen_p_i_126_io_x_sub),
    .io_sel(gen_p_i_126_io_sel),
    .io_p(gen_p_i_126_io_p)
  );
  gen_p_i gen_p_i_127 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_127_io_x),
    .io_x_sub(gen_p_i_127_io_x_sub),
    .io_sel(gen_p_i_127_io_sel),
    .io_p(gen_p_i_127_io_p)
  );
  gen_p_i gen_p_i_128 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_128_io_x),
    .io_x_sub(gen_p_i_128_io_x_sub),
    .io_sel(gen_p_i_128_io_sel),
    .io_p(gen_p_i_128_io_p)
  );
  gen_p_i gen_p_i_129 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_129_io_x),
    .io_x_sub(gen_p_i_129_io_x_sub),
    .io_sel(gen_p_i_129_io_sel),
    .io_p(gen_p_i_129_io_p)
  );
  gen_p_i gen_p_i_130 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_130_io_x),
    .io_x_sub(gen_p_i_130_io_x_sub),
    .io_sel(gen_p_i_130_io_sel),
    .io_p(gen_p_i_130_io_p)
  );
  gen_p_i gen_p_i_131 ( // @[WallaceTest.scala 76:29]
    .io_x(gen_p_i_131_io_x),
    .io_x_sub(gen_p_i_131_io_x_sub),
    .io_sel(gen_p_i_131_io_sel),
    .io_p(gen_p_i_131_io_p)
  );
  assign io_p = {io_p_hi,io_p_lo}; // @[Cat.scala 33:92]
  assign io_c = gen_sel_io_out[0] | gen_sel_io_out[2]; // @[WallaceTest.scala 92:21]
  assign gen_sel_io_src = io_src; // @[WallaceTest.scala 78:10]
  assign gen_p_i_io_x = io_x[0]; // @[WallaceTest.scala 80:16]
  assign gen_p_i_io_x_sub = 1'h0; // @[WallaceTest.scala 81:14]
  assign gen_p_i_io_sel = gen_sel_io_out; // @[WallaceTest.scala 82:11]
  assign gen_p_i_1_io_x = io_x[1]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_1_io_x_sub = io_x[0]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_1_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_2_io_x = io_x[2]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_2_io_x_sub = io_x[1]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_2_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_3_io_x = io_x[3]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_3_io_x_sub = io_x[2]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_3_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_4_io_x = io_x[4]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_4_io_x_sub = io_x[3]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_4_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_5_io_x = io_x[5]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_5_io_x_sub = io_x[4]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_5_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_6_io_x = io_x[6]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_6_io_x_sub = io_x[5]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_6_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_7_io_x = io_x[7]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_7_io_x_sub = io_x[6]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_7_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_8_io_x = io_x[8]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_8_io_x_sub = io_x[7]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_8_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_9_io_x = io_x[9]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_9_io_x_sub = io_x[8]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_9_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_10_io_x = io_x[10]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_10_io_x_sub = io_x[9]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_10_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_11_io_x = io_x[11]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_11_io_x_sub = io_x[10]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_11_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_12_io_x = io_x[12]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_12_io_x_sub = io_x[11]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_12_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_13_io_x = io_x[13]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_13_io_x_sub = io_x[12]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_13_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_14_io_x = io_x[14]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_14_io_x_sub = io_x[13]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_14_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_15_io_x = io_x[15]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_15_io_x_sub = io_x[14]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_15_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_16_io_x = io_x[16]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_16_io_x_sub = io_x[15]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_16_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_17_io_x = io_x[17]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_17_io_x_sub = io_x[16]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_17_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_18_io_x = io_x[18]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_18_io_x_sub = io_x[17]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_18_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_19_io_x = io_x[19]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_19_io_x_sub = io_x[18]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_19_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_20_io_x = io_x[20]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_20_io_x_sub = io_x[19]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_20_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_21_io_x = io_x[21]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_21_io_x_sub = io_x[20]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_21_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_22_io_x = io_x[22]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_22_io_x_sub = io_x[21]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_22_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_23_io_x = io_x[23]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_23_io_x_sub = io_x[22]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_23_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_24_io_x = io_x[24]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_24_io_x_sub = io_x[23]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_24_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_25_io_x = io_x[25]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_25_io_x_sub = io_x[24]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_25_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_26_io_x = io_x[26]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_26_io_x_sub = io_x[25]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_26_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_27_io_x = io_x[27]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_27_io_x_sub = io_x[26]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_27_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_28_io_x = io_x[28]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_28_io_x_sub = io_x[27]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_28_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_29_io_x = io_x[29]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_29_io_x_sub = io_x[28]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_29_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_30_io_x = io_x[30]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_30_io_x_sub = io_x[29]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_30_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_31_io_x = io_x[31]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_31_io_x_sub = io_x[30]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_31_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_32_io_x = io_x[32]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_32_io_x_sub = io_x[31]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_32_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_33_io_x = io_x[33]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_33_io_x_sub = io_x[32]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_33_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_34_io_x = io_x[34]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_34_io_x_sub = io_x[33]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_34_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_35_io_x = io_x[35]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_35_io_x_sub = io_x[34]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_35_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_36_io_x = io_x[36]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_36_io_x_sub = io_x[35]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_36_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_37_io_x = io_x[37]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_37_io_x_sub = io_x[36]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_37_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_38_io_x = io_x[38]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_38_io_x_sub = io_x[37]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_38_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_39_io_x = io_x[39]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_39_io_x_sub = io_x[38]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_39_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_40_io_x = io_x[40]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_40_io_x_sub = io_x[39]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_40_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_41_io_x = io_x[41]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_41_io_x_sub = io_x[40]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_41_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_42_io_x = io_x[42]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_42_io_x_sub = io_x[41]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_42_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_43_io_x = io_x[43]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_43_io_x_sub = io_x[42]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_43_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_44_io_x = io_x[44]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_44_io_x_sub = io_x[43]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_44_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_45_io_x = io_x[45]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_45_io_x_sub = io_x[44]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_45_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_46_io_x = io_x[46]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_46_io_x_sub = io_x[45]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_46_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_47_io_x = io_x[47]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_47_io_x_sub = io_x[46]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_47_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_48_io_x = io_x[48]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_48_io_x_sub = io_x[47]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_48_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_49_io_x = io_x[49]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_49_io_x_sub = io_x[48]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_49_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_50_io_x = io_x[50]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_50_io_x_sub = io_x[49]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_50_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_51_io_x = io_x[51]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_51_io_x_sub = io_x[50]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_51_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_52_io_x = io_x[52]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_52_io_x_sub = io_x[51]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_52_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_53_io_x = io_x[53]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_53_io_x_sub = io_x[52]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_53_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_54_io_x = io_x[54]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_54_io_x_sub = io_x[53]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_54_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_55_io_x = io_x[55]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_55_io_x_sub = io_x[54]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_55_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_56_io_x = io_x[56]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_56_io_x_sub = io_x[55]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_56_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_57_io_x = io_x[57]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_57_io_x_sub = io_x[56]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_57_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_58_io_x = io_x[58]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_58_io_x_sub = io_x[57]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_58_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_59_io_x = io_x[59]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_59_io_x_sub = io_x[58]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_59_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_60_io_x = io_x[60]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_60_io_x_sub = io_x[59]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_60_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_61_io_x = io_x[61]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_61_io_x_sub = io_x[60]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_61_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_62_io_x = io_x[62]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_62_io_x_sub = io_x[61]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_62_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_63_io_x = io_x[63]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_63_io_x_sub = io_x[62]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_63_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_64_io_x = io_x[64]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_64_io_x_sub = io_x[63]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_64_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_65_io_x = io_x[65]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_65_io_x_sub = io_x[64]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_65_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_66_io_x = io_x[66]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_66_io_x_sub = io_x[65]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_66_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_67_io_x = io_x[67]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_67_io_x_sub = io_x[66]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_67_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_68_io_x = io_x[68]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_68_io_x_sub = io_x[67]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_68_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_69_io_x = io_x[69]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_69_io_x_sub = io_x[68]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_69_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_70_io_x = io_x[70]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_70_io_x_sub = io_x[69]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_70_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_71_io_x = io_x[71]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_71_io_x_sub = io_x[70]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_71_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_72_io_x = io_x[72]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_72_io_x_sub = io_x[71]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_72_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_73_io_x = io_x[73]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_73_io_x_sub = io_x[72]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_73_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_74_io_x = io_x[74]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_74_io_x_sub = io_x[73]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_74_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_75_io_x = io_x[75]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_75_io_x_sub = io_x[74]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_75_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_76_io_x = io_x[76]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_76_io_x_sub = io_x[75]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_76_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_77_io_x = io_x[77]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_77_io_x_sub = io_x[76]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_77_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_78_io_x = io_x[78]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_78_io_x_sub = io_x[77]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_78_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_79_io_x = io_x[79]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_79_io_x_sub = io_x[78]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_79_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_80_io_x = io_x[80]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_80_io_x_sub = io_x[79]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_80_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_81_io_x = io_x[81]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_81_io_x_sub = io_x[80]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_81_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_82_io_x = io_x[82]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_82_io_x_sub = io_x[81]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_82_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_83_io_x = io_x[83]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_83_io_x_sub = io_x[82]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_83_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_84_io_x = io_x[84]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_84_io_x_sub = io_x[83]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_84_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_85_io_x = io_x[85]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_85_io_x_sub = io_x[84]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_85_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_86_io_x = io_x[86]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_86_io_x_sub = io_x[85]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_86_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_87_io_x = io_x[87]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_87_io_x_sub = io_x[86]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_87_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_88_io_x = io_x[88]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_88_io_x_sub = io_x[87]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_88_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_89_io_x = io_x[89]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_89_io_x_sub = io_x[88]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_89_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_90_io_x = io_x[90]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_90_io_x_sub = io_x[89]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_90_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_91_io_x = io_x[91]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_91_io_x_sub = io_x[90]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_91_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_92_io_x = io_x[92]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_92_io_x_sub = io_x[91]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_92_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_93_io_x = io_x[93]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_93_io_x_sub = io_x[92]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_93_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_94_io_x = io_x[94]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_94_io_x_sub = io_x[93]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_94_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_95_io_x = io_x[95]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_95_io_x_sub = io_x[94]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_95_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_96_io_x = io_x[96]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_96_io_x_sub = io_x[95]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_96_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_97_io_x = io_x[97]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_97_io_x_sub = io_x[96]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_97_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_98_io_x = io_x[98]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_98_io_x_sub = io_x[97]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_98_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_99_io_x = io_x[99]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_99_io_x_sub = io_x[98]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_99_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_100_io_x = io_x[100]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_100_io_x_sub = io_x[99]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_100_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_101_io_x = io_x[101]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_101_io_x_sub = io_x[100]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_101_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_102_io_x = io_x[102]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_102_io_x_sub = io_x[101]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_102_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_103_io_x = io_x[103]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_103_io_x_sub = io_x[102]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_103_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_104_io_x = io_x[104]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_104_io_x_sub = io_x[103]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_104_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_105_io_x = io_x[105]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_105_io_x_sub = io_x[104]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_105_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_106_io_x = io_x[106]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_106_io_x_sub = io_x[105]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_106_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_107_io_x = io_x[107]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_107_io_x_sub = io_x[106]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_107_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_108_io_x = io_x[108]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_108_io_x_sub = io_x[107]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_108_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_109_io_x = io_x[109]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_109_io_x_sub = io_x[108]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_109_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_110_io_x = io_x[110]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_110_io_x_sub = io_x[109]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_110_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_111_io_x = io_x[111]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_111_io_x_sub = io_x[110]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_111_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_112_io_x = io_x[112]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_112_io_x_sub = io_x[111]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_112_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_113_io_x = io_x[113]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_113_io_x_sub = io_x[112]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_113_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_114_io_x = io_x[114]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_114_io_x_sub = io_x[113]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_114_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_115_io_x = io_x[115]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_115_io_x_sub = io_x[114]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_115_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_116_io_x = io_x[116]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_116_io_x_sub = io_x[115]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_116_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_117_io_x = io_x[117]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_117_io_x_sub = io_x[116]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_117_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_118_io_x = io_x[118]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_118_io_x_sub = io_x[117]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_118_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_119_io_x = io_x[119]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_119_io_x_sub = io_x[118]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_119_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_120_io_x = io_x[120]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_120_io_x_sub = io_x[119]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_120_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_121_io_x = io_x[121]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_121_io_x_sub = io_x[120]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_121_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_122_io_x = io_x[122]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_122_io_x_sub = io_x[121]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_122_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_123_io_x = io_x[123]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_123_io_x_sub = io_x[122]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_123_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_124_io_x = io_x[124]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_124_io_x_sub = io_x[123]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_124_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_125_io_x = io_x[125]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_125_io_x_sub = io_x[124]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_125_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_126_io_x = io_x[126]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_126_io_x_sub = io_x[125]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_126_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_127_io_x = io_x[127]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_127_io_x_sub = io_x[126]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_127_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_128_io_x = io_x[128]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_128_io_x_sub = io_x[127]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_128_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_129_io_x = io_x[129]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_129_io_x_sub = io_x[128]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_129_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_130_io_x = io_x[130]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_130_io_x_sub = io_x[129]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_130_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
  assign gen_p_i_131_io_x = io_x[131]; // @[WallaceTest.scala 85:18]
  assign gen_p_i_131_io_x_sub = io_x[130]; // @[WallaceTest.scala 86:23]
  assign gen_p_i_131_io_sel = gen_sel_io_out; // @[WallaceTest.scala 87:13]
endmodule
module switch(
  input          clock,
  input          reset,
  input  [131:0] io_in_0,
  input  [131:0] io_in_1,
  input  [131:0] io_in_2,
  input  [131:0] io_in_3,
  input  [131:0] io_in_4,
  input  [131:0] io_in_5,
  input  [131:0] io_in_6,
  input  [131:0] io_in_7,
  input  [131:0] io_in_8,
  input  [131:0] io_in_9,
  input  [131:0] io_in_10,
  input  [131:0] io_in_11,
  input  [131:0] io_in_12,
  input  [131:0] io_in_13,
  input  [131:0] io_in_14,
  input  [131:0] io_in_15,
  input  [131:0] io_in_16,
  input  [131:0] io_in_17,
  input  [131:0] io_in_18,
  input  [131:0] io_in_19,
  input  [131:0] io_in_20,
  input  [131:0] io_in_21,
  input  [131:0] io_in_22,
  input  [131:0] io_in_23,
  input  [131:0] io_in_24,
  input  [131:0] io_in_25,
  input  [131:0] io_in_26,
  input  [131:0] io_in_27,
  input  [131:0] io_in_28,
  input  [131:0] io_in_29,
  input  [131:0] io_in_30,
  input  [131:0] io_in_31,
  input  [131:0] io_in_32,
  output [32:0]  io_out_0,
  output [32:0]  io_out_1,
  output [32:0]  io_out_2,
  output [32:0]  io_out_3,
  output [32:0]  io_out_4,
  output [32:0]  io_out_5,
  output [32:0]  io_out_6,
  output [32:0]  io_out_7,
  output [32:0]  io_out_8,
  output [32:0]  io_out_9,
  output [32:0]  io_out_10,
  output [32:0]  io_out_11,
  output [32:0]  io_out_12,
  output [32:0]  io_out_13,
  output [32:0]  io_out_14,
  output [32:0]  io_out_15,
  output [32:0]  io_out_16,
  output [32:0]  io_out_17,
  output [32:0]  io_out_18,
  output [32:0]  io_out_19,
  output [32:0]  io_out_20,
  output [32:0]  io_out_21,
  output [32:0]  io_out_22,
  output [32:0]  io_out_23,
  output [32:0]  io_out_24,
  output [32:0]  io_out_25,
  output [32:0]  io_out_26,
  output [32:0]  io_out_27,
  output [32:0]  io_out_28,
  output [32:0]  io_out_29,
  output [32:0]  io_out_30,
  output [32:0]  io_out_31,
  output [32:0]  io_out_32,
  output [32:0]  io_out_33,
  output [32:0]  io_out_34,
  output [32:0]  io_out_35,
  output [32:0]  io_out_36,
  output [32:0]  io_out_37,
  output [32:0]  io_out_38,
  output [32:0]  io_out_39,
  output [32:0]  io_out_40,
  output [32:0]  io_out_41,
  output [32:0]  io_out_42,
  output [32:0]  io_out_43,
  output [32:0]  io_out_44,
  output [32:0]  io_out_45,
  output [32:0]  io_out_46,
  output [32:0]  io_out_47,
  output [32:0]  io_out_48,
  output [32:0]  io_out_49,
  output [32:0]  io_out_50,
  output [32:0]  io_out_51,
  output [32:0]  io_out_52,
  output [32:0]  io_out_53,
  output [32:0]  io_out_54,
  output [32:0]  io_out_55,
  output [32:0]  io_out_56,
  output [32:0]  io_out_57,
  output [32:0]  io_out_58,
  output [32:0]  io_out_59,
  output [32:0]  io_out_60,
  output [32:0]  io_out_61,
  output [32:0]  io_out_62,
  output [32:0]  io_out_63,
  output [32:0]  io_out_64,
  output [32:0]  io_out_65,
  output [32:0]  io_out_66,
  output [32:0]  io_out_67,
  output [32:0]  io_out_68,
  output [32:0]  io_out_69,
  output [32:0]  io_out_70,
  output [32:0]  io_out_71,
  output [32:0]  io_out_72,
  output [32:0]  io_out_73,
  output [32:0]  io_out_74,
  output [32:0]  io_out_75,
  output [32:0]  io_out_76,
  output [32:0]  io_out_77,
  output [32:0]  io_out_78,
  output [32:0]  io_out_79,
  output [32:0]  io_out_80,
  output [32:0]  io_out_81,
  output [32:0]  io_out_82,
  output [32:0]  io_out_83,
  output [32:0]  io_out_84,
  output [32:0]  io_out_85,
  output [32:0]  io_out_86,
  output [32:0]  io_out_87,
  output [32:0]  io_out_88,
  output [32:0]  io_out_89,
  output [32:0]  io_out_90,
  output [32:0]  io_out_91,
  output [32:0]  io_out_92,
  output [32:0]  io_out_93,
  output [32:0]  io_out_94,
  output [32:0]  io_out_95,
  output [32:0]  io_out_96,
  output [32:0]  io_out_97,
  output [32:0]  io_out_98,
  output [32:0]  io_out_99,
  output [32:0]  io_out_100,
  output [32:0]  io_out_101,
  output [32:0]  io_out_102,
  output [32:0]  io_out_103,
  output [32:0]  io_out_104,
  output [32:0]  io_out_105,
  output [32:0]  io_out_106,
  output [32:0]  io_out_107,
  output [32:0]  io_out_108,
  output [32:0]  io_out_109,
  output [32:0]  io_out_110,
  output [32:0]  io_out_111,
  output [32:0]  io_out_112,
  output [32:0]  io_out_113,
  output [32:0]  io_out_114,
  output [32:0]  io_out_115,
  output [32:0]  io_out_116,
  output [32:0]  io_out_117,
  output [32:0]  io_out_118,
  output [32:0]  io_out_119,
  output [32:0]  io_out_120,
  output [32:0]  io_out_121,
  output [32:0]  io_out_122,
  output [32:0]  io_out_123,
  output [32:0]  io_out_124,
  output [32:0]  io_out_125,
  output [32:0]  io_out_126,
  output [32:0]  io_out_127,
  output [32:0]  io_out_128,
  output [32:0]  io_out_129,
  output [32:0]  io_out_130,
  output [32:0]  io_out_131,
  input          io_cin_0,
  input          io_cin_1,
  input          io_cin_2,
  input          io_cin_3,
  input          io_cin_4,
  input          io_cin_5,
  input          io_cin_6,
  input          io_cin_7,
  input          io_cin_8,
  input          io_cin_9,
  input          io_cin_10,
  input          io_cin_11,
  input          io_cin_12,
  input          io_cin_13,
  input          io_cin_14,
  input          io_cin_15,
  input          io_cin_16,
  input          io_cin_17,
  input          io_cin_18,
  input          io_cin_19,
  input          io_cin_20,
  input          io_cin_21,
  input          io_cin_22,
  input          io_cin_23,
  input          io_cin_24,
  input          io_cin_25,
  input          io_cin_26,
  input          io_cin_27,
  input          io_cin_28,
  input          io_cin_29,
  input          io_cin_30,
  input          io_cin_31,
  input          io_cin_32,
  output [31:0]  io_cout
);
  wire  c__0 = io_in_0[0]; // @[WallaceTest.scala 105:23]
  wire  c__1 = io_in_1[0]; // @[WallaceTest.scala 105:23]
  wire  c__2 = io_in_2[0]; // @[WallaceTest.scala 105:23]
  wire  c__3 = io_in_3[0]; // @[WallaceTest.scala 105:23]
  wire  c__4 = io_in_4[0]; // @[WallaceTest.scala 105:23]
  wire  c__5 = io_in_5[0]; // @[WallaceTest.scala 105:23]
  wire  c__6 = io_in_6[0]; // @[WallaceTest.scala 105:23]
  wire  c__7 = io_in_7[0]; // @[WallaceTest.scala 105:23]
  wire  c__8 = io_in_8[0]; // @[WallaceTest.scala 105:23]
  wire  c__9 = io_in_9[0]; // @[WallaceTest.scala 105:23]
  wire  c__10 = io_in_10[0]; // @[WallaceTest.scala 105:23]
  wire  c__11 = io_in_11[0]; // @[WallaceTest.scala 105:23]
  wire  c__12 = io_in_12[0]; // @[WallaceTest.scala 105:23]
  wire  c__13 = io_in_13[0]; // @[WallaceTest.scala 105:23]
  wire  c__14 = io_in_14[0]; // @[WallaceTest.scala 105:23]
  wire  c__15 = io_in_15[0]; // @[WallaceTest.scala 105:23]
  wire  c__16 = io_in_16[0]; // @[WallaceTest.scala 105:23]
  wire  c__17 = io_in_17[0]; // @[WallaceTest.scala 105:23]
  wire  c__18 = io_in_18[0]; // @[WallaceTest.scala 105:23]
  wire  c__19 = io_in_19[0]; // @[WallaceTest.scala 105:23]
  wire  c__20 = io_in_20[0]; // @[WallaceTest.scala 105:23]
  wire  c__21 = io_in_21[0]; // @[WallaceTest.scala 105:23]
  wire  c__22 = io_in_22[0]; // @[WallaceTest.scala 105:23]
  wire  c__23 = io_in_23[0]; // @[WallaceTest.scala 105:23]
  wire  c__24 = io_in_24[0]; // @[WallaceTest.scala 105:23]
  wire  c__25 = io_in_25[0]; // @[WallaceTest.scala 105:23]
  wire  c__26 = io_in_26[0]; // @[WallaceTest.scala 105:23]
  wire  c__27 = io_in_27[0]; // @[WallaceTest.scala 105:23]
  wire  c__28 = io_in_28[0]; // @[WallaceTest.scala 105:23]
  wire  c__29 = io_in_29[0]; // @[WallaceTest.scala 105:23]
  wire  c__30 = io_in_30[0]; // @[WallaceTest.scala 105:23]
  wire  c__31 = io_in_31[0]; // @[WallaceTest.scala 105:23]
  wire  c__32 = io_in_32[0]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_0_lo_lo = {c__7,c__6,c__5,c__4,c__3,c__2,c__1,c__0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_0_lo = {c__15,c__14,c__13,c__12,c__11,c__10,c__9,c__8,io_out_0_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_0_hi_lo = {c__23,c__22,c__21,c__20,c__19,c__18,c__17,c__16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_0_hi = {c__32,c__31,c__30,c__29,c__28,c__27,c__26,c__25,c__24,io_out_0_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_1_0 = io_in_0[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_1 = io_in_1[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_2 = io_in_2[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_3 = io_in_3[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_4 = io_in_4[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_5 = io_in_5[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_6 = io_in_6[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_7 = io_in_7[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_8 = io_in_8[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_9 = io_in_9[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_10 = io_in_10[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_11 = io_in_11[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_12 = io_in_12[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_13 = io_in_13[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_14 = io_in_14[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_15 = io_in_15[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_16 = io_in_16[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_17 = io_in_17[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_18 = io_in_18[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_19 = io_in_19[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_20 = io_in_20[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_21 = io_in_21[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_22 = io_in_22[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_23 = io_in_23[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_24 = io_in_24[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_25 = io_in_25[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_26 = io_in_26[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_27 = io_in_27[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_28 = io_in_28[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_29 = io_in_29[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_30 = io_in_30[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_31 = io_in_31[1]; // @[WallaceTest.scala 105:23]
  wire  c_1_32 = io_in_32[1]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_1_lo_lo = {c_1_7,c_1_6,c_1_5,c_1_4,c_1_3,c_1_2,c_1_1,c_1_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_1_lo = {c_1_15,c_1_14,c_1_13,c_1_12,c_1_11,c_1_10,c_1_9,c_1_8,io_out_1_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_1_hi_lo = {c_1_23,c_1_22,c_1_21,c_1_20,c_1_19,c_1_18,c_1_17,c_1_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_1_hi = {c_1_32,c_1_31,c_1_30,c_1_29,c_1_28,c_1_27,c_1_26,c_1_25,c_1_24,io_out_1_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_2_0 = io_in_0[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_1 = io_in_1[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_2 = io_in_2[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_3 = io_in_3[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_4 = io_in_4[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_5 = io_in_5[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_6 = io_in_6[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_7 = io_in_7[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_8 = io_in_8[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_9 = io_in_9[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_10 = io_in_10[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_11 = io_in_11[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_12 = io_in_12[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_13 = io_in_13[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_14 = io_in_14[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_15 = io_in_15[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_16 = io_in_16[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_17 = io_in_17[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_18 = io_in_18[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_19 = io_in_19[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_20 = io_in_20[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_21 = io_in_21[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_22 = io_in_22[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_23 = io_in_23[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_24 = io_in_24[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_25 = io_in_25[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_26 = io_in_26[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_27 = io_in_27[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_28 = io_in_28[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_29 = io_in_29[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_30 = io_in_30[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_31 = io_in_31[2]; // @[WallaceTest.scala 105:23]
  wire  c_2_32 = io_in_32[2]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_2_lo_lo = {c_2_7,c_2_6,c_2_5,c_2_4,c_2_3,c_2_2,c_2_1,c_2_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_2_lo = {c_2_15,c_2_14,c_2_13,c_2_12,c_2_11,c_2_10,c_2_9,c_2_8,io_out_2_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_2_hi_lo = {c_2_23,c_2_22,c_2_21,c_2_20,c_2_19,c_2_18,c_2_17,c_2_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_2_hi = {c_2_32,c_2_31,c_2_30,c_2_29,c_2_28,c_2_27,c_2_26,c_2_25,c_2_24,io_out_2_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_3_0 = io_in_0[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_1 = io_in_1[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_2 = io_in_2[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_3 = io_in_3[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_4 = io_in_4[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_5 = io_in_5[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_6 = io_in_6[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_7 = io_in_7[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_8 = io_in_8[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_9 = io_in_9[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_10 = io_in_10[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_11 = io_in_11[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_12 = io_in_12[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_13 = io_in_13[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_14 = io_in_14[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_15 = io_in_15[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_16 = io_in_16[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_17 = io_in_17[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_18 = io_in_18[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_19 = io_in_19[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_20 = io_in_20[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_21 = io_in_21[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_22 = io_in_22[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_23 = io_in_23[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_24 = io_in_24[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_25 = io_in_25[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_26 = io_in_26[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_27 = io_in_27[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_28 = io_in_28[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_29 = io_in_29[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_30 = io_in_30[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_31 = io_in_31[3]; // @[WallaceTest.scala 105:23]
  wire  c_3_32 = io_in_32[3]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_3_lo_lo = {c_3_7,c_3_6,c_3_5,c_3_4,c_3_3,c_3_2,c_3_1,c_3_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_3_lo = {c_3_15,c_3_14,c_3_13,c_3_12,c_3_11,c_3_10,c_3_9,c_3_8,io_out_3_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_3_hi_lo = {c_3_23,c_3_22,c_3_21,c_3_20,c_3_19,c_3_18,c_3_17,c_3_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_3_hi = {c_3_32,c_3_31,c_3_30,c_3_29,c_3_28,c_3_27,c_3_26,c_3_25,c_3_24,io_out_3_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_4_0 = io_in_0[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_1 = io_in_1[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_2 = io_in_2[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_3 = io_in_3[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_4 = io_in_4[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_5 = io_in_5[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_6 = io_in_6[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_7 = io_in_7[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_8 = io_in_8[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_9 = io_in_9[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_10 = io_in_10[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_11 = io_in_11[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_12 = io_in_12[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_13 = io_in_13[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_14 = io_in_14[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_15 = io_in_15[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_16 = io_in_16[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_17 = io_in_17[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_18 = io_in_18[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_19 = io_in_19[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_20 = io_in_20[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_21 = io_in_21[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_22 = io_in_22[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_23 = io_in_23[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_24 = io_in_24[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_25 = io_in_25[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_26 = io_in_26[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_27 = io_in_27[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_28 = io_in_28[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_29 = io_in_29[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_30 = io_in_30[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_31 = io_in_31[4]; // @[WallaceTest.scala 105:23]
  wire  c_4_32 = io_in_32[4]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_4_lo_lo = {c_4_7,c_4_6,c_4_5,c_4_4,c_4_3,c_4_2,c_4_1,c_4_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_4_lo = {c_4_15,c_4_14,c_4_13,c_4_12,c_4_11,c_4_10,c_4_9,c_4_8,io_out_4_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_4_hi_lo = {c_4_23,c_4_22,c_4_21,c_4_20,c_4_19,c_4_18,c_4_17,c_4_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_4_hi = {c_4_32,c_4_31,c_4_30,c_4_29,c_4_28,c_4_27,c_4_26,c_4_25,c_4_24,io_out_4_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_5_0 = io_in_0[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_1 = io_in_1[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_2 = io_in_2[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_3 = io_in_3[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_4 = io_in_4[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_5 = io_in_5[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_6 = io_in_6[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_7 = io_in_7[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_8 = io_in_8[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_9 = io_in_9[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_10 = io_in_10[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_11 = io_in_11[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_12 = io_in_12[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_13 = io_in_13[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_14 = io_in_14[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_15 = io_in_15[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_16 = io_in_16[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_17 = io_in_17[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_18 = io_in_18[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_19 = io_in_19[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_20 = io_in_20[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_21 = io_in_21[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_22 = io_in_22[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_23 = io_in_23[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_24 = io_in_24[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_25 = io_in_25[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_26 = io_in_26[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_27 = io_in_27[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_28 = io_in_28[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_29 = io_in_29[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_30 = io_in_30[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_31 = io_in_31[5]; // @[WallaceTest.scala 105:23]
  wire  c_5_32 = io_in_32[5]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_5_lo_lo = {c_5_7,c_5_6,c_5_5,c_5_4,c_5_3,c_5_2,c_5_1,c_5_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_5_lo = {c_5_15,c_5_14,c_5_13,c_5_12,c_5_11,c_5_10,c_5_9,c_5_8,io_out_5_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_5_hi_lo = {c_5_23,c_5_22,c_5_21,c_5_20,c_5_19,c_5_18,c_5_17,c_5_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_5_hi = {c_5_32,c_5_31,c_5_30,c_5_29,c_5_28,c_5_27,c_5_26,c_5_25,c_5_24,io_out_5_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_6_0 = io_in_0[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_1 = io_in_1[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_2 = io_in_2[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_3 = io_in_3[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_4 = io_in_4[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_5 = io_in_5[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_6 = io_in_6[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_7 = io_in_7[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_8 = io_in_8[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_9 = io_in_9[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_10 = io_in_10[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_11 = io_in_11[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_12 = io_in_12[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_13 = io_in_13[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_14 = io_in_14[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_15 = io_in_15[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_16 = io_in_16[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_17 = io_in_17[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_18 = io_in_18[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_19 = io_in_19[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_20 = io_in_20[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_21 = io_in_21[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_22 = io_in_22[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_23 = io_in_23[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_24 = io_in_24[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_25 = io_in_25[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_26 = io_in_26[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_27 = io_in_27[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_28 = io_in_28[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_29 = io_in_29[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_30 = io_in_30[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_31 = io_in_31[6]; // @[WallaceTest.scala 105:23]
  wire  c_6_32 = io_in_32[6]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_6_lo_lo = {c_6_7,c_6_6,c_6_5,c_6_4,c_6_3,c_6_2,c_6_1,c_6_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_6_lo = {c_6_15,c_6_14,c_6_13,c_6_12,c_6_11,c_6_10,c_6_9,c_6_8,io_out_6_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_6_hi_lo = {c_6_23,c_6_22,c_6_21,c_6_20,c_6_19,c_6_18,c_6_17,c_6_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_6_hi = {c_6_32,c_6_31,c_6_30,c_6_29,c_6_28,c_6_27,c_6_26,c_6_25,c_6_24,io_out_6_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_7_0 = io_in_0[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_1 = io_in_1[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_2 = io_in_2[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_3 = io_in_3[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_4 = io_in_4[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_5 = io_in_5[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_6 = io_in_6[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_7 = io_in_7[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_8 = io_in_8[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_9 = io_in_9[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_10 = io_in_10[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_11 = io_in_11[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_12 = io_in_12[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_13 = io_in_13[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_14 = io_in_14[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_15 = io_in_15[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_16 = io_in_16[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_17 = io_in_17[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_18 = io_in_18[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_19 = io_in_19[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_20 = io_in_20[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_21 = io_in_21[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_22 = io_in_22[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_23 = io_in_23[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_24 = io_in_24[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_25 = io_in_25[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_26 = io_in_26[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_27 = io_in_27[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_28 = io_in_28[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_29 = io_in_29[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_30 = io_in_30[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_31 = io_in_31[7]; // @[WallaceTest.scala 105:23]
  wire  c_7_32 = io_in_32[7]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_7_lo_lo = {c_7_7,c_7_6,c_7_5,c_7_4,c_7_3,c_7_2,c_7_1,c_7_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_7_lo = {c_7_15,c_7_14,c_7_13,c_7_12,c_7_11,c_7_10,c_7_9,c_7_8,io_out_7_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_7_hi_lo = {c_7_23,c_7_22,c_7_21,c_7_20,c_7_19,c_7_18,c_7_17,c_7_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_7_hi = {c_7_32,c_7_31,c_7_30,c_7_29,c_7_28,c_7_27,c_7_26,c_7_25,c_7_24,io_out_7_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_8_0 = io_in_0[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_1 = io_in_1[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_2 = io_in_2[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_3 = io_in_3[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_4 = io_in_4[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_5 = io_in_5[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_6 = io_in_6[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_7 = io_in_7[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_8 = io_in_8[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_9 = io_in_9[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_10 = io_in_10[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_11 = io_in_11[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_12 = io_in_12[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_13 = io_in_13[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_14 = io_in_14[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_15 = io_in_15[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_16 = io_in_16[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_17 = io_in_17[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_18 = io_in_18[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_19 = io_in_19[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_20 = io_in_20[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_21 = io_in_21[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_22 = io_in_22[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_23 = io_in_23[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_24 = io_in_24[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_25 = io_in_25[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_26 = io_in_26[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_27 = io_in_27[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_28 = io_in_28[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_29 = io_in_29[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_30 = io_in_30[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_31 = io_in_31[8]; // @[WallaceTest.scala 105:23]
  wire  c_8_32 = io_in_32[8]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_8_lo_lo = {c_8_7,c_8_6,c_8_5,c_8_4,c_8_3,c_8_2,c_8_1,c_8_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_8_lo = {c_8_15,c_8_14,c_8_13,c_8_12,c_8_11,c_8_10,c_8_9,c_8_8,io_out_8_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_8_hi_lo = {c_8_23,c_8_22,c_8_21,c_8_20,c_8_19,c_8_18,c_8_17,c_8_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_8_hi = {c_8_32,c_8_31,c_8_30,c_8_29,c_8_28,c_8_27,c_8_26,c_8_25,c_8_24,io_out_8_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_9_0 = io_in_0[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_1 = io_in_1[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_2 = io_in_2[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_3 = io_in_3[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_4 = io_in_4[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_5 = io_in_5[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_6 = io_in_6[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_7 = io_in_7[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_8 = io_in_8[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_9 = io_in_9[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_10 = io_in_10[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_11 = io_in_11[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_12 = io_in_12[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_13 = io_in_13[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_14 = io_in_14[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_15 = io_in_15[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_16 = io_in_16[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_17 = io_in_17[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_18 = io_in_18[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_19 = io_in_19[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_20 = io_in_20[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_21 = io_in_21[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_22 = io_in_22[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_23 = io_in_23[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_24 = io_in_24[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_25 = io_in_25[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_26 = io_in_26[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_27 = io_in_27[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_28 = io_in_28[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_29 = io_in_29[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_30 = io_in_30[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_31 = io_in_31[9]; // @[WallaceTest.scala 105:23]
  wire  c_9_32 = io_in_32[9]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_9_lo_lo = {c_9_7,c_9_6,c_9_5,c_9_4,c_9_3,c_9_2,c_9_1,c_9_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_9_lo = {c_9_15,c_9_14,c_9_13,c_9_12,c_9_11,c_9_10,c_9_9,c_9_8,io_out_9_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_9_hi_lo = {c_9_23,c_9_22,c_9_21,c_9_20,c_9_19,c_9_18,c_9_17,c_9_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_9_hi = {c_9_32,c_9_31,c_9_30,c_9_29,c_9_28,c_9_27,c_9_26,c_9_25,c_9_24,io_out_9_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_10_0 = io_in_0[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_1 = io_in_1[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_2 = io_in_2[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_3 = io_in_3[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_4 = io_in_4[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_5 = io_in_5[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_6 = io_in_6[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_7 = io_in_7[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_8 = io_in_8[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_9 = io_in_9[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_10 = io_in_10[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_11 = io_in_11[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_12 = io_in_12[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_13 = io_in_13[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_14 = io_in_14[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_15 = io_in_15[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_16 = io_in_16[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_17 = io_in_17[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_18 = io_in_18[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_19 = io_in_19[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_20 = io_in_20[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_21 = io_in_21[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_22 = io_in_22[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_23 = io_in_23[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_24 = io_in_24[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_25 = io_in_25[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_26 = io_in_26[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_27 = io_in_27[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_28 = io_in_28[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_29 = io_in_29[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_30 = io_in_30[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_31 = io_in_31[10]; // @[WallaceTest.scala 105:23]
  wire  c_10_32 = io_in_32[10]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_10_lo_lo = {c_10_7,c_10_6,c_10_5,c_10_4,c_10_3,c_10_2,c_10_1,c_10_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_10_lo = {c_10_15,c_10_14,c_10_13,c_10_12,c_10_11,c_10_10,c_10_9,c_10_8,io_out_10_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_10_hi_lo = {c_10_23,c_10_22,c_10_21,c_10_20,c_10_19,c_10_18,c_10_17,c_10_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_10_hi = {c_10_32,c_10_31,c_10_30,c_10_29,c_10_28,c_10_27,c_10_26,c_10_25,c_10_24,io_out_10_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_11_0 = io_in_0[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_1 = io_in_1[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_2 = io_in_2[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_3 = io_in_3[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_4 = io_in_4[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_5 = io_in_5[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_6 = io_in_6[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_7 = io_in_7[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_8 = io_in_8[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_9 = io_in_9[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_10 = io_in_10[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_11 = io_in_11[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_12 = io_in_12[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_13 = io_in_13[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_14 = io_in_14[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_15 = io_in_15[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_16 = io_in_16[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_17 = io_in_17[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_18 = io_in_18[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_19 = io_in_19[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_20 = io_in_20[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_21 = io_in_21[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_22 = io_in_22[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_23 = io_in_23[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_24 = io_in_24[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_25 = io_in_25[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_26 = io_in_26[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_27 = io_in_27[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_28 = io_in_28[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_29 = io_in_29[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_30 = io_in_30[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_31 = io_in_31[11]; // @[WallaceTest.scala 105:23]
  wire  c_11_32 = io_in_32[11]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_11_lo_lo = {c_11_7,c_11_6,c_11_5,c_11_4,c_11_3,c_11_2,c_11_1,c_11_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_11_lo = {c_11_15,c_11_14,c_11_13,c_11_12,c_11_11,c_11_10,c_11_9,c_11_8,io_out_11_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_11_hi_lo = {c_11_23,c_11_22,c_11_21,c_11_20,c_11_19,c_11_18,c_11_17,c_11_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_11_hi = {c_11_32,c_11_31,c_11_30,c_11_29,c_11_28,c_11_27,c_11_26,c_11_25,c_11_24,io_out_11_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_12_0 = io_in_0[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_1 = io_in_1[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_2 = io_in_2[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_3 = io_in_3[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_4 = io_in_4[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_5 = io_in_5[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_6 = io_in_6[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_7 = io_in_7[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_8 = io_in_8[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_9 = io_in_9[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_10 = io_in_10[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_11 = io_in_11[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_12 = io_in_12[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_13 = io_in_13[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_14 = io_in_14[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_15 = io_in_15[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_16 = io_in_16[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_17 = io_in_17[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_18 = io_in_18[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_19 = io_in_19[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_20 = io_in_20[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_21 = io_in_21[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_22 = io_in_22[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_23 = io_in_23[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_24 = io_in_24[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_25 = io_in_25[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_26 = io_in_26[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_27 = io_in_27[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_28 = io_in_28[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_29 = io_in_29[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_30 = io_in_30[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_31 = io_in_31[12]; // @[WallaceTest.scala 105:23]
  wire  c_12_32 = io_in_32[12]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_12_lo_lo = {c_12_7,c_12_6,c_12_5,c_12_4,c_12_3,c_12_2,c_12_1,c_12_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_12_lo = {c_12_15,c_12_14,c_12_13,c_12_12,c_12_11,c_12_10,c_12_9,c_12_8,io_out_12_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_12_hi_lo = {c_12_23,c_12_22,c_12_21,c_12_20,c_12_19,c_12_18,c_12_17,c_12_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_12_hi = {c_12_32,c_12_31,c_12_30,c_12_29,c_12_28,c_12_27,c_12_26,c_12_25,c_12_24,io_out_12_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_13_0 = io_in_0[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_1 = io_in_1[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_2 = io_in_2[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_3 = io_in_3[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_4 = io_in_4[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_5 = io_in_5[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_6 = io_in_6[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_7 = io_in_7[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_8 = io_in_8[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_9 = io_in_9[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_10 = io_in_10[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_11 = io_in_11[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_12 = io_in_12[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_13 = io_in_13[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_14 = io_in_14[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_15 = io_in_15[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_16 = io_in_16[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_17 = io_in_17[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_18 = io_in_18[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_19 = io_in_19[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_20 = io_in_20[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_21 = io_in_21[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_22 = io_in_22[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_23 = io_in_23[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_24 = io_in_24[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_25 = io_in_25[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_26 = io_in_26[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_27 = io_in_27[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_28 = io_in_28[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_29 = io_in_29[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_30 = io_in_30[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_31 = io_in_31[13]; // @[WallaceTest.scala 105:23]
  wire  c_13_32 = io_in_32[13]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_13_lo_lo = {c_13_7,c_13_6,c_13_5,c_13_4,c_13_3,c_13_2,c_13_1,c_13_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_13_lo = {c_13_15,c_13_14,c_13_13,c_13_12,c_13_11,c_13_10,c_13_9,c_13_8,io_out_13_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_13_hi_lo = {c_13_23,c_13_22,c_13_21,c_13_20,c_13_19,c_13_18,c_13_17,c_13_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_13_hi = {c_13_32,c_13_31,c_13_30,c_13_29,c_13_28,c_13_27,c_13_26,c_13_25,c_13_24,io_out_13_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_14_0 = io_in_0[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_1 = io_in_1[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_2 = io_in_2[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_3 = io_in_3[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_4 = io_in_4[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_5 = io_in_5[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_6 = io_in_6[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_7 = io_in_7[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_8 = io_in_8[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_9 = io_in_9[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_10 = io_in_10[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_11 = io_in_11[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_12 = io_in_12[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_13 = io_in_13[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_14 = io_in_14[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_15 = io_in_15[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_16 = io_in_16[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_17 = io_in_17[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_18 = io_in_18[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_19 = io_in_19[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_20 = io_in_20[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_21 = io_in_21[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_22 = io_in_22[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_23 = io_in_23[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_24 = io_in_24[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_25 = io_in_25[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_26 = io_in_26[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_27 = io_in_27[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_28 = io_in_28[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_29 = io_in_29[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_30 = io_in_30[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_31 = io_in_31[14]; // @[WallaceTest.scala 105:23]
  wire  c_14_32 = io_in_32[14]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_14_lo_lo = {c_14_7,c_14_6,c_14_5,c_14_4,c_14_3,c_14_2,c_14_1,c_14_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_14_lo = {c_14_15,c_14_14,c_14_13,c_14_12,c_14_11,c_14_10,c_14_9,c_14_8,io_out_14_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_14_hi_lo = {c_14_23,c_14_22,c_14_21,c_14_20,c_14_19,c_14_18,c_14_17,c_14_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_14_hi = {c_14_32,c_14_31,c_14_30,c_14_29,c_14_28,c_14_27,c_14_26,c_14_25,c_14_24,io_out_14_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_15_0 = io_in_0[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_1 = io_in_1[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_2 = io_in_2[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_3 = io_in_3[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_4 = io_in_4[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_5 = io_in_5[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_6 = io_in_6[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_7 = io_in_7[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_8 = io_in_8[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_9 = io_in_9[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_10 = io_in_10[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_11 = io_in_11[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_12 = io_in_12[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_13 = io_in_13[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_14 = io_in_14[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_15 = io_in_15[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_16 = io_in_16[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_17 = io_in_17[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_18 = io_in_18[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_19 = io_in_19[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_20 = io_in_20[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_21 = io_in_21[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_22 = io_in_22[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_23 = io_in_23[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_24 = io_in_24[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_25 = io_in_25[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_26 = io_in_26[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_27 = io_in_27[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_28 = io_in_28[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_29 = io_in_29[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_30 = io_in_30[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_31 = io_in_31[15]; // @[WallaceTest.scala 105:23]
  wire  c_15_32 = io_in_32[15]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_15_lo_lo = {c_15_7,c_15_6,c_15_5,c_15_4,c_15_3,c_15_2,c_15_1,c_15_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_15_lo = {c_15_15,c_15_14,c_15_13,c_15_12,c_15_11,c_15_10,c_15_9,c_15_8,io_out_15_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_15_hi_lo = {c_15_23,c_15_22,c_15_21,c_15_20,c_15_19,c_15_18,c_15_17,c_15_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_15_hi = {c_15_32,c_15_31,c_15_30,c_15_29,c_15_28,c_15_27,c_15_26,c_15_25,c_15_24,io_out_15_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_16_0 = io_in_0[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_1 = io_in_1[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_2 = io_in_2[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_3 = io_in_3[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_4 = io_in_4[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_5 = io_in_5[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_6 = io_in_6[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_7 = io_in_7[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_8 = io_in_8[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_9 = io_in_9[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_10 = io_in_10[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_11 = io_in_11[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_12 = io_in_12[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_13 = io_in_13[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_14 = io_in_14[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_15 = io_in_15[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_16 = io_in_16[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_17 = io_in_17[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_18 = io_in_18[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_19 = io_in_19[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_20 = io_in_20[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_21 = io_in_21[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_22 = io_in_22[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_23 = io_in_23[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_24 = io_in_24[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_25 = io_in_25[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_26 = io_in_26[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_27 = io_in_27[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_28 = io_in_28[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_29 = io_in_29[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_30 = io_in_30[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_31 = io_in_31[16]; // @[WallaceTest.scala 105:23]
  wire  c_16_32 = io_in_32[16]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_16_lo_lo = {c_16_7,c_16_6,c_16_5,c_16_4,c_16_3,c_16_2,c_16_1,c_16_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_16_lo = {c_16_15,c_16_14,c_16_13,c_16_12,c_16_11,c_16_10,c_16_9,c_16_8,io_out_16_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_16_hi_lo = {c_16_23,c_16_22,c_16_21,c_16_20,c_16_19,c_16_18,c_16_17,c_16_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_16_hi = {c_16_32,c_16_31,c_16_30,c_16_29,c_16_28,c_16_27,c_16_26,c_16_25,c_16_24,io_out_16_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_17_0 = io_in_0[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_1 = io_in_1[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_2 = io_in_2[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_3 = io_in_3[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_4 = io_in_4[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_5 = io_in_5[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_6 = io_in_6[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_7 = io_in_7[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_8 = io_in_8[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_9 = io_in_9[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_10 = io_in_10[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_11 = io_in_11[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_12 = io_in_12[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_13 = io_in_13[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_14 = io_in_14[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_15 = io_in_15[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_16 = io_in_16[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_17 = io_in_17[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_18 = io_in_18[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_19 = io_in_19[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_20 = io_in_20[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_21 = io_in_21[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_22 = io_in_22[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_23 = io_in_23[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_24 = io_in_24[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_25 = io_in_25[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_26 = io_in_26[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_27 = io_in_27[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_28 = io_in_28[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_29 = io_in_29[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_30 = io_in_30[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_31 = io_in_31[17]; // @[WallaceTest.scala 105:23]
  wire  c_17_32 = io_in_32[17]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_17_lo_lo = {c_17_7,c_17_6,c_17_5,c_17_4,c_17_3,c_17_2,c_17_1,c_17_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_17_lo = {c_17_15,c_17_14,c_17_13,c_17_12,c_17_11,c_17_10,c_17_9,c_17_8,io_out_17_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_17_hi_lo = {c_17_23,c_17_22,c_17_21,c_17_20,c_17_19,c_17_18,c_17_17,c_17_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_17_hi = {c_17_32,c_17_31,c_17_30,c_17_29,c_17_28,c_17_27,c_17_26,c_17_25,c_17_24,io_out_17_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_18_0 = io_in_0[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_1 = io_in_1[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_2 = io_in_2[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_3 = io_in_3[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_4 = io_in_4[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_5 = io_in_5[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_6 = io_in_6[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_7 = io_in_7[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_8 = io_in_8[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_9 = io_in_9[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_10 = io_in_10[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_11 = io_in_11[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_12 = io_in_12[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_13 = io_in_13[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_14 = io_in_14[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_15 = io_in_15[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_16 = io_in_16[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_17 = io_in_17[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_18 = io_in_18[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_19 = io_in_19[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_20 = io_in_20[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_21 = io_in_21[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_22 = io_in_22[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_23 = io_in_23[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_24 = io_in_24[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_25 = io_in_25[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_26 = io_in_26[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_27 = io_in_27[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_28 = io_in_28[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_29 = io_in_29[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_30 = io_in_30[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_31 = io_in_31[18]; // @[WallaceTest.scala 105:23]
  wire  c_18_32 = io_in_32[18]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_18_lo_lo = {c_18_7,c_18_6,c_18_5,c_18_4,c_18_3,c_18_2,c_18_1,c_18_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_18_lo = {c_18_15,c_18_14,c_18_13,c_18_12,c_18_11,c_18_10,c_18_9,c_18_8,io_out_18_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_18_hi_lo = {c_18_23,c_18_22,c_18_21,c_18_20,c_18_19,c_18_18,c_18_17,c_18_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_18_hi = {c_18_32,c_18_31,c_18_30,c_18_29,c_18_28,c_18_27,c_18_26,c_18_25,c_18_24,io_out_18_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_19_0 = io_in_0[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_1 = io_in_1[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_2 = io_in_2[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_3 = io_in_3[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_4 = io_in_4[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_5 = io_in_5[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_6 = io_in_6[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_7 = io_in_7[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_8 = io_in_8[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_9 = io_in_9[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_10 = io_in_10[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_11 = io_in_11[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_12 = io_in_12[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_13 = io_in_13[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_14 = io_in_14[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_15 = io_in_15[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_16 = io_in_16[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_17 = io_in_17[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_18 = io_in_18[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_19 = io_in_19[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_20 = io_in_20[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_21 = io_in_21[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_22 = io_in_22[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_23 = io_in_23[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_24 = io_in_24[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_25 = io_in_25[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_26 = io_in_26[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_27 = io_in_27[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_28 = io_in_28[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_29 = io_in_29[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_30 = io_in_30[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_31 = io_in_31[19]; // @[WallaceTest.scala 105:23]
  wire  c_19_32 = io_in_32[19]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_19_lo_lo = {c_19_7,c_19_6,c_19_5,c_19_4,c_19_3,c_19_2,c_19_1,c_19_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_19_lo = {c_19_15,c_19_14,c_19_13,c_19_12,c_19_11,c_19_10,c_19_9,c_19_8,io_out_19_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_19_hi_lo = {c_19_23,c_19_22,c_19_21,c_19_20,c_19_19,c_19_18,c_19_17,c_19_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_19_hi = {c_19_32,c_19_31,c_19_30,c_19_29,c_19_28,c_19_27,c_19_26,c_19_25,c_19_24,io_out_19_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_20_0 = io_in_0[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_1 = io_in_1[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_2 = io_in_2[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_3 = io_in_3[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_4 = io_in_4[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_5 = io_in_5[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_6 = io_in_6[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_7 = io_in_7[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_8 = io_in_8[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_9 = io_in_9[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_10 = io_in_10[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_11 = io_in_11[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_12 = io_in_12[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_13 = io_in_13[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_14 = io_in_14[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_15 = io_in_15[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_16 = io_in_16[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_17 = io_in_17[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_18 = io_in_18[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_19 = io_in_19[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_20 = io_in_20[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_21 = io_in_21[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_22 = io_in_22[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_23 = io_in_23[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_24 = io_in_24[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_25 = io_in_25[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_26 = io_in_26[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_27 = io_in_27[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_28 = io_in_28[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_29 = io_in_29[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_30 = io_in_30[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_31 = io_in_31[20]; // @[WallaceTest.scala 105:23]
  wire  c_20_32 = io_in_32[20]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_20_lo_lo = {c_20_7,c_20_6,c_20_5,c_20_4,c_20_3,c_20_2,c_20_1,c_20_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_20_lo = {c_20_15,c_20_14,c_20_13,c_20_12,c_20_11,c_20_10,c_20_9,c_20_8,io_out_20_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_20_hi_lo = {c_20_23,c_20_22,c_20_21,c_20_20,c_20_19,c_20_18,c_20_17,c_20_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_20_hi = {c_20_32,c_20_31,c_20_30,c_20_29,c_20_28,c_20_27,c_20_26,c_20_25,c_20_24,io_out_20_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_21_0 = io_in_0[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_1 = io_in_1[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_2 = io_in_2[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_3 = io_in_3[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_4 = io_in_4[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_5 = io_in_5[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_6 = io_in_6[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_7 = io_in_7[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_8 = io_in_8[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_9 = io_in_9[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_10 = io_in_10[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_11 = io_in_11[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_12 = io_in_12[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_13 = io_in_13[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_14 = io_in_14[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_15 = io_in_15[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_16 = io_in_16[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_17 = io_in_17[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_18 = io_in_18[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_19 = io_in_19[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_20 = io_in_20[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_21 = io_in_21[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_22 = io_in_22[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_23 = io_in_23[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_24 = io_in_24[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_25 = io_in_25[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_26 = io_in_26[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_27 = io_in_27[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_28 = io_in_28[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_29 = io_in_29[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_30 = io_in_30[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_31 = io_in_31[21]; // @[WallaceTest.scala 105:23]
  wire  c_21_32 = io_in_32[21]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_21_lo_lo = {c_21_7,c_21_6,c_21_5,c_21_4,c_21_3,c_21_2,c_21_1,c_21_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_21_lo = {c_21_15,c_21_14,c_21_13,c_21_12,c_21_11,c_21_10,c_21_9,c_21_8,io_out_21_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_21_hi_lo = {c_21_23,c_21_22,c_21_21,c_21_20,c_21_19,c_21_18,c_21_17,c_21_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_21_hi = {c_21_32,c_21_31,c_21_30,c_21_29,c_21_28,c_21_27,c_21_26,c_21_25,c_21_24,io_out_21_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_22_0 = io_in_0[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_1 = io_in_1[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_2 = io_in_2[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_3 = io_in_3[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_4 = io_in_4[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_5 = io_in_5[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_6 = io_in_6[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_7 = io_in_7[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_8 = io_in_8[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_9 = io_in_9[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_10 = io_in_10[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_11 = io_in_11[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_12 = io_in_12[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_13 = io_in_13[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_14 = io_in_14[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_15 = io_in_15[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_16 = io_in_16[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_17 = io_in_17[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_18 = io_in_18[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_19 = io_in_19[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_20 = io_in_20[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_21 = io_in_21[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_22 = io_in_22[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_23 = io_in_23[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_24 = io_in_24[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_25 = io_in_25[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_26 = io_in_26[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_27 = io_in_27[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_28 = io_in_28[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_29 = io_in_29[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_30 = io_in_30[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_31 = io_in_31[22]; // @[WallaceTest.scala 105:23]
  wire  c_22_32 = io_in_32[22]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_22_lo_lo = {c_22_7,c_22_6,c_22_5,c_22_4,c_22_3,c_22_2,c_22_1,c_22_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_22_lo = {c_22_15,c_22_14,c_22_13,c_22_12,c_22_11,c_22_10,c_22_9,c_22_8,io_out_22_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_22_hi_lo = {c_22_23,c_22_22,c_22_21,c_22_20,c_22_19,c_22_18,c_22_17,c_22_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_22_hi = {c_22_32,c_22_31,c_22_30,c_22_29,c_22_28,c_22_27,c_22_26,c_22_25,c_22_24,io_out_22_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_23_0 = io_in_0[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_1 = io_in_1[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_2 = io_in_2[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_3 = io_in_3[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_4 = io_in_4[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_5 = io_in_5[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_6 = io_in_6[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_7 = io_in_7[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_8 = io_in_8[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_9 = io_in_9[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_10 = io_in_10[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_11 = io_in_11[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_12 = io_in_12[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_13 = io_in_13[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_14 = io_in_14[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_15 = io_in_15[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_16 = io_in_16[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_17 = io_in_17[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_18 = io_in_18[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_19 = io_in_19[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_20 = io_in_20[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_21 = io_in_21[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_22 = io_in_22[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_23 = io_in_23[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_24 = io_in_24[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_25 = io_in_25[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_26 = io_in_26[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_27 = io_in_27[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_28 = io_in_28[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_29 = io_in_29[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_30 = io_in_30[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_31 = io_in_31[23]; // @[WallaceTest.scala 105:23]
  wire  c_23_32 = io_in_32[23]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_23_lo_lo = {c_23_7,c_23_6,c_23_5,c_23_4,c_23_3,c_23_2,c_23_1,c_23_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_23_lo = {c_23_15,c_23_14,c_23_13,c_23_12,c_23_11,c_23_10,c_23_9,c_23_8,io_out_23_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_23_hi_lo = {c_23_23,c_23_22,c_23_21,c_23_20,c_23_19,c_23_18,c_23_17,c_23_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_23_hi = {c_23_32,c_23_31,c_23_30,c_23_29,c_23_28,c_23_27,c_23_26,c_23_25,c_23_24,io_out_23_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_24_0 = io_in_0[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_1 = io_in_1[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_2 = io_in_2[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_3 = io_in_3[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_4 = io_in_4[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_5 = io_in_5[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_6 = io_in_6[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_7 = io_in_7[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_8 = io_in_8[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_9 = io_in_9[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_10 = io_in_10[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_11 = io_in_11[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_12 = io_in_12[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_13 = io_in_13[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_14 = io_in_14[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_15 = io_in_15[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_16 = io_in_16[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_17 = io_in_17[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_18 = io_in_18[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_19 = io_in_19[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_20 = io_in_20[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_21 = io_in_21[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_22 = io_in_22[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_23 = io_in_23[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_24 = io_in_24[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_25 = io_in_25[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_26 = io_in_26[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_27 = io_in_27[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_28 = io_in_28[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_29 = io_in_29[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_30 = io_in_30[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_31 = io_in_31[24]; // @[WallaceTest.scala 105:23]
  wire  c_24_32 = io_in_32[24]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_24_lo_lo = {c_24_7,c_24_6,c_24_5,c_24_4,c_24_3,c_24_2,c_24_1,c_24_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_24_lo = {c_24_15,c_24_14,c_24_13,c_24_12,c_24_11,c_24_10,c_24_9,c_24_8,io_out_24_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_24_hi_lo = {c_24_23,c_24_22,c_24_21,c_24_20,c_24_19,c_24_18,c_24_17,c_24_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_24_hi = {c_24_32,c_24_31,c_24_30,c_24_29,c_24_28,c_24_27,c_24_26,c_24_25,c_24_24,io_out_24_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_25_0 = io_in_0[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_1 = io_in_1[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_2 = io_in_2[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_3 = io_in_3[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_4 = io_in_4[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_5 = io_in_5[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_6 = io_in_6[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_7 = io_in_7[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_8 = io_in_8[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_9 = io_in_9[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_10 = io_in_10[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_11 = io_in_11[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_12 = io_in_12[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_13 = io_in_13[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_14 = io_in_14[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_15 = io_in_15[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_16 = io_in_16[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_17 = io_in_17[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_18 = io_in_18[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_19 = io_in_19[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_20 = io_in_20[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_21 = io_in_21[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_22 = io_in_22[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_23 = io_in_23[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_24 = io_in_24[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_25 = io_in_25[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_26 = io_in_26[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_27 = io_in_27[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_28 = io_in_28[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_29 = io_in_29[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_30 = io_in_30[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_31 = io_in_31[25]; // @[WallaceTest.scala 105:23]
  wire  c_25_32 = io_in_32[25]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_25_lo_lo = {c_25_7,c_25_6,c_25_5,c_25_4,c_25_3,c_25_2,c_25_1,c_25_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_25_lo = {c_25_15,c_25_14,c_25_13,c_25_12,c_25_11,c_25_10,c_25_9,c_25_8,io_out_25_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_25_hi_lo = {c_25_23,c_25_22,c_25_21,c_25_20,c_25_19,c_25_18,c_25_17,c_25_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_25_hi = {c_25_32,c_25_31,c_25_30,c_25_29,c_25_28,c_25_27,c_25_26,c_25_25,c_25_24,io_out_25_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_26_0 = io_in_0[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_1 = io_in_1[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_2 = io_in_2[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_3 = io_in_3[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_4 = io_in_4[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_5 = io_in_5[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_6 = io_in_6[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_7 = io_in_7[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_8 = io_in_8[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_9 = io_in_9[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_10 = io_in_10[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_11 = io_in_11[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_12 = io_in_12[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_13 = io_in_13[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_14 = io_in_14[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_15 = io_in_15[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_16 = io_in_16[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_17 = io_in_17[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_18 = io_in_18[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_19 = io_in_19[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_20 = io_in_20[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_21 = io_in_21[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_22 = io_in_22[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_23 = io_in_23[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_24 = io_in_24[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_25 = io_in_25[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_26 = io_in_26[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_27 = io_in_27[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_28 = io_in_28[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_29 = io_in_29[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_30 = io_in_30[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_31 = io_in_31[26]; // @[WallaceTest.scala 105:23]
  wire  c_26_32 = io_in_32[26]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_26_lo_lo = {c_26_7,c_26_6,c_26_5,c_26_4,c_26_3,c_26_2,c_26_1,c_26_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_26_lo = {c_26_15,c_26_14,c_26_13,c_26_12,c_26_11,c_26_10,c_26_9,c_26_8,io_out_26_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_26_hi_lo = {c_26_23,c_26_22,c_26_21,c_26_20,c_26_19,c_26_18,c_26_17,c_26_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_26_hi = {c_26_32,c_26_31,c_26_30,c_26_29,c_26_28,c_26_27,c_26_26,c_26_25,c_26_24,io_out_26_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_27_0 = io_in_0[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_1 = io_in_1[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_2 = io_in_2[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_3 = io_in_3[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_4 = io_in_4[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_5 = io_in_5[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_6 = io_in_6[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_7 = io_in_7[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_8 = io_in_8[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_9 = io_in_9[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_10 = io_in_10[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_11 = io_in_11[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_12 = io_in_12[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_13 = io_in_13[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_14 = io_in_14[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_15 = io_in_15[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_16 = io_in_16[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_17 = io_in_17[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_18 = io_in_18[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_19 = io_in_19[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_20 = io_in_20[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_21 = io_in_21[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_22 = io_in_22[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_23 = io_in_23[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_24 = io_in_24[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_25 = io_in_25[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_26 = io_in_26[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_27 = io_in_27[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_28 = io_in_28[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_29 = io_in_29[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_30 = io_in_30[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_31 = io_in_31[27]; // @[WallaceTest.scala 105:23]
  wire  c_27_32 = io_in_32[27]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_27_lo_lo = {c_27_7,c_27_6,c_27_5,c_27_4,c_27_3,c_27_2,c_27_1,c_27_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_27_lo = {c_27_15,c_27_14,c_27_13,c_27_12,c_27_11,c_27_10,c_27_9,c_27_8,io_out_27_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_27_hi_lo = {c_27_23,c_27_22,c_27_21,c_27_20,c_27_19,c_27_18,c_27_17,c_27_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_27_hi = {c_27_32,c_27_31,c_27_30,c_27_29,c_27_28,c_27_27,c_27_26,c_27_25,c_27_24,io_out_27_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_28_0 = io_in_0[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_1 = io_in_1[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_2 = io_in_2[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_3 = io_in_3[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_4 = io_in_4[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_5 = io_in_5[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_6 = io_in_6[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_7 = io_in_7[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_8 = io_in_8[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_9 = io_in_9[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_10 = io_in_10[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_11 = io_in_11[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_12 = io_in_12[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_13 = io_in_13[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_14 = io_in_14[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_15 = io_in_15[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_16 = io_in_16[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_17 = io_in_17[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_18 = io_in_18[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_19 = io_in_19[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_20 = io_in_20[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_21 = io_in_21[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_22 = io_in_22[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_23 = io_in_23[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_24 = io_in_24[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_25 = io_in_25[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_26 = io_in_26[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_27 = io_in_27[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_28 = io_in_28[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_29 = io_in_29[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_30 = io_in_30[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_31 = io_in_31[28]; // @[WallaceTest.scala 105:23]
  wire  c_28_32 = io_in_32[28]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_28_lo_lo = {c_28_7,c_28_6,c_28_5,c_28_4,c_28_3,c_28_2,c_28_1,c_28_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_28_lo = {c_28_15,c_28_14,c_28_13,c_28_12,c_28_11,c_28_10,c_28_9,c_28_8,io_out_28_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_28_hi_lo = {c_28_23,c_28_22,c_28_21,c_28_20,c_28_19,c_28_18,c_28_17,c_28_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_28_hi = {c_28_32,c_28_31,c_28_30,c_28_29,c_28_28,c_28_27,c_28_26,c_28_25,c_28_24,io_out_28_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_29_0 = io_in_0[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_1 = io_in_1[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_2 = io_in_2[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_3 = io_in_3[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_4 = io_in_4[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_5 = io_in_5[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_6 = io_in_6[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_7 = io_in_7[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_8 = io_in_8[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_9 = io_in_9[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_10 = io_in_10[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_11 = io_in_11[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_12 = io_in_12[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_13 = io_in_13[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_14 = io_in_14[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_15 = io_in_15[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_16 = io_in_16[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_17 = io_in_17[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_18 = io_in_18[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_19 = io_in_19[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_20 = io_in_20[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_21 = io_in_21[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_22 = io_in_22[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_23 = io_in_23[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_24 = io_in_24[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_25 = io_in_25[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_26 = io_in_26[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_27 = io_in_27[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_28 = io_in_28[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_29 = io_in_29[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_30 = io_in_30[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_31 = io_in_31[29]; // @[WallaceTest.scala 105:23]
  wire  c_29_32 = io_in_32[29]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_29_lo_lo = {c_29_7,c_29_6,c_29_5,c_29_4,c_29_3,c_29_2,c_29_1,c_29_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_29_lo = {c_29_15,c_29_14,c_29_13,c_29_12,c_29_11,c_29_10,c_29_9,c_29_8,io_out_29_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_29_hi_lo = {c_29_23,c_29_22,c_29_21,c_29_20,c_29_19,c_29_18,c_29_17,c_29_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_29_hi = {c_29_32,c_29_31,c_29_30,c_29_29,c_29_28,c_29_27,c_29_26,c_29_25,c_29_24,io_out_29_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_30_0 = io_in_0[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_1 = io_in_1[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_2 = io_in_2[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_3 = io_in_3[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_4 = io_in_4[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_5 = io_in_5[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_6 = io_in_6[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_7 = io_in_7[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_8 = io_in_8[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_9 = io_in_9[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_10 = io_in_10[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_11 = io_in_11[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_12 = io_in_12[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_13 = io_in_13[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_14 = io_in_14[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_15 = io_in_15[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_16 = io_in_16[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_17 = io_in_17[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_18 = io_in_18[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_19 = io_in_19[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_20 = io_in_20[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_21 = io_in_21[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_22 = io_in_22[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_23 = io_in_23[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_24 = io_in_24[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_25 = io_in_25[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_26 = io_in_26[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_27 = io_in_27[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_28 = io_in_28[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_29 = io_in_29[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_30 = io_in_30[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_31 = io_in_31[30]; // @[WallaceTest.scala 105:23]
  wire  c_30_32 = io_in_32[30]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_30_lo_lo = {c_30_7,c_30_6,c_30_5,c_30_4,c_30_3,c_30_2,c_30_1,c_30_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_30_lo = {c_30_15,c_30_14,c_30_13,c_30_12,c_30_11,c_30_10,c_30_9,c_30_8,io_out_30_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_30_hi_lo = {c_30_23,c_30_22,c_30_21,c_30_20,c_30_19,c_30_18,c_30_17,c_30_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_30_hi = {c_30_32,c_30_31,c_30_30,c_30_29,c_30_28,c_30_27,c_30_26,c_30_25,c_30_24,io_out_30_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_31_0 = io_in_0[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_1 = io_in_1[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_2 = io_in_2[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_3 = io_in_3[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_4 = io_in_4[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_5 = io_in_5[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_6 = io_in_6[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_7 = io_in_7[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_8 = io_in_8[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_9 = io_in_9[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_10 = io_in_10[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_11 = io_in_11[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_12 = io_in_12[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_13 = io_in_13[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_14 = io_in_14[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_15 = io_in_15[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_16 = io_in_16[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_17 = io_in_17[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_18 = io_in_18[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_19 = io_in_19[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_20 = io_in_20[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_21 = io_in_21[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_22 = io_in_22[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_23 = io_in_23[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_24 = io_in_24[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_25 = io_in_25[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_26 = io_in_26[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_27 = io_in_27[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_28 = io_in_28[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_29 = io_in_29[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_30 = io_in_30[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_31 = io_in_31[31]; // @[WallaceTest.scala 105:23]
  wire  c_31_32 = io_in_32[31]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_31_lo_lo = {c_31_7,c_31_6,c_31_5,c_31_4,c_31_3,c_31_2,c_31_1,c_31_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_31_lo = {c_31_15,c_31_14,c_31_13,c_31_12,c_31_11,c_31_10,c_31_9,c_31_8,io_out_31_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_31_hi_lo = {c_31_23,c_31_22,c_31_21,c_31_20,c_31_19,c_31_18,c_31_17,c_31_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_31_hi = {c_31_32,c_31_31,c_31_30,c_31_29,c_31_28,c_31_27,c_31_26,c_31_25,c_31_24,io_out_31_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_32_0 = io_in_0[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_1 = io_in_1[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_2 = io_in_2[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_3 = io_in_3[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_4 = io_in_4[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_5 = io_in_5[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_6 = io_in_6[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_7 = io_in_7[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_8 = io_in_8[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_9 = io_in_9[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_10 = io_in_10[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_11 = io_in_11[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_12 = io_in_12[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_13 = io_in_13[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_14 = io_in_14[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_15 = io_in_15[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_16 = io_in_16[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_17 = io_in_17[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_18 = io_in_18[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_19 = io_in_19[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_20 = io_in_20[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_21 = io_in_21[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_22 = io_in_22[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_23 = io_in_23[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_24 = io_in_24[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_25 = io_in_25[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_26 = io_in_26[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_27 = io_in_27[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_28 = io_in_28[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_29 = io_in_29[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_30 = io_in_30[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_31 = io_in_31[32]; // @[WallaceTest.scala 105:23]
  wire  c_32_32 = io_in_32[32]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_32_lo_lo = {c_32_7,c_32_6,c_32_5,c_32_4,c_32_3,c_32_2,c_32_1,c_32_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_32_lo = {c_32_15,c_32_14,c_32_13,c_32_12,c_32_11,c_32_10,c_32_9,c_32_8,io_out_32_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_32_hi_lo = {c_32_23,c_32_22,c_32_21,c_32_20,c_32_19,c_32_18,c_32_17,c_32_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_32_hi = {c_32_32,c_32_31,c_32_30,c_32_29,c_32_28,c_32_27,c_32_26,c_32_25,c_32_24,io_out_32_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_33_0 = io_in_0[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_1 = io_in_1[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_2 = io_in_2[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_3 = io_in_3[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_4 = io_in_4[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_5 = io_in_5[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_6 = io_in_6[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_7 = io_in_7[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_8 = io_in_8[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_9 = io_in_9[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_10 = io_in_10[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_11 = io_in_11[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_12 = io_in_12[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_13 = io_in_13[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_14 = io_in_14[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_15 = io_in_15[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_16 = io_in_16[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_17 = io_in_17[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_18 = io_in_18[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_19 = io_in_19[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_20 = io_in_20[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_21 = io_in_21[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_22 = io_in_22[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_23 = io_in_23[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_24 = io_in_24[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_25 = io_in_25[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_26 = io_in_26[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_27 = io_in_27[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_28 = io_in_28[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_29 = io_in_29[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_30 = io_in_30[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_31 = io_in_31[33]; // @[WallaceTest.scala 105:23]
  wire  c_33_32 = io_in_32[33]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_33_lo_lo = {c_33_7,c_33_6,c_33_5,c_33_4,c_33_3,c_33_2,c_33_1,c_33_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_33_lo = {c_33_15,c_33_14,c_33_13,c_33_12,c_33_11,c_33_10,c_33_9,c_33_8,io_out_33_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_33_hi_lo = {c_33_23,c_33_22,c_33_21,c_33_20,c_33_19,c_33_18,c_33_17,c_33_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_33_hi = {c_33_32,c_33_31,c_33_30,c_33_29,c_33_28,c_33_27,c_33_26,c_33_25,c_33_24,io_out_33_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_34_0 = io_in_0[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_1 = io_in_1[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_2 = io_in_2[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_3 = io_in_3[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_4 = io_in_4[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_5 = io_in_5[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_6 = io_in_6[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_7 = io_in_7[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_8 = io_in_8[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_9 = io_in_9[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_10 = io_in_10[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_11 = io_in_11[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_12 = io_in_12[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_13 = io_in_13[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_14 = io_in_14[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_15 = io_in_15[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_16 = io_in_16[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_17 = io_in_17[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_18 = io_in_18[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_19 = io_in_19[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_20 = io_in_20[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_21 = io_in_21[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_22 = io_in_22[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_23 = io_in_23[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_24 = io_in_24[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_25 = io_in_25[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_26 = io_in_26[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_27 = io_in_27[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_28 = io_in_28[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_29 = io_in_29[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_30 = io_in_30[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_31 = io_in_31[34]; // @[WallaceTest.scala 105:23]
  wire  c_34_32 = io_in_32[34]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_34_lo_lo = {c_34_7,c_34_6,c_34_5,c_34_4,c_34_3,c_34_2,c_34_1,c_34_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_34_lo = {c_34_15,c_34_14,c_34_13,c_34_12,c_34_11,c_34_10,c_34_9,c_34_8,io_out_34_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_34_hi_lo = {c_34_23,c_34_22,c_34_21,c_34_20,c_34_19,c_34_18,c_34_17,c_34_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_34_hi = {c_34_32,c_34_31,c_34_30,c_34_29,c_34_28,c_34_27,c_34_26,c_34_25,c_34_24,io_out_34_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_35_0 = io_in_0[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_1 = io_in_1[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_2 = io_in_2[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_3 = io_in_3[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_4 = io_in_4[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_5 = io_in_5[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_6 = io_in_6[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_7 = io_in_7[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_8 = io_in_8[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_9 = io_in_9[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_10 = io_in_10[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_11 = io_in_11[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_12 = io_in_12[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_13 = io_in_13[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_14 = io_in_14[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_15 = io_in_15[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_16 = io_in_16[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_17 = io_in_17[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_18 = io_in_18[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_19 = io_in_19[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_20 = io_in_20[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_21 = io_in_21[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_22 = io_in_22[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_23 = io_in_23[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_24 = io_in_24[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_25 = io_in_25[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_26 = io_in_26[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_27 = io_in_27[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_28 = io_in_28[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_29 = io_in_29[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_30 = io_in_30[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_31 = io_in_31[35]; // @[WallaceTest.scala 105:23]
  wire  c_35_32 = io_in_32[35]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_35_lo_lo = {c_35_7,c_35_6,c_35_5,c_35_4,c_35_3,c_35_2,c_35_1,c_35_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_35_lo = {c_35_15,c_35_14,c_35_13,c_35_12,c_35_11,c_35_10,c_35_9,c_35_8,io_out_35_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_35_hi_lo = {c_35_23,c_35_22,c_35_21,c_35_20,c_35_19,c_35_18,c_35_17,c_35_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_35_hi = {c_35_32,c_35_31,c_35_30,c_35_29,c_35_28,c_35_27,c_35_26,c_35_25,c_35_24,io_out_35_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_36_0 = io_in_0[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_1 = io_in_1[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_2 = io_in_2[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_3 = io_in_3[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_4 = io_in_4[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_5 = io_in_5[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_6 = io_in_6[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_7 = io_in_7[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_8 = io_in_8[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_9 = io_in_9[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_10 = io_in_10[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_11 = io_in_11[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_12 = io_in_12[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_13 = io_in_13[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_14 = io_in_14[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_15 = io_in_15[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_16 = io_in_16[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_17 = io_in_17[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_18 = io_in_18[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_19 = io_in_19[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_20 = io_in_20[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_21 = io_in_21[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_22 = io_in_22[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_23 = io_in_23[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_24 = io_in_24[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_25 = io_in_25[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_26 = io_in_26[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_27 = io_in_27[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_28 = io_in_28[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_29 = io_in_29[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_30 = io_in_30[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_31 = io_in_31[36]; // @[WallaceTest.scala 105:23]
  wire  c_36_32 = io_in_32[36]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_36_lo_lo = {c_36_7,c_36_6,c_36_5,c_36_4,c_36_3,c_36_2,c_36_1,c_36_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_36_lo = {c_36_15,c_36_14,c_36_13,c_36_12,c_36_11,c_36_10,c_36_9,c_36_8,io_out_36_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_36_hi_lo = {c_36_23,c_36_22,c_36_21,c_36_20,c_36_19,c_36_18,c_36_17,c_36_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_36_hi = {c_36_32,c_36_31,c_36_30,c_36_29,c_36_28,c_36_27,c_36_26,c_36_25,c_36_24,io_out_36_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_37_0 = io_in_0[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_1 = io_in_1[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_2 = io_in_2[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_3 = io_in_3[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_4 = io_in_4[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_5 = io_in_5[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_6 = io_in_6[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_7 = io_in_7[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_8 = io_in_8[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_9 = io_in_9[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_10 = io_in_10[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_11 = io_in_11[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_12 = io_in_12[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_13 = io_in_13[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_14 = io_in_14[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_15 = io_in_15[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_16 = io_in_16[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_17 = io_in_17[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_18 = io_in_18[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_19 = io_in_19[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_20 = io_in_20[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_21 = io_in_21[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_22 = io_in_22[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_23 = io_in_23[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_24 = io_in_24[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_25 = io_in_25[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_26 = io_in_26[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_27 = io_in_27[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_28 = io_in_28[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_29 = io_in_29[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_30 = io_in_30[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_31 = io_in_31[37]; // @[WallaceTest.scala 105:23]
  wire  c_37_32 = io_in_32[37]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_37_lo_lo = {c_37_7,c_37_6,c_37_5,c_37_4,c_37_3,c_37_2,c_37_1,c_37_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_37_lo = {c_37_15,c_37_14,c_37_13,c_37_12,c_37_11,c_37_10,c_37_9,c_37_8,io_out_37_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_37_hi_lo = {c_37_23,c_37_22,c_37_21,c_37_20,c_37_19,c_37_18,c_37_17,c_37_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_37_hi = {c_37_32,c_37_31,c_37_30,c_37_29,c_37_28,c_37_27,c_37_26,c_37_25,c_37_24,io_out_37_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_38_0 = io_in_0[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_1 = io_in_1[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_2 = io_in_2[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_3 = io_in_3[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_4 = io_in_4[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_5 = io_in_5[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_6 = io_in_6[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_7 = io_in_7[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_8 = io_in_8[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_9 = io_in_9[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_10 = io_in_10[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_11 = io_in_11[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_12 = io_in_12[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_13 = io_in_13[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_14 = io_in_14[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_15 = io_in_15[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_16 = io_in_16[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_17 = io_in_17[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_18 = io_in_18[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_19 = io_in_19[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_20 = io_in_20[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_21 = io_in_21[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_22 = io_in_22[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_23 = io_in_23[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_24 = io_in_24[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_25 = io_in_25[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_26 = io_in_26[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_27 = io_in_27[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_28 = io_in_28[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_29 = io_in_29[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_30 = io_in_30[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_31 = io_in_31[38]; // @[WallaceTest.scala 105:23]
  wire  c_38_32 = io_in_32[38]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_38_lo_lo = {c_38_7,c_38_6,c_38_5,c_38_4,c_38_3,c_38_2,c_38_1,c_38_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_38_lo = {c_38_15,c_38_14,c_38_13,c_38_12,c_38_11,c_38_10,c_38_9,c_38_8,io_out_38_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_38_hi_lo = {c_38_23,c_38_22,c_38_21,c_38_20,c_38_19,c_38_18,c_38_17,c_38_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_38_hi = {c_38_32,c_38_31,c_38_30,c_38_29,c_38_28,c_38_27,c_38_26,c_38_25,c_38_24,io_out_38_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_39_0 = io_in_0[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_1 = io_in_1[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_2 = io_in_2[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_3 = io_in_3[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_4 = io_in_4[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_5 = io_in_5[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_6 = io_in_6[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_7 = io_in_7[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_8 = io_in_8[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_9 = io_in_9[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_10 = io_in_10[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_11 = io_in_11[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_12 = io_in_12[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_13 = io_in_13[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_14 = io_in_14[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_15 = io_in_15[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_16 = io_in_16[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_17 = io_in_17[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_18 = io_in_18[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_19 = io_in_19[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_20 = io_in_20[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_21 = io_in_21[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_22 = io_in_22[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_23 = io_in_23[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_24 = io_in_24[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_25 = io_in_25[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_26 = io_in_26[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_27 = io_in_27[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_28 = io_in_28[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_29 = io_in_29[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_30 = io_in_30[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_31 = io_in_31[39]; // @[WallaceTest.scala 105:23]
  wire  c_39_32 = io_in_32[39]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_39_lo_lo = {c_39_7,c_39_6,c_39_5,c_39_4,c_39_3,c_39_2,c_39_1,c_39_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_39_lo = {c_39_15,c_39_14,c_39_13,c_39_12,c_39_11,c_39_10,c_39_9,c_39_8,io_out_39_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_39_hi_lo = {c_39_23,c_39_22,c_39_21,c_39_20,c_39_19,c_39_18,c_39_17,c_39_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_39_hi = {c_39_32,c_39_31,c_39_30,c_39_29,c_39_28,c_39_27,c_39_26,c_39_25,c_39_24,io_out_39_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_40_0 = io_in_0[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_1 = io_in_1[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_2 = io_in_2[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_3 = io_in_3[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_4 = io_in_4[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_5 = io_in_5[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_6 = io_in_6[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_7 = io_in_7[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_8 = io_in_8[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_9 = io_in_9[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_10 = io_in_10[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_11 = io_in_11[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_12 = io_in_12[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_13 = io_in_13[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_14 = io_in_14[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_15 = io_in_15[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_16 = io_in_16[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_17 = io_in_17[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_18 = io_in_18[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_19 = io_in_19[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_20 = io_in_20[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_21 = io_in_21[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_22 = io_in_22[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_23 = io_in_23[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_24 = io_in_24[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_25 = io_in_25[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_26 = io_in_26[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_27 = io_in_27[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_28 = io_in_28[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_29 = io_in_29[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_30 = io_in_30[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_31 = io_in_31[40]; // @[WallaceTest.scala 105:23]
  wire  c_40_32 = io_in_32[40]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_40_lo_lo = {c_40_7,c_40_6,c_40_5,c_40_4,c_40_3,c_40_2,c_40_1,c_40_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_40_lo = {c_40_15,c_40_14,c_40_13,c_40_12,c_40_11,c_40_10,c_40_9,c_40_8,io_out_40_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_40_hi_lo = {c_40_23,c_40_22,c_40_21,c_40_20,c_40_19,c_40_18,c_40_17,c_40_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_40_hi = {c_40_32,c_40_31,c_40_30,c_40_29,c_40_28,c_40_27,c_40_26,c_40_25,c_40_24,io_out_40_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_41_0 = io_in_0[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_1 = io_in_1[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_2 = io_in_2[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_3 = io_in_3[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_4 = io_in_4[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_5 = io_in_5[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_6 = io_in_6[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_7 = io_in_7[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_8 = io_in_8[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_9 = io_in_9[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_10 = io_in_10[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_11 = io_in_11[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_12 = io_in_12[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_13 = io_in_13[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_14 = io_in_14[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_15 = io_in_15[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_16 = io_in_16[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_17 = io_in_17[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_18 = io_in_18[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_19 = io_in_19[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_20 = io_in_20[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_21 = io_in_21[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_22 = io_in_22[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_23 = io_in_23[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_24 = io_in_24[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_25 = io_in_25[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_26 = io_in_26[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_27 = io_in_27[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_28 = io_in_28[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_29 = io_in_29[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_30 = io_in_30[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_31 = io_in_31[41]; // @[WallaceTest.scala 105:23]
  wire  c_41_32 = io_in_32[41]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_41_lo_lo = {c_41_7,c_41_6,c_41_5,c_41_4,c_41_3,c_41_2,c_41_1,c_41_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_41_lo = {c_41_15,c_41_14,c_41_13,c_41_12,c_41_11,c_41_10,c_41_9,c_41_8,io_out_41_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_41_hi_lo = {c_41_23,c_41_22,c_41_21,c_41_20,c_41_19,c_41_18,c_41_17,c_41_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_41_hi = {c_41_32,c_41_31,c_41_30,c_41_29,c_41_28,c_41_27,c_41_26,c_41_25,c_41_24,io_out_41_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_42_0 = io_in_0[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_1 = io_in_1[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_2 = io_in_2[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_3 = io_in_3[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_4 = io_in_4[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_5 = io_in_5[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_6 = io_in_6[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_7 = io_in_7[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_8 = io_in_8[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_9 = io_in_9[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_10 = io_in_10[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_11 = io_in_11[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_12 = io_in_12[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_13 = io_in_13[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_14 = io_in_14[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_15 = io_in_15[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_16 = io_in_16[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_17 = io_in_17[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_18 = io_in_18[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_19 = io_in_19[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_20 = io_in_20[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_21 = io_in_21[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_22 = io_in_22[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_23 = io_in_23[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_24 = io_in_24[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_25 = io_in_25[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_26 = io_in_26[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_27 = io_in_27[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_28 = io_in_28[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_29 = io_in_29[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_30 = io_in_30[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_31 = io_in_31[42]; // @[WallaceTest.scala 105:23]
  wire  c_42_32 = io_in_32[42]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_42_lo_lo = {c_42_7,c_42_6,c_42_5,c_42_4,c_42_3,c_42_2,c_42_1,c_42_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_42_lo = {c_42_15,c_42_14,c_42_13,c_42_12,c_42_11,c_42_10,c_42_9,c_42_8,io_out_42_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_42_hi_lo = {c_42_23,c_42_22,c_42_21,c_42_20,c_42_19,c_42_18,c_42_17,c_42_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_42_hi = {c_42_32,c_42_31,c_42_30,c_42_29,c_42_28,c_42_27,c_42_26,c_42_25,c_42_24,io_out_42_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_43_0 = io_in_0[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_1 = io_in_1[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_2 = io_in_2[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_3 = io_in_3[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_4 = io_in_4[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_5 = io_in_5[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_6 = io_in_6[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_7 = io_in_7[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_8 = io_in_8[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_9 = io_in_9[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_10 = io_in_10[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_11 = io_in_11[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_12 = io_in_12[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_13 = io_in_13[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_14 = io_in_14[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_15 = io_in_15[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_16 = io_in_16[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_17 = io_in_17[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_18 = io_in_18[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_19 = io_in_19[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_20 = io_in_20[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_21 = io_in_21[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_22 = io_in_22[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_23 = io_in_23[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_24 = io_in_24[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_25 = io_in_25[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_26 = io_in_26[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_27 = io_in_27[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_28 = io_in_28[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_29 = io_in_29[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_30 = io_in_30[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_31 = io_in_31[43]; // @[WallaceTest.scala 105:23]
  wire  c_43_32 = io_in_32[43]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_43_lo_lo = {c_43_7,c_43_6,c_43_5,c_43_4,c_43_3,c_43_2,c_43_1,c_43_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_43_lo = {c_43_15,c_43_14,c_43_13,c_43_12,c_43_11,c_43_10,c_43_9,c_43_8,io_out_43_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_43_hi_lo = {c_43_23,c_43_22,c_43_21,c_43_20,c_43_19,c_43_18,c_43_17,c_43_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_43_hi = {c_43_32,c_43_31,c_43_30,c_43_29,c_43_28,c_43_27,c_43_26,c_43_25,c_43_24,io_out_43_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_44_0 = io_in_0[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_1 = io_in_1[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_2 = io_in_2[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_3 = io_in_3[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_4 = io_in_4[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_5 = io_in_5[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_6 = io_in_6[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_7 = io_in_7[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_8 = io_in_8[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_9 = io_in_9[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_10 = io_in_10[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_11 = io_in_11[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_12 = io_in_12[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_13 = io_in_13[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_14 = io_in_14[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_15 = io_in_15[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_16 = io_in_16[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_17 = io_in_17[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_18 = io_in_18[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_19 = io_in_19[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_20 = io_in_20[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_21 = io_in_21[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_22 = io_in_22[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_23 = io_in_23[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_24 = io_in_24[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_25 = io_in_25[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_26 = io_in_26[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_27 = io_in_27[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_28 = io_in_28[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_29 = io_in_29[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_30 = io_in_30[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_31 = io_in_31[44]; // @[WallaceTest.scala 105:23]
  wire  c_44_32 = io_in_32[44]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_44_lo_lo = {c_44_7,c_44_6,c_44_5,c_44_4,c_44_3,c_44_2,c_44_1,c_44_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_44_lo = {c_44_15,c_44_14,c_44_13,c_44_12,c_44_11,c_44_10,c_44_9,c_44_8,io_out_44_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_44_hi_lo = {c_44_23,c_44_22,c_44_21,c_44_20,c_44_19,c_44_18,c_44_17,c_44_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_44_hi = {c_44_32,c_44_31,c_44_30,c_44_29,c_44_28,c_44_27,c_44_26,c_44_25,c_44_24,io_out_44_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_45_0 = io_in_0[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_1 = io_in_1[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_2 = io_in_2[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_3 = io_in_3[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_4 = io_in_4[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_5 = io_in_5[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_6 = io_in_6[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_7 = io_in_7[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_8 = io_in_8[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_9 = io_in_9[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_10 = io_in_10[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_11 = io_in_11[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_12 = io_in_12[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_13 = io_in_13[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_14 = io_in_14[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_15 = io_in_15[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_16 = io_in_16[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_17 = io_in_17[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_18 = io_in_18[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_19 = io_in_19[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_20 = io_in_20[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_21 = io_in_21[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_22 = io_in_22[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_23 = io_in_23[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_24 = io_in_24[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_25 = io_in_25[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_26 = io_in_26[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_27 = io_in_27[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_28 = io_in_28[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_29 = io_in_29[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_30 = io_in_30[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_31 = io_in_31[45]; // @[WallaceTest.scala 105:23]
  wire  c_45_32 = io_in_32[45]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_45_lo_lo = {c_45_7,c_45_6,c_45_5,c_45_4,c_45_3,c_45_2,c_45_1,c_45_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_45_lo = {c_45_15,c_45_14,c_45_13,c_45_12,c_45_11,c_45_10,c_45_9,c_45_8,io_out_45_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_45_hi_lo = {c_45_23,c_45_22,c_45_21,c_45_20,c_45_19,c_45_18,c_45_17,c_45_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_45_hi = {c_45_32,c_45_31,c_45_30,c_45_29,c_45_28,c_45_27,c_45_26,c_45_25,c_45_24,io_out_45_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_46_0 = io_in_0[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_1 = io_in_1[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_2 = io_in_2[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_3 = io_in_3[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_4 = io_in_4[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_5 = io_in_5[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_6 = io_in_6[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_7 = io_in_7[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_8 = io_in_8[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_9 = io_in_9[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_10 = io_in_10[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_11 = io_in_11[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_12 = io_in_12[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_13 = io_in_13[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_14 = io_in_14[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_15 = io_in_15[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_16 = io_in_16[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_17 = io_in_17[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_18 = io_in_18[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_19 = io_in_19[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_20 = io_in_20[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_21 = io_in_21[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_22 = io_in_22[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_23 = io_in_23[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_24 = io_in_24[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_25 = io_in_25[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_26 = io_in_26[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_27 = io_in_27[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_28 = io_in_28[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_29 = io_in_29[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_30 = io_in_30[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_31 = io_in_31[46]; // @[WallaceTest.scala 105:23]
  wire  c_46_32 = io_in_32[46]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_46_lo_lo = {c_46_7,c_46_6,c_46_5,c_46_4,c_46_3,c_46_2,c_46_1,c_46_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_46_lo = {c_46_15,c_46_14,c_46_13,c_46_12,c_46_11,c_46_10,c_46_9,c_46_8,io_out_46_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_46_hi_lo = {c_46_23,c_46_22,c_46_21,c_46_20,c_46_19,c_46_18,c_46_17,c_46_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_46_hi = {c_46_32,c_46_31,c_46_30,c_46_29,c_46_28,c_46_27,c_46_26,c_46_25,c_46_24,io_out_46_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_47_0 = io_in_0[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_1 = io_in_1[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_2 = io_in_2[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_3 = io_in_3[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_4 = io_in_4[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_5 = io_in_5[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_6 = io_in_6[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_7 = io_in_7[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_8 = io_in_8[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_9 = io_in_9[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_10 = io_in_10[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_11 = io_in_11[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_12 = io_in_12[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_13 = io_in_13[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_14 = io_in_14[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_15 = io_in_15[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_16 = io_in_16[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_17 = io_in_17[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_18 = io_in_18[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_19 = io_in_19[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_20 = io_in_20[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_21 = io_in_21[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_22 = io_in_22[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_23 = io_in_23[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_24 = io_in_24[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_25 = io_in_25[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_26 = io_in_26[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_27 = io_in_27[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_28 = io_in_28[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_29 = io_in_29[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_30 = io_in_30[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_31 = io_in_31[47]; // @[WallaceTest.scala 105:23]
  wire  c_47_32 = io_in_32[47]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_47_lo_lo = {c_47_7,c_47_6,c_47_5,c_47_4,c_47_3,c_47_2,c_47_1,c_47_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_47_lo = {c_47_15,c_47_14,c_47_13,c_47_12,c_47_11,c_47_10,c_47_9,c_47_8,io_out_47_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_47_hi_lo = {c_47_23,c_47_22,c_47_21,c_47_20,c_47_19,c_47_18,c_47_17,c_47_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_47_hi = {c_47_32,c_47_31,c_47_30,c_47_29,c_47_28,c_47_27,c_47_26,c_47_25,c_47_24,io_out_47_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_48_0 = io_in_0[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_1 = io_in_1[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_2 = io_in_2[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_3 = io_in_3[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_4 = io_in_4[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_5 = io_in_5[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_6 = io_in_6[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_7 = io_in_7[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_8 = io_in_8[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_9 = io_in_9[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_10 = io_in_10[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_11 = io_in_11[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_12 = io_in_12[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_13 = io_in_13[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_14 = io_in_14[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_15 = io_in_15[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_16 = io_in_16[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_17 = io_in_17[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_18 = io_in_18[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_19 = io_in_19[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_20 = io_in_20[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_21 = io_in_21[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_22 = io_in_22[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_23 = io_in_23[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_24 = io_in_24[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_25 = io_in_25[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_26 = io_in_26[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_27 = io_in_27[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_28 = io_in_28[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_29 = io_in_29[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_30 = io_in_30[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_31 = io_in_31[48]; // @[WallaceTest.scala 105:23]
  wire  c_48_32 = io_in_32[48]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_48_lo_lo = {c_48_7,c_48_6,c_48_5,c_48_4,c_48_3,c_48_2,c_48_1,c_48_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_48_lo = {c_48_15,c_48_14,c_48_13,c_48_12,c_48_11,c_48_10,c_48_9,c_48_8,io_out_48_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_48_hi_lo = {c_48_23,c_48_22,c_48_21,c_48_20,c_48_19,c_48_18,c_48_17,c_48_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_48_hi = {c_48_32,c_48_31,c_48_30,c_48_29,c_48_28,c_48_27,c_48_26,c_48_25,c_48_24,io_out_48_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_49_0 = io_in_0[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_1 = io_in_1[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_2 = io_in_2[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_3 = io_in_3[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_4 = io_in_4[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_5 = io_in_5[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_6 = io_in_6[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_7 = io_in_7[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_8 = io_in_8[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_9 = io_in_9[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_10 = io_in_10[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_11 = io_in_11[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_12 = io_in_12[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_13 = io_in_13[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_14 = io_in_14[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_15 = io_in_15[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_16 = io_in_16[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_17 = io_in_17[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_18 = io_in_18[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_19 = io_in_19[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_20 = io_in_20[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_21 = io_in_21[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_22 = io_in_22[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_23 = io_in_23[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_24 = io_in_24[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_25 = io_in_25[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_26 = io_in_26[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_27 = io_in_27[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_28 = io_in_28[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_29 = io_in_29[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_30 = io_in_30[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_31 = io_in_31[49]; // @[WallaceTest.scala 105:23]
  wire  c_49_32 = io_in_32[49]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_49_lo_lo = {c_49_7,c_49_6,c_49_5,c_49_4,c_49_3,c_49_2,c_49_1,c_49_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_49_lo = {c_49_15,c_49_14,c_49_13,c_49_12,c_49_11,c_49_10,c_49_9,c_49_8,io_out_49_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_49_hi_lo = {c_49_23,c_49_22,c_49_21,c_49_20,c_49_19,c_49_18,c_49_17,c_49_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_49_hi = {c_49_32,c_49_31,c_49_30,c_49_29,c_49_28,c_49_27,c_49_26,c_49_25,c_49_24,io_out_49_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_50_0 = io_in_0[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_1 = io_in_1[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_2 = io_in_2[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_3 = io_in_3[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_4 = io_in_4[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_5 = io_in_5[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_6 = io_in_6[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_7 = io_in_7[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_8 = io_in_8[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_9 = io_in_9[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_10 = io_in_10[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_11 = io_in_11[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_12 = io_in_12[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_13 = io_in_13[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_14 = io_in_14[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_15 = io_in_15[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_16 = io_in_16[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_17 = io_in_17[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_18 = io_in_18[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_19 = io_in_19[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_20 = io_in_20[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_21 = io_in_21[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_22 = io_in_22[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_23 = io_in_23[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_24 = io_in_24[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_25 = io_in_25[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_26 = io_in_26[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_27 = io_in_27[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_28 = io_in_28[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_29 = io_in_29[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_30 = io_in_30[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_31 = io_in_31[50]; // @[WallaceTest.scala 105:23]
  wire  c_50_32 = io_in_32[50]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_50_lo_lo = {c_50_7,c_50_6,c_50_5,c_50_4,c_50_3,c_50_2,c_50_1,c_50_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_50_lo = {c_50_15,c_50_14,c_50_13,c_50_12,c_50_11,c_50_10,c_50_9,c_50_8,io_out_50_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_50_hi_lo = {c_50_23,c_50_22,c_50_21,c_50_20,c_50_19,c_50_18,c_50_17,c_50_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_50_hi = {c_50_32,c_50_31,c_50_30,c_50_29,c_50_28,c_50_27,c_50_26,c_50_25,c_50_24,io_out_50_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_51_0 = io_in_0[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_1 = io_in_1[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_2 = io_in_2[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_3 = io_in_3[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_4 = io_in_4[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_5 = io_in_5[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_6 = io_in_6[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_7 = io_in_7[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_8 = io_in_8[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_9 = io_in_9[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_10 = io_in_10[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_11 = io_in_11[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_12 = io_in_12[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_13 = io_in_13[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_14 = io_in_14[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_15 = io_in_15[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_16 = io_in_16[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_17 = io_in_17[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_18 = io_in_18[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_19 = io_in_19[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_20 = io_in_20[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_21 = io_in_21[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_22 = io_in_22[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_23 = io_in_23[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_24 = io_in_24[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_25 = io_in_25[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_26 = io_in_26[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_27 = io_in_27[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_28 = io_in_28[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_29 = io_in_29[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_30 = io_in_30[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_31 = io_in_31[51]; // @[WallaceTest.scala 105:23]
  wire  c_51_32 = io_in_32[51]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_51_lo_lo = {c_51_7,c_51_6,c_51_5,c_51_4,c_51_3,c_51_2,c_51_1,c_51_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_51_lo = {c_51_15,c_51_14,c_51_13,c_51_12,c_51_11,c_51_10,c_51_9,c_51_8,io_out_51_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_51_hi_lo = {c_51_23,c_51_22,c_51_21,c_51_20,c_51_19,c_51_18,c_51_17,c_51_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_51_hi = {c_51_32,c_51_31,c_51_30,c_51_29,c_51_28,c_51_27,c_51_26,c_51_25,c_51_24,io_out_51_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_52_0 = io_in_0[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_1 = io_in_1[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_2 = io_in_2[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_3 = io_in_3[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_4 = io_in_4[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_5 = io_in_5[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_6 = io_in_6[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_7 = io_in_7[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_8 = io_in_8[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_9 = io_in_9[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_10 = io_in_10[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_11 = io_in_11[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_12 = io_in_12[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_13 = io_in_13[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_14 = io_in_14[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_15 = io_in_15[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_16 = io_in_16[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_17 = io_in_17[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_18 = io_in_18[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_19 = io_in_19[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_20 = io_in_20[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_21 = io_in_21[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_22 = io_in_22[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_23 = io_in_23[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_24 = io_in_24[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_25 = io_in_25[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_26 = io_in_26[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_27 = io_in_27[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_28 = io_in_28[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_29 = io_in_29[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_30 = io_in_30[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_31 = io_in_31[52]; // @[WallaceTest.scala 105:23]
  wire  c_52_32 = io_in_32[52]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_52_lo_lo = {c_52_7,c_52_6,c_52_5,c_52_4,c_52_3,c_52_2,c_52_1,c_52_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_52_lo = {c_52_15,c_52_14,c_52_13,c_52_12,c_52_11,c_52_10,c_52_9,c_52_8,io_out_52_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_52_hi_lo = {c_52_23,c_52_22,c_52_21,c_52_20,c_52_19,c_52_18,c_52_17,c_52_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_52_hi = {c_52_32,c_52_31,c_52_30,c_52_29,c_52_28,c_52_27,c_52_26,c_52_25,c_52_24,io_out_52_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_53_0 = io_in_0[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_1 = io_in_1[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_2 = io_in_2[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_3 = io_in_3[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_4 = io_in_4[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_5 = io_in_5[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_6 = io_in_6[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_7 = io_in_7[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_8 = io_in_8[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_9 = io_in_9[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_10 = io_in_10[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_11 = io_in_11[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_12 = io_in_12[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_13 = io_in_13[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_14 = io_in_14[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_15 = io_in_15[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_16 = io_in_16[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_17 = io_in_17[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_18 = io_in_18[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_19 = io_in_19[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_20 = io_in_20[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_21 = io_in_21[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_22 = io_in_22[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_23 = io_in_23[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_24 = io_in_24[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_25 = io_in_25[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_26 = io_in_26[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_27 = io_in_27[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_28 = io_in_28[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_29 = io_in_29[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_30 = io_in_30[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_31 = io_in_31[53]; // @[WallaceTest.scala 105:23]
  wire  c_53_32 = io_in_32[53]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_53_lo_lo = {c_53_7,c_53_6,c_53_5,c_53_4,c_53_3,c_53_2,c_53_1,c_53_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_53_lo = {c_53_15,c_53_14,c_53_13,c_53_12,c_53_11,c_53_10,c_53_9,c_53_8,io_out_53_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_53_hi_lo = {c_53_23,c_53_22,c_53_21,c_53_20,c_53_19,c_53_18,c_53_17,c_53_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_53_hi = {c_53_32,c_53_31,c_53_30,c_53_29,c_53_28,c_53_27,c_53_26,c_53_25,c_53_24,io_out_53_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_54_0 = io_in_0[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_1 = io_in_1[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_2 = io_in_2[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_3 = io_in_3[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_4 = io_in_4[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_5 = io_in_5[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_6 = io_in_6[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_7 = io_in_7[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_8 = io_in_8[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_9 = io_in_9[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_10 = io_in_10[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_11 = io_in_11[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_12 = io_in_12[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_13 = io_in_13[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_14 = io_in_14[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_15 = io_in_15[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_16 = io_in_16[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_17 = io_in_17[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_18 = io_in_18[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_19 = io_in_19[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_20 = io_in_20[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_21 = io_in_21[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_22 = io_in_22[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_23 = io_in_23[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_24 = io_in_24[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_25 = io_in_25[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_26 = io_in_26[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_27 = io_in_27[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_28 = io_in_28[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_29 = io_in_29[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_30 = io_in_30[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_31 = io_in_31[54]; // @[WallaceTest.scala 105:23]
  wire  c_54_32 = io_in_32[54]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_54_lo_lo = {c_54_7,c_54_6,c_54_5,c_54_4,c_54_3,c_54_2,c_54_1,c_54_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_54_lo = {c_54_15,c_54_14,c_54_13,c_54_12,c_54_11,c_54_10,c_54_9,c_54_8,io_out_54_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_54_hi_lo = {c_54_23,c_54_22,c_54_21,c_54_20,c_54_19,c_54_18,c_54_17,c_54_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_54_hi = {c_54_32,c_54_31,c_54_30,c_54_29,c_54_28,c_54_27,c_54_26,c_54_25,c_54_24,io_out_54_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_55_0 = io_in_0[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_1 = io_in_1[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_2 = io_in_2[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_3 = io_in_3[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_4 = io_in_4[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_5 = io_in_5[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_6 = io_in_6[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_7 = io_in_7[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_8 = io_in_8[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_9 = io_in_9[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_10 = io_in_10[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_11 = io_in_11[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_12 = io_in_12[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_13 = io_in_13[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_14 = io_in_14[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_15 = io_in_15[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_16 = io_in_16[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_17 = io_in_17[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_18 = io_in_18[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_19 = io_in_19[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_20 = io_in_20[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_21 = io_in_21[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_22 = io_in_22[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_23 = io_in_23[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_24 = io_in_24[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_25 = io_in_25[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_26 = io_in_26[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_27 = io_in_27[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_28 = io_in_28[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_29 = io_in_29[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_30 = io_in_30[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_31 = io_in_31[55]; // @[WallaceTest.scala 105:23]
  wire  c_55_32 = io_in_32[55]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_55_lo_lo = {c_55_7,c_55_6,c_55_5,c_55_4,c_55_3,c_55_2,c_55_1,c_55_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_55_lo = {c_55_15,c_55_14,c_55_13,c_55_12,c_55_11,c_55_10,c_55_9,c_55_8,io_out_55_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_55_hi_lo = {c_55_23,c_55_22,c_55_21,c_55_20,c_55_19,c_55_18,c_55_17,c_55_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_55_hi = {c_55_32,c_55_31,c_55_30,c_55_29,c_55_28,c_55_27,c_55_26,c_55_25,c_55_24,io_out_55_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_56_0 = io_in_0[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_1 = io_in_1[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_2 = io_in_2[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_3 = io_in_3[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_4 = io_in_4[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_5 = io_in_5[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_6 = io_in_6[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_7 = io_in_7[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_8 = io_in_8[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_9 = io_in_9[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_10 = io_in_10[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_11 = io_in_11[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_12 = io_in_12[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_13 = io_in_13[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_14 = io_in_14[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_15 = io_in_15[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_16 = io_in_16[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_17 = io_in_17[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_18 = io_in_18[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_19 = io_in_19[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_20 = io_in_20[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_21 = io_in_21[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_22 = io_in_22[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_23 = io_in_23[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_24 = io_in_24[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_25 = io_in_25[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_26 = io_in_26[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_27 = io_in_27[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_28 = io_in_28[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_29 = io_in_29[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_30 = io_in_30[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_31 = io_in_31[56]; // @[WallaceTest.scala 105:23]
  wire  c_56_32 = io_in_32[56]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_56_lo_lo = {c_56_7,c_56_6,c_56_5,c_56_4,c_56_3,c_56_2,c_56_1,c_56_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_56_lo = {c_56_15,c_56_14,c_56_13,c_56_12,c_56_11,c_56_10,c_56_9,c_56_8,io_out_56_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_56_hi_lo = {c_56_23,c_56_22,c_56_21,c_56_20,c_56_19,c_56_18,c_56_17,c_56_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_56_hi = {c_56_32,c_56_31,c_56_30,c_56_29,c_56_28,c_56_27,c_56_26,c_56_25,c_56_24,io_out_56_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_57_0 = io_in_0[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_1 = io_in_1[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_2 = io_in_2[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_3 = io_in_3[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_4 = io_in_4[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_5 = io_in_5[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_6 = io_in_6[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_7 = io_in_7[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_8 = io_in_8[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_9 = io_in_9[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_10 = io_in_10[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_11 = io_in_11[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_12 = io_in_12[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_13 = io_in_13[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_14 = io_in_14[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_15 = io_in_15[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_16 = io_in_16[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_17 = io_in_17[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_18 = io_in_18[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_19 = io_in_19[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_20 = io_in_20[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_21 = io_in_21[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_22 = io_in_22[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_23 = io_in_23[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_24 = io_in_24[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_25 = io_in_25[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_26 = io_in_26[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_27 = io_in_27[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_28 = io_in_28[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_29 = io_in_29[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_30 = io_in_30[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_31 = io_in_31[57]; // @[WallaceTest.scala 105:23]
  wire  c_57_32 = io_in_32[57]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_57_lo_lo = {c_57_7,c_57_6,c_57_5,c_57_4,c_57_3,c_57_2,c_57_1,c_57_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_57_lo = {c_57_15,c_57_14,c_57_13,c_57_12,c_57_11,c_57_10,c_57_9,c_57_8,io_out_57_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_57_hi_lo = {c_57_23,c_57_22,c_57_21,c_57_20,c_57_19,c_57_18,c_57_17,c_57_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_57_hi = {c_57_32,c_57_31,c_57_30,c_57_29,c_57_28,c_57_27,c_57_26,c_57_25,c_57_24,io_out_57_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_58_0 = io_in_0[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_1 = io_in_1[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_2 = io_in_2[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_3 = io_in_3[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_4 = io_in_4[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_5 = io_in_5[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_6 = io_in_6[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_7 = io_in_7[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_8 = io_in_8[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_9 = io_in_9[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_10 = io_in_10[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_11 = io_in_11[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_12 = io_in_12[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_13 = io_in_13[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_14 = io_in_14[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_15 = io_in_15[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_16 = io_in_16[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_17 = io_in_17[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_18 = io_in_18[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_19 = io_in_19[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_20 = io_in_20[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_21 = io_in_21[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_22 = io_in_22[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_23 = io_in_23[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_24 = io_in_24[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_25 = io_in_25[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_26 = io_in_26[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_27 = io_in_27[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_28 = io_in_28[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_29 = io_in_29[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_30 = io_in_30[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_31 = io_in_31[58]; // @[WallaceTest.scala 105:23]
  wire  c_58_32 = io_in_32[58]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_58_lo_lo = {c_58_7,c_58_6,c_58_5,c_58_4,c_58_3,c_58_2,c_58_1,c_58_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_58_lo = {c_58_15,c_58_14,c_58_13,c_58_12,c_58_11,c_58_10,c_58_9,c_58_8,io_out_58_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_58_hi_lo = {c_58_23,c_58_22,c_58_21,c_58_20,c_58_19,c_58_18,c_58_17,c_58_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_58_hi = {c_58_32,c_58_31,c_58_30,c_58_29,c_58_28,c_58_27,c_58_26,c_58_25,c_58_24,io_out_58_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_59_0 = io_in_0[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_1 = io_in_1[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_2 = io_in_2[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_3 = io_in_3[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_4 = io_in_4[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_5 = io_in_5[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_6 = io_in_6[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_7 = io_in_7[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_8 = io_in_8[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_9 = io_in_9[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_10 = io_in_10[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_11 = io_in_11[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_12 = io_in_12[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_13 = io_in_13[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_14 = io_in_14[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_15 = io_in_15[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_16 = io_in_16[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_17 = io_in_17[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_18 = io_in_18[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_19 = io_in_19[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_20 = io_in_20[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_21 = io_in_21[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_22 = io_in_22[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_23 = io_in_23[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_24 = io_in_24[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_25 = io_in_25[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_26 = io_in_26[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_27 = io_in_27[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_28 = io_in_28[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_29 = io_in_29[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_30 = io_in_30[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_31 = io_in_31[59]; // @[WallaceTest.scala 105:23]
  wire  c_59_32 = io_in_32[59]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_59_lo_lo = {c_59_7,c_59_6,c_59_5,c_59_4,c_59_3,c_59_2,c_59_1,c_59_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_59_lo = {c_59_15,c_59_14,c_59_13,c_59_12,c_59_11,c_59_10,c_59_9,c_59_8,io_out_59_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_59_hi_lo = {c_59_23,c_59_22,c_59_21,c_59_20,c_59_19,c_59_18,c_59_17,c_59_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_59_hi = {c_59_32,c_59_31,c_59_30,c_59_29,c_59_28,c_59_27,c_59_26,c_59_25,c_59_24,io_out_59_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_60_0 = io_in_0[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_1 = io_in_1[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_2 = io_in_2[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_3 = io_in_3[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_4 = io_in_4[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_5 = io_in_5[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_6 = io_in_6[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_7 = io_in_7[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_8 = io_in_8[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_9 = io_in_9[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_10 = io_in_10[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_11 = io_in_11[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_12 = io_in_12[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_13 = io_in_13[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_14 = io_in_14[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_15 = io_in_15[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_16 = io_in_16[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_17 = io_in_17[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_18 = io_in_18[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_19 = io_in_19[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_20 = io_in_20[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_21 = io_in_21[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_22 = io_in_22[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_23 = io_in_23[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_24 = io_in_24[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_25 = io_in_25[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_26 = io_in_26[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_27 = io_in_27[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_28 = io_in_28[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_29 = io_in_29[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_30 = io_in_30[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_31 = io_in_31[60]; // @[WallaceTest.scala 105:23]
  wire  c_60_32 = io_in_32[60]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_60_lo_lo = {c_60_7,c_60_6,c_60_5,c_60_4,c_60_3,c_60_2,c_60_1,c_60_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_60_lo = {c_60_15,c_60_14,c_60_13,c_60_12,c_60_11,c_60_10,c_60_9,c_60_8,io_out_60_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_60_hi_lo = {c_60_23,c_60_22,c_60_21,c_60_20,c_60_19,c_60_18,c_60_17,c_60_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_60_hi = {c_60_32,c_60_31,c_60_30,c_60_29,c_60_28,c_60_27,c_60_26,c_60_25,c_60_24,io_out_60_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_61_0 = io_in_0[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_1 = io_in_1[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_2 = io_in_2[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_3 = io_in_3[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_4 = io_in_4[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_5 = io_in_5[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_6 = io_in_6[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_7 = io_in_7[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_8 = io_in_8[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_9 = io_in_9[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_10 = io_in_10[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_11 = io_in_11[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_12 = io_in_12[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_13 = io_in_13[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_14 = io_in_14[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_15 = io_in_15[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_16 = io_in_16[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_17 = io_in_17[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_18 = io_in_18[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_19 = io_in_19[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_20 = io_in_20[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_21 = io_in_21[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_22 = io_in_22[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_23 = io_in_23[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_24 = io_in_24[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_25 = io_in_25[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_26 = io_in_26[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_27 = io_in_27[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_28 = io_in_28[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_29 = io_in_29[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_30 = io_in_30[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_31 = io_in_31[61]; // @[WallaceTest.scala 105:23]
  wire  c_61_32 = io_in_32[61]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_61_lo_lo = {c_61_7,c_61_6,c_61_5,c_61_4,c_61_3,c_61_2,c_61_1,c_61_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_61_lo = {c_61_15,c_61_14,c_61_13,c_61_12,c_61_11,c_61_10,c_61_9,c_61_8,io_out_61_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_61_hi_lo = {c_61_23,c_61_22,c_61_21,c_61_20,c_61_19,c_61_18,c_61_17,c_61_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_61_hi = {c_61_32,c_61_31,c_61_30,c_61_29,c_61_28,c_61_27,c_61_26,c_61_25,c_61_24,io_out_61_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_62_0 = io_in_0[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_1 = io_in_1[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_2 = io_in_2[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_3 = io_in_3[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_4 = io_in_4[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_5 = io_in_5[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_6 = io_in_6[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_7 = io_in_7[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_8 = io_in_8[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_9 = io_in_9[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_10 = io_in_10[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_11 = io_in_11[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_12 = io_in_12[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_13 = io_in_13[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_14 = io_in_14[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_15 = io_in_15[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_16 = io_in_16[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_17 = io_in_17[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_18 = io_in_18[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_19 = io_in_19[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_20 = io_in_20[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_21 = io_in_21[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_22 = io_in_22[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_23 = io_in_23[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_24 = io_in_24[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_25 = io_in_25[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_26 = io_in_26[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_27 = io_in_27[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_28 = io_in_28[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_29 = io_in_29[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_30 = io_in_30[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_31 = io_in_31[62]; // @[WallaceTest.scala 105:23]
  wire  c_62_32 = io_in_32[62]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_62_lo_lo = {c_62_7,c_62_6,c_62_5,c_62_4,c_62_3,c_62_2,c_62_1,c_62_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_62_lo = {c_62_15,c_62_14,c_62_13,c_62_12,c_62_11,c_62_10,c_62_9,c_62_8,io_out_62_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_62_hi_lo = {c_62_23,c_62_22,c_62_21,c_62_20,c_62_19,c_62_18,c_62_17,c_62_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_62_hi = {c_62_32,c_62_31,c_62_30,c_62_29,c_62_28,c_62_27,c_62_26,c_62_25,c_62_24,io_out_62_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_63_0 = io_in_0[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_1 = io_in_1[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_2 = io_in_2[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_3 = io_in_3[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_4 = io_in_4[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_5 = io_in_5[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_6 = io_in_6[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_7 = io_in_7[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_8 = io_in_8[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_9 = io_in_9[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_10 = io_in_10[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_11 = io_in_11[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_12 = io_in_12[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_13 = io_in_13[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_14 = io_in_14[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_15 = io_in_15[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_16 = io_in_16[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_17 = io_in_17[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_18 = io_in_18[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_19 = io_in_19[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_20 = io_in_20[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_21 = io_in_21[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_22 = io_in_22[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_23 = io_in_23[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_24 = io_in_24[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_25 = io_in_25[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_26 = io_in_26[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_27 = io_in_27[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_28 = io_in_28[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_29 = io_in_29[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_30 = io_in_30[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_31 = io_in_31[63]; // @[WallaceTest.scala 105:23]
  wire  c_63_32 = io_in_32[63]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_63_lo_lo = {c_63_7,c_63_6,c_63_5,c_63_4,c_63_3,c_63_2,c_63_1,c_63_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_63_lo = {c_63_15,c_63_14,c_63_13,c_63_12,c_63_11,c_63_10,c_63_9,c_63_8,io_out_63_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_63_hi_lo = {c_63_23,c_63_22,c_63_21,c_63_20,c_63_19,c_63_18,c_63_17,c_63_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_63_hi = {c_63_32,c_63_31,c_63_30,c_63_29,c_63_28,c_63_27,c_63_26,c_63_25,c_63_24,io_out_63_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_64_0 = io_in_0[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_1 = io_in_1[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_2 = io_in_2[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_3 = io_in_3[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_4 = io_in_4[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_5 = io_in_5[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_6 = io_in_6[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_7 = io_in_7[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_8 = io_in_8[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_9 = io_in_9[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_10 = io_in_10[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_11 = io_in_11[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_12 = io_in_12[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_13 = io_in_13[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_14 = io_in_14[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_15 = io_in_15[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_16 = io_in_16[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_17 = io_in_17[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_18 = io_in_18[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_19 = io_in_19[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_20 = io_in_20[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_21 = io_in_21[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_22 = io_in_22[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_23 = io_in_23[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_24 = io_in_24[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_25 = io_in_25[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_26 = io_in_26[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_27 = io_in_27[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_28 = io_in_28[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_29 = io_in_29[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_30 = io_in_30[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_31 = io_in_31[64]; // @[WallaceTest.scala 105:23]
  wire  c_64_32 = io_in_32[64]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_64_lo_lo = {c_64_7,c_64_6,c_64_5,c_64_4,c_64_3,c_64_2,c_64_1,c_64_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_64_lo = {c_64_15,c_64_14,c_64_13,c_64_12,c_64_11,c_64_10,c_64_9,c_64_8,io_out_64_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_64_hi_lo = {c_64_23,c_64_22,c_64_21,c_64_20,c_64_19,c_64_18,c_64_17,c_64_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_64_hi = {c_64_32,c_64_31,c_64_30,c_64_29,c_64_28,c_64_27,c_64_26,c_64_25,c_64_24,io_out_64_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_65_0 = io_in_0[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_1 = io_in_1[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_2 = io_in_2[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_3 = io_in_3[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_4 = io_in_4[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_5 = io_in_5[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_6 = io_in_6[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_7 = io_in_7[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_8 = io_in_8[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_9 = io_in_9[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_10 = io_in_10[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_11 = io_in_11[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_12 = io_in_12[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_13 = io_in_13[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_14 = io_in_14[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_15 = io_in_15[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_16 = io_in_16[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_17 = io_in_17[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_18 = io_in_18[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_19 = io_in_19[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_20 = io_in_20[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_21 = io_in_21[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_22 = io_in_22[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_23 = io_in_23[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_24 = io_in_24[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_25 = io_in_25[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_26 = io_in_26[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_27 = io_in_27[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_28 = io_in_28[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_29 = io_in_29[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_30 = io_in_30[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_31 = io_in_31[65]; // @[WallaceTest.scala 105:23]
  wire  c_65_32 = io_in_32[65]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_65_lo_lo = {c_65_7,c_65_6,c_65_5,c_65_4,c_65_3,c_65_2,c_65_1,c_65_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_65_lo = {c_65_15,c_65_14,c_65_13,c_65_12,c_65_11,c_65_10,c_65_9,c_65_8,io_out_65_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_65_hi_lo = {c_65_23,c_65_22,c_65_21,c_65_20,c_65_19,c_65_18,c_65_17,c_65_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_65_hi = {c_65_32,c_65_31,c_65_30,c_65_29,c_65_28,c_65_27,c_65_26,c_65_25,c_65_24,io_out_65_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_66_0 = io_in_0[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_1 = io_in_1[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_2 = io_in_2[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_3 = io_in_3[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_4 = io_in_4[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_5 = io_in_5[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_6 = io_in_6[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_7 = io_in_7[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_8 = io_in_8[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_9 = io_in_9[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_10 = io_in_10[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_11 = io_in_11[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_12 = io_in_12[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_13 = io_in_13[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_14 = io_in_14[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_15 = io_in_15[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_16 = io_in_16[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_17 = io_in_17[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_18 = io_in_18[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_19 = io_in_19[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_20 = io_in_20[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_21 = io_in_21[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_22 = io_in_22[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_23 = io_in_23[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_24 = io_in_24[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_25 = io_in_25[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_26 = io_in_26[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_27 = io_in_27[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_28 = io_in_28[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_29 = io_in_29[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_30 = io_in_30[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_31 = io_in_31[66]; // @[WallaceTest.scala 105:23]
  wire  c_66_32 = io_in_32[66]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_66_lo_lo = {c_66_7,c_66_6,c_66_5,c_66_4,c_66_3,c_66_2,c_66_1,c_66_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_66_lo = {c_66_15,c_66_14,c_66_13,c_66_12,c_66_11,c_66_10,c_66_9,c_66_8,io_out_66_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_66_hi_lo = {c_66_23,c_66_22,c_66_21,c_66_20,c_66_19,c_66_18,c_66_17,c_66_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_66_hi = {c_66_32,c_66_31,c_66_30,c_66_29,c_66_28,c_66_27,c_66_26,c_66_25,c_66_24,io_out_66_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_67_0 = io_in_0[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_1 = io_in_1[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_2 = io_in_2[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_3 = io_in_3[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_4 = io_in_4[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_5 = io_in_5[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_6 = io_in_6[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_7 = io_in_7[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_8 = io_in_8[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_9 = io_in_9[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_10 = io_in_10[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_11 = io_in_11[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_12 = io_in_12[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_13 = io_in_13[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_14 = io_in_14[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_15 = io_in_15[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_16 = io_in_16[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_17 = io_in_17[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_18 = io_in_18[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_19 = io_in_19[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_20 = io_in_20[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_21 = io_in_21[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_22 = io_in_22[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_23 = io_in_23[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_24 = io_in_24[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_25 = io_in_25[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_26 = io_in_26[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_27 = io_in_27[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_28 = io_in_28[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_29 = io_in_29[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_30 = io_in_30[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_31 = io_in_31[67]; // @[WallaceTest.scala 105:23]
  wire  c_67_32 = io_in_32[67]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_67_lo_lo = {c_67_7,c_67_6,c_67_5,c_67_4,c_67_3,c_67_2,c_67_1,c_67_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_67_lo = {c_67_15,c_67_14,c_67_13,c_67_12,c_67_11,c_67_10,c_67_9,c_67_8,io_out_67_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_67_hi_lo = {c_67_23,c_67_22,c_67_21,c_67_20,c_67_19,c_67_18,c_67_17,c_67_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_67_hi = {c_67_32,c_67_31,c_67_30,c_67_29,c_67_28,c_67_27,c_67_26,c_67_25,c_67_24,io_out_67_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_68_0 = io_in_0[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_1 = io_in_1[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_2 = io_in_2[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_3 = io_in_3[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_4 = io_in_4[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_5 = io_in_5[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_6 = io_in_6[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_7 = io_in_7[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_8 = io_in_8[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_9 = io_in_9[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_10 = io_in_10[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_11 = io_in_11[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_12 = io_in_12[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_13 = io_in_13[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_14 = io_in_14[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_15 = io_in_15[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_16 = io_in_16[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_17 = io_in_17[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_18 = io_in_18[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_19 = io_in_19[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_20 = io_in_20[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_21 = io_in_21[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_22 = io_in_22[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_23 = io_in_23[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_24 = io_in_24[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_25 = io_in_25[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_26 = io_in_26[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_27 = io_in_27[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_28 = io_in_28[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_29 = io_in_29[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_30 = io_in_30[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_31 = io_in_31[68]; // @[WallaceTest.scala 105:23]
  wire  c_68_32 = io_in_32[68]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_68_lo_lo = {c_68_7,c_68_6,c_68_5,c_68_4,c_68_3,c_68_2,c_68_1,c_68_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_68_lo = {c_68_15,c_68_14,c_68_13,c_68_12,c_68_11,c_68_10,c_68_9,c_68_8,io_out_68_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_68_hi_lo = {c_68_23,c_68_22,c_68_21,c_68_20,c_68_19,c_68_18,c_68_17,c_68_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_68_hi = {c_68_32,c_68_31,c_68_30,c_68_29,c_68_28,c_68_27,c_68_26,c_68_25,c_68_24,io_out_68_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_69_0 = io_in_0[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_1 = io_in_1[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_2 = io_in_2[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_3 = io_in_3[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_4 = io_in_4[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_5 = io_in_5[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_6 = io_in_6[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_7 = io_in_7[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_8 = io_in_8[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_9 = io_in_9[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_10 = io_in_10[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_11 = io_in_11[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_12 = io_in_12[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_13 = io_in_13[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_14 = io_in_14[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_15 = io_in_15[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_16 = io_in_16[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_17 = io_in_17[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_18 = io_in_18[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_19 = io_in_19[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_20 = io_in_20[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_21 = io_in_21[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_22 = io_in_22[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_23 = io_in_23[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_24 = io_in_24[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_25 = io_in_25[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_26 = io_in_26[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_27 = io_in_27[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_28 = io_in_28[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_29 = io_in_29[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_30 = io_in_30[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_31 = io_in_31[69]; // @[WallaceTest.scala 105:23]
  wire  c_69_32 = io_in_32[69]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_69_lo_lo = {c_69_7,c_69_6,c_69_5,c_69_4,c_69_3,c_69_2,c_69_1,c_69_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_69_lo = {c_69_15,c_69_14,c_69_13,c_69_12,c_69_11,c_69_10,c_69_9,c_69_8,io_out_69_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_69_hi_lo = {c_69_23,c_69_22,c_69_21,c_69_20,c_69_19,c_69_18,c_69_17,c_69_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_69_hi = {c_69_32,c_69_31,c_69_30,c_69_29,c_69_28,c_69_27,c_69_26,c_69_25,c_69_24,io_out_69_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_70_0 = io_in_0[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_1 = io_in_1[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_2 = io_in_2[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_3 = io_in_3[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_4 = io_in_4[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_5 = io_in_5[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_6 = io_in_6[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_7 = io_in_7[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_8 = io_in_8[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_9 = io_in_9[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_10 = io_in_10[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_11 = io_in_11[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_12 = io_in_12[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_13 = io_in_13[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_14 = io_in_14[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_15 = io_in_15[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_16 = io_in_16[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_17 = io_in_17[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_18 = io_in_18[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_19 = io_in_19[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_20 = io_in_20[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_21 = io_in_21[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_22 = io_in_22[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_23 = io_in_23[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_24 = io_in_24[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_25 = io_in_25[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_26 = io_in_26[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_27 = io_in_27[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_28 = io_in_28[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_29 = io_in_29[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_30 = io_in_30[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_31 = io_in_31[70]; // @[WallaceTest.scala 105:23]
  wire  c_70_32 = io_in_32[70]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_70_lo_lo = {c_70_7,c_70_6,c_70_5,c_70_4,c_70_3,c_70_2,c_70_1,c_70_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_70_lo = {c_70_15,c_70_14,c_70_13,c_70_12,c_70_11,c_70_10,c_70_9,c_70_8,io_out_70_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_70_hi_lo = {c_70_23,c_70_22,c_70_21,c_70_20,c_70_19,c_70_18,c_70_17,c_70_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_70_hi = {c_70_32,c_70_31,c_70_30,c_70_29,c_70_28,c_70_27,c_70_26,c_70_25,c_70_24,io_out_70_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_71_0 = io_in_0[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_1 = io_in_1[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_2 = io_in_2[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_3 = io_in_3[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_4 = io_in_4[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_5 = io_in_5[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_6 = io_in_6[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_7 = io_in_7[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_8 = io_in_8[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_9 = io_in_9[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_10 = io_in_10[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_11 = io_in_11[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_12 = io_in_12[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_13 = io_in_13[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_14 = io_in_14[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_15 = io_in_15[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_16 = io_in_16[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_17 = io_in_17[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_18 = io_in_18[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_19 = io_in_19[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_20 = io_in_20[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_21 = io_in_21[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_22 = io_in_22[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_23 = io_in_23[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_24 = io_in_24[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_25 = io_in_25[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_26 = io_in_26[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_27 = io_in_27[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_28 = io_in_28[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_29 = io_in_29[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_30 = io_in_30[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_31 = io_in_31[71]; // @[WallaceTest.scala 105:23]
  wire  c_71_32 = io_in_32[71]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_71_lo_lo = {c_71_7,c_71_6,c_71_5,c_71_4,c_71_3,c_71_2,c_71_1,c_71_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_71_lo = {c_71_15,c_71_14,c_71_13,c_71_12,c_71_11,c_71_10,c_71_9,c_71_8,io_out_71_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_71_hi_lo = {c_71_23,c_71_22,c_71_21,c_71_20,c_71_19,c_71_18,c_71_17,c_71_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_71_hi = {c_71_32,c_71_31,c_71_30,c_71_29,c_71_28,c_71_27,c_71_26,c_71_25,c_71_24,io_out_71_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_72_0 = io_in_0[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_1 = io_in_1[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_2 = io_in_2[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_3 = io_in_3[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_4 = io_in_4[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_5 = io_in_5[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_6 = io_in_6[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_7 = io_in_7[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_8 = io_in_8[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_9 = io_in_9[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_10 = io_in_10[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_11 = io_in_11[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_12 = io_in_12[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_13 = io_in_13[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_14 = io_in_14[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_15 = io_in_15[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_16 = io_in_16[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_17 = io_in_17[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_18 = io_in_18[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_19 = io_in_19[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_20 = io_in_20[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_21 = io_in_21[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_22 = io_in_22[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_23 = io_in_23[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_24 = io_in_24[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_25 = io_in_25[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_26 = io_in_26[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_27 = io_in_27[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_28 = io_in_28[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_29 = io_in_29[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_30 = io_in_30[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_31 = io_in_31[72]; // @[WallaceTest.scala 105:23]
  wire  c_72_32 = io_in_32[72]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_72_lo_lo = {c_72_7,c_72_6,c_72_5,c_72_4,c_72_3,c_72_2,c_72_1,c_72_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_72_lo = {c_72_15,c_72_14,c_72_13,c_72_12,c_72_11,c_72_10,c_72_9,c_72_8,io_out_72_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_72_hi_lo = {c_72_23,c_72_22,c_72_21,c_72_20,c_72_19,c_72_18,c_72_17,c_72_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_72_hi = {c_72_32,c_72_31,c_72_30,c_72_29,c_72_28,c_72_27,c_72_26,c_72_25,c_72_24,io_out_72_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_73_0 = io_in_0[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_1 = io_in_1[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_2 = io_in_2[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_3 = io_in_3[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_4 = io_in_4[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_5 = io_in_5[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_6 = io_in_6[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_7 = io_in_7[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_8 = io_in_8[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_9 = io_in_9[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_10 = io_in_10[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_11 = io_in_11[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_12 = io_in_12[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_13 = io_in_13[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_14 = io_in_14[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_15 = io_in_15[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_16 = io_in_16[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_17 = io_in_17[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_18 = io_in_18[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_19 = io_in_19[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_20 = io_in_20[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_21 = io_in_21[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_22 = io_in_22[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_23 = io_in_23[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_24 = io_in_24[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_25 = io_in_25[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_26 = io_in_26[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_27 = io_in_27[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_28 = io_in_28[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_29 = io_in_29[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_30 = io_in_30[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_31 = io_in_31[73]; // @[WallaceTest.scala 105:23]
  wire  c_73_32 = io_in_32[73]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_73_lo_lo = {c_73_7,c_73_6,c_73_5,c_73_4,c_73_3,c_73_2,c_73_1,c_73_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_73_lo = {c_73_15,c_73_14,c_73_13,c_73_12,c_73_11,c_73_10,c_73_9,c_73_8,io_out_73_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_73_hi_lo = {c_73_23,c_73_22,c_73_21,c_73_20,c_73_19,c_73_18,c_73_17,c_73_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_73_hi = {c_73_32,c_73_31,c_73_30,c_73_29,c_73_28,c_73_27,c_73_26,c_73_25,c_73_24,io_out_73_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_74_0 = io_in_0[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_1 = io_in_1[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_2 = io_in_2[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_3 = io_in_3[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_4 = io_in_4[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_5 = io_in_5[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_6 = io_in_6[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_7 = io_in_7[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_8 = io_in_8[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_9 = io_in_9[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_10 = io_in_10[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_11 = io_in_11[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_12 = io_in_12[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_13 = io_in_13[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_14 = io_in_14[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_15 = io_in_15[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_16 = io_in_16[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_17 = io_in_17[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_18 = io_in_18[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_19 = io_in_19[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_20 = io_in_20[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_21 = io_in_21[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_22 = io_in_22[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_23 = io_in_23[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_24 = io_in_24[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_25 = io_in_25[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_26 = io_in_26[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_27 = io_in_27[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_28 = io_in_28[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_29 = io_in_29[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_30 = io_in_30[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_31 = io_in_31[74]; // @[WallaceTest.scala 105:23]
  wire  c_74_32 = io_in_32[74]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_74_lo_lo = {c_74_7,c_74_6,c_74_5,c_74_4,c_74_3,c_74_2,c_74_1,c_74_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_74_lo = {c_74_15,c_74_14,c_74_13,c_74_12,c_74_11,c_74_10,c_74_9,c_74_8,io_out_74_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_74_hi_lo = {c_74_23,c_74_22,c_74_21,c_74_20,c_74_19,c_74_18,c_74_17,c_74_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_74_hi = {c_74_32,c_74_31,c_74_30,c_74_29,c_74_28,c_74_27,c_74_26,c_74_25,c_74_24,io_out_74_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_75_0 = io_in_0[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_1 = io_in_1[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_2 = io_in_2[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_3 = io_in_3[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_4 = io_in_4[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_5 = io_in_5[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_6 = io_in_6[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_7 = io_in_7[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_8 = io_in_8[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_9 = io_in_9[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_10 = io_in_10[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_11 = io_in_11[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_12 = io_in_12[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_13 = io_in_13[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_14 = io_in_14[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_15 = io_in_15[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_16 = io_in_16[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_17 = io_in_17[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_18 = io_in_18[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_19 = io_in_19[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_20 = io_in_20[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_21 = io_in_21[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_22 = io_in_22[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_23 = io_in_23[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_24 = io_in_24[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_25 = io_in_25[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_26 = io_in_26[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_27 = io_in_27[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_28 = io_in_28[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_29 = io_in_29[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_30 = io_in_30[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_31 = io_in_31[75]; // @[WallaceTest.scala 105:23]
  wire  c_75_32 = io_in_32[75]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_75_lo_lo = {c_75_7,c_75_6,c_75_5,c_75_4,c_75_3,c_75_2,c_75_1,c_75_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_75_lo = {c_75_15,c_75_14,c_75_13,c_75_12,c_75_11,c_75_10,c_75_9,c_75_8,io_out_75_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_75_hi_lo = {c_75_23,c_75_22,c_75_21,c_75_20,c_75_19,c_75_18,c_75_17,c_75_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_75_hi = {c_75_32,c_75_31,c_75_30,c_75_29,c_75_28,c_75_27,c_75_26,c_75_25,c_75_24,io_out_75_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_76_0 = io_in_0[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_1 = io_in_1[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_2 = io_in_2[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_3 = io_in_3[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_4 = io_in_4[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_5 = io_in_5[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_6 = io_in_6[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_7 = io_in_7[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_8 = io_in_8[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_9 = io_in_9[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_10 = io_in_10[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_11 = io_in_11[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_12 = io_in_12[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_13 = io_in_13[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_14 = io_in_14[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_15 = io_in_15[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_16 = io_in_16[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_17 = io_in_17[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_18 = io_in_18[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_19 = io_in_19[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_20 = io_in_20[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_21 = io_in_21[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_22 = io_in_22[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_23 = io_in_23[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_24 = io_in_24[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_25 = io_in_25[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_26 = io_in_26[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_27 = io_in_27[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_28 = io_in_28[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_29 = io_in_29[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_30 = io_in_30[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_31 = io_in_31[76]; // @[WallaceTest.scala 105:23]
  wire  c_76_32 = io_in_32[76]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_76_lo_lo = {c_76_7,c_76_6,c_76_5,c_76_4,c_76_3,c_76_2,c_76_1,c_76_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_76_lo = {c_76_15,c_76_14,c_76_13,c_76_12,c_76_11,c_76_10,c_76_9,c_76_8,io_out_76_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_76_hi_lo = {c_76_23,c_76_22,c_76_21,c_76_20,c_76_19,c_76_18,c_76_17,c_76_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_76_hi = {c_76_32,c_76_31,c_76_30,c_76_29,c_76_28,c_76_27,c_76_26,c_76_25,c_76_24,io_out_76_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_77_0 = io_in_0[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_1 = io_in_1[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_2 = io_in_2[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_3 = io_in_3[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_4 = io_in_4[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_5 = io_in_5[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_6 = io_in_6[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_7 = io_in_7[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_8 = io_in_8[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_9 = io_in_9[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_10 = io_in_10[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_11 = io_in_11[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_12 = io_in_12[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_13 = io_in_13[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_14 = io_in_14[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_15 = io_in_15[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_16 = io_in_16[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_17 = io_in_17[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_18 = io_in_18[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_19 = io_in_19[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_20 = io_in_20[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_21 = io_in_21[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_22 = io_in_22[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_23 = io_in_23[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_24 = io_in_24[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_25 = io_in_25[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_26 = io_in_26[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_27 = io_in_27[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_28 = io_in_28[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_29 = io_in_29[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_30 = io_in_30[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_31 = io_in_31[77]; // @[WallaceTest.scala 105:23]
  wire  c_77_32 = io_in_32[77]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_77_lo_lo = {c_77_7,c_77_6,c_77_5,c_77_4,c_77_3,c_77_2,c_77_1,c_77_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_77_lo = {c_77_15,c_77_14,c_77_13,c_77_12,c_77_11,c_77_10,c_77_9,c_77_8,io_out_77_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_77_hi_lo = {c_77_23,c_77_22,c_77_21,c_77_20,c_77_19,c_77_18,c_77_17,c_77_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_77_hi = {c_77_32,c_77_31,c_77_30,c_77_29,c_77_28,c_77_27,c_77_26,c_77_25,c_77_24,io_out_77_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_78_0 = io_in_0[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_1 = io_in_1[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_2 = io_in_2[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_3 = io_in_3[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_4 = io_in_4[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_5 = io_in_5[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_6 = io_in_6[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_7 = io_in_7[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_8 = io_in_8[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_9 = io_in_9[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_10 = io_in_10[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_11 = io_in_11[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_12 = io_in_12[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_13 = io_in_13[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_14 = io_in_14[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_15 = io_in_15[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_16 = io_in_16[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_17 = io_in_17[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_18 = io_in_18[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_19 = io_in_19[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_20 = io_in_20[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_21 = io_in_21[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_22 = io_in_22[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_23 = io_in_23[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_24 = io_in_24[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_25 = io_in_25[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_26 = io_in_26[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_27 = io_in_27[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_28 = io_in_28[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_29 = io_in_29[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_30 = io_in_30[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_31 = io_in_31[78]; // @[WallaceTest.scala 105:23]
  wire  c_78_32 = io_in_32[78]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_78_lo_lo = {c_78_7,c_78_6,c_78_5,c_78_4,c_78_3,c_78_2,c_78_1,c_78_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_78_lo = {c_78_15,c_78_14,c_78_13,c_78_12,c_78_11,c_78_10,c_78_9,c_78_8,io_out_78_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_78_hi_lo = {c_78_23,c_78_22,c_78_21,c_78_20,c_78_19,c_78_18,c_78_17,c_78_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_78_hi = {c_78_32,c_78_31,c_78_30,c_78_29,c_78_28,c_78_27,c_78_26,c_78_25,c_78_24,io_out_78_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_79_0 = io_in_0[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_1 = io_in_1[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_2 = io_in_2[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_3 = io_in_3[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_4 = io_in_4[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_5 = io_in_5[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_6 = io_in_6[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_7 = io_in_7[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_8 = io_in_8[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_9 = io_in_9[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_10 = io_in_10[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_11 = io_in_11[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_12 = io_in_12[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_13 = io_in_13[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_14 = io_in_14[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_15 = io_in_15[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_16 = io_in_16[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_17 = io_in_17[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_18 = io_in_18[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_19 = io_in_19[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_20 = io_in_20[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_21 = io_in_21[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_22 = io_in_22[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_23 = io_in_23[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_24 = io_in_24[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_25 = io_in_25[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_26 = io_in_26[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_27 = io_in_27[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_28 = io_in_28[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_29 = io_in_29[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_30 = io_in_30[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_31 = io_in_31[79]; // @[WallaceTest.scala 105:23]
  wire  c_79_32 = io_in_32[79]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_79_lo_lo = {c_79_7,c_79_6,c_79_5,c_79_4,c_79_3,c_79_2,c_79_1,c_79_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_79_lo = {c_79_15,c_79_14,c_79_13,c_79_12,c_79_11,c_79_10,c_79_9,c_79_8,io_out_79_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_79_hi_lo = {c_79_23,c_79_22,c_79_21,c_79_20,c_79_19,c_79_18,c_79_17,c_79_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_79_hi = {c_79_32,c_79_31,c_79_30,c_79_29,c_79_28,c_79_27,c_79_26,c_79_25,c_79_24,io_out_79_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_80_0 = io_in_0[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_1 = io_in_1[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_2 = io_in_2[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_3 = io_in_3[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_4 = io_in_4[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_5 = io_in_5[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_6 = io_in_6[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_7 = io_in_7[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_8 = io_in_8[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_9 = io_in_9[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_10 = io_in_10[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_11 = io_in_11[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_12 = io_in_12[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_13 = io_in_13[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_14 = io_in_14[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_15 = io_in_15[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_16 = io_in_16[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_17 = io_in_17[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_18 = io_in_18[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_19 = io_in_19[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_20 = io_in_20[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_21 = io_in_21[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_22 = io_in_22[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_23 = io_in_23[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_24 = io_in_24[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_25 = io_in_25[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_26 = io_in_26[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_27 = io_in_27[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_28 = io_in_28[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_29 = io_in_29[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_30 = io_in_30[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_31 = io_in_31[80]; // @[WallaceTest.scala 105:23]
  wire  c_80_32 = io_in_32[80]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_80_lo_lo = {c_80_7,c_80_6,c_80_5,c_80_4,c_80_3,c_80_2,c_80_1,c_80_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_80_lo = {c_80_15,c_80_14,c_80_13,c_80_12,c_80_11,c_80_10,c_80_9,c_80_8,io_out_80_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_80_hi_lo = {c_80_23,c_80_22,c_80_21,c_80_20,c_80_19,c_80_18,c_80_17,c_80_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_80_hi = {c_80_32,c_80_31,c_80_30,c_80_29,c_80_28,c_80_27,c_80_26,c_80_25,c_80_24,io_out_80_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_81_0 = io_in_0[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_1 = io_in_1[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_2 = io_in_2[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_3 = io_in_3[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_4 = io_in_4[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_5 = io_in_5[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_6 = io_in_6[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_7 = io_in_7[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_8 = io_in_8[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_9 = io_in_9[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_10 = io_in_10[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_11 = io_in_11[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_12 = io_in_12[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_13 = io_in_13[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_14 = io_in_14[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_15 = io_in_15[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_16 = io_in_16[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_17 = io_in_17[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_18 = io_in_18[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_19 = io_in_19[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_20 = io_in_20[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_21 = io_in_21[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_22 = io_in_22[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_23 = io_in_23[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_24 = io_in_24[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_25 = io_in_25[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_26 = io_in_26[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_27 = io_in_27[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_28 = io_in_28[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_29 = io_in_29[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_30 = io_in_30[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_31 = io_in_31[81]; // @[WallaceTest.scala 105:23]
  wire  c_81_32 = io_in_32[81]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_81_lo_lo = {c_81_7,c_81_6,c_81_5,c_81_4,c_81_3,c_81_2,c_81_1,c_81_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_81_lo = {c_81_15,c_81_14,c_81_13,c_81_12,c_81_11,c_81_10,c_81_9,c_81_8,io_out_81_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_81_hi_lo = {c_81_23,c_81_22,c_81_21,c_81_20,c_81_19,c_81_18,c_81_17,c_81_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_81_hi = {c_81_32,c_81_31,c_81_30,c_81_29,c_81_28,c_81_27,c_81_26,c_81_25,c_81_24,io_out_81_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_82_0 = io_in_0[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_1 = io_in_1[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_2 = io_in_2[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_3 = io_in_3[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_4 = io_in_4[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_5 = io_in_5[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_6 = io_in_6[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_7 = io_in_7[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_8 = io_in_8[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_9 = io_in_9[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_10 = io_in_10[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_11 = io_in_11[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_12 = io_in_12[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_13 = io_in_13[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_14 = io_in_14[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_15 = io_in_15[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_16 = io_in_16[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_17 = io_in_17[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_18 = io_in_18[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_19 = io_in_19[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_20 = io_in_20[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_21 = io_in_21[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_22 = io_in_22[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_23 = io_in_23[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_24 = io_in_24[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_25 = io_in_25[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_26 = io_in_26[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_27 = io_in_27[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_28 = io_in_28[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_29 = io_in_29[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_30 = io_in_30[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_31 = io_in_31[82]; // @[WallaceTest.scala 105:23]
  wire  c_82_32 = io_in_32[82]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_82_lo_lo = {c_82_7,c_82_6,c_82_5,c_82_4,c_82_3,c_82_2,c_82_1,c_82_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_82_lo = {c_82_15,c_82_14,c_82_13,c_82_12,c_82_11,c_82_10,c_82_9,c_82_8,io_out_82_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_82_hi_lo = {c_82_23,c_82_22,c_82_21,c_82_20,c_82_19,c_82_18,c_82_17,c_82_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_82_hi = {c_82_32,c_82_31,c_82_30,c_82_29,c_82_28,c_82_27,c_82_26,c_82_25,c_82_24,io_out_82_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_83_0 = io_in_0[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_1 = io_in_1[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_2 = io_in_2[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_3 = io_in_3[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_4 = io_in_4[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_5 = io_in_5[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_6 = io_in_6[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_7 = io_in_7[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_8 = io_in_8[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_9 = io_in_9[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_10 = io_in_10[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_11 = io_in_11[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_12 = io_in_12[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_13 = io_in_13[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_14 = io_in_14[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_15 = io_in_15[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_16 = io_in_16[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_17 = io_in_17[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_18 = io_in_18[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_19 = io_in_19[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_20 = io_in_20[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_21 = io_in_21[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_22 = io_in_22[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_23 = io_in_23[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_24 = io_in_24[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_25 = io_in_25[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_26 = io_in_26[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_27 = io_in_27[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_28 = io_in_28[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_29 = io_in_29[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_30 = io_in_30[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_31 = io_in_31[83]; // @[WallaceTest.scala 105:23]
  wire  c_83_32 = io_in_32[83]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_83_lo_lo = {c_83_7,c_83_6,c_83_5,c_83_4,c_83_3,c_83_2,c_83_1,c_83_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_83_lo = {c_83_15,c_83_14,c_83_13,c_83_12,c_83_11,c_83_10,c_83_9,c_83_8,io_out_83_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_83_hi_lo = {c_83_23,c_83_22,c_83_21,c_83_20,c_83_19,c_83_18,c_83_17,c_83_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_83_hi = {c_83_32,c_83_31,c_83_30,c_83_29,c_83_28,c_83_27,c_83_26,c_83_25,c_83_24,io_out_83_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_84_0 = io_in_0[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_1 = io_in_1[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_2 = io_in_2[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_3 = io_in_3[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_4 = io_in_4[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_5 = io_in_5[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_6 = io_in_6[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_7 = io_in_7[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_8 = io_in_8[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_9 = io_in_9[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_10 = io_in_10[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_11 = io_in_11[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_12 = io_in_12[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_13 = io_in_13[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_14 = io_in_14[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_15 = io_in_15[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_16 = io_in_16[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_17 = io_in_17[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_18 = io_in_18[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_19 = io_in_19[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_20 = io_in_20[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_21 = io_in_21[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_22 = io_in_22[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_23 = io_in_23[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_24 = io_in_24[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_25 = io_in_25[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_26 = io_in_26[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_27 = io_in_27[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_28 = io_in_28[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_29 = io_in_29[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_30 = io_in_30[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_31 = io_in_31[84]; // @[WallaceTest.scala 105:23]
  wire  c_84_32 = io_in_32[84]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_84_lo_lo = {c_84_7,c_84_6,c_84_5,c_84_4,c_84_3,c_84_2,c_84_1,c_84_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_84_lo = {c_84_15,c_84_14,c_84_13,c_84_12,c_84_11,c_84_10,c_84_9,c_84_8,io_out_84_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_84_hi_lo = {c_84_23,c_84_22,c_84_21,c_84_20,c_84_19,c_84_18,c_84_17,c_84_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_84_hi = {c_84_32,c_84_31,c_84_30,c_84_29,c_84_28,c_84_27,c_84_26,c_84_25,c_84_24,io_out_84_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_85_0 = io_in_0[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_1 = io_in_1[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_2 = io_in_2[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_3 = io_in_3[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_4 = io_in_4[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_5 = io_in_5[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_6 = io_in_6[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_7 = io_in_7[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_8 = io_in_8[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_9 = io_in_9[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_10 = io_in_10[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_11 = io_in_11[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_12 = io_in_12[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_13 = io_in_13[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_14 = io_in_14[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_15 = io_in_15[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_16 = io_in_16[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_17 = io_in_17[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_18 = io_in_18[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_19 = io_in_19[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_20 = io_in_20[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_21 = io_in_21[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_22 = io_in_22[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_23 = io_in_23[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_24 = io_in_24[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_25 = io_in_25[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_26 = io_in_26[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_27 = io_in_27[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_28 = io_in_28[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_29 = io_in_29[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_30 = io_in_30[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_31 = io_in_31[85]; // @[WallaceTest.scala 105:23]
  wire  c_85_32 = io_in_32[85]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_85_lo_lo = {c_85_7,c_85_6,c_85_5,c_85_4,c_85_3,c_85_2,c_85_1,c_85_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_85_lo = {c_85_15,c_85_14,c_85_13,c_85_12,c_85_11,c_85_10,c_85_9,c_85_8,io_out_85_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_85_hi_lo = {c_85_23,c_85_22,c_85_21,c_85_20,c_85_19,c_85_18,c_85_17,c_85_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_85_hi = {c_85_32,c_85_31,c_85_30,c_85_29,c_85_28,c_85_27,c_85_26,c_85_25,c_85_24,io_out_85_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_86_0 = io_in_0[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_1 = io_in_1[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_2 = io_in_2[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_3 = io_in_3[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_4 = io_in_4[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_5 = io_in_5[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_6 = io_in_6[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_7 = io_in_7[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_8 = io_in_8[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_9 = io_in_9[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_10 = io_in_10[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_11 = io_in_11[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_12 = io_in_12[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_13 = io_in_13[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_14 = io_in_14[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_15 = io_in_15[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_16 = io_in_16[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_17 = io_in_17[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_18 = io_in_18[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_19 = io_in_19[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_20 = io_in_20[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_21 = io_in_21[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_22 = io_in_22[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_23 = io_in_23[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_24 = io_in_24[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_25 = io_in_25[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_26 = io_in_26[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_27 = io_in_27[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_28 = io_in_28[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_29 = io_in_29[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_30 = io_in_30[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_31 = io_in_31[86]; // @[WallaceTest.scala 105:23]
  wire  c_86_32 = io_in_32[86]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_86_lo_lo = {c_86_7,c_86_6,c_86_5,c_86_4,c_86_3,c_86_2,c_86_1,c_86_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_86_lo = {c_86_15,c_86_14,c_86_13,c_86_12,c_86_11,c_86_10,c_86_9,c_86_8,io_out_86_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_86_hi_lo = {c_86_23,c_86_22,c_86_21,c_86_20,c_86_19,c_86_18,c_86_17,c_86_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_86_hi = {c_86_32,c_86_31,c_86_30,c_86_29,c_86_28,c_86_27,c_86_26,c_86_25,c_86_24,io_out_86_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_87_0 = io_in_0[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_1 = io_in_1[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_2 = io_in_2[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_3 = io_in_3[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_4 = io_in_4[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_5 = io_in_5[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_6 = io_in_6[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_7 = io_in_7[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_8 = io_in_8[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_9 = io_in_9[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_10 = io_in_10[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_11 = io_in_11[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_12 = io_in_12[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_13 = io_in_13[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_14 = io_in_14[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_15 = io_in_15[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_16 = io_in_16[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_17 = io_in_17[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_18 = io_in_18[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_19 = io_in_19[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_20 = io_in_20[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_21 = io_in_21[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_22 = io_in_22[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_23 = io_in_23[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_24 = io_in_24[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_25 = io_in_25[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_26 = io_in_26[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_27 = io_in_27[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_28 = io_in_28[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_29 = io_in_29[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_30 = io_in_30[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_31 = io_in_31[87]; // @[WallaceTest.scala 105:23]
  wire  c_87_32 = io_in_32[87]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_87_lo_lo = {c_87_7,c_87_6,c_87_5,c_87_4,c_87_3,c_87_2,c_87_1,c_87_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_87_lo = {c_87_15,c_87_14,c_87_13,c_87_12,c_87_11,c_87_10,c_87_9,c_87_8,io_out_87_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_87_hi_lo = {c_87_23,c_87_22,c_87_21,c_87_20,c_87_19,c_87_18,c_87_17,c_87_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_87_hi = {c_87_32,c_87_31,c_87_30,c_87_29,c_87_28,c_87_27,c_87_26,c_87_25,c_87_24,io_out_87_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_88_0 = io_in_0[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_1 = io_in_1[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_2 = io_in_2[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_3 = io_in_3[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_4 = io_in_4[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_5 = io_in_5[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_6 = io_in_6[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_7 = io_in_7[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_8 = io_in_8[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_9 = io_in_9[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_10 = io_in_10[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_11 = io_in_11[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_12 = io_in_12[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_13 = io_in_13[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_14 = io_in_14[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_15 = io_in_15[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_16 = io_in_16[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_17 = io_in_17[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_18 = io_in_18[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_19 = io_in_19[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_20 = io_in_20[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_21 = io_in_21[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_22 = io_in_22[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_23 = io_in_23[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_24 = io_in_24[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_25 = io_in_25[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_26 = io_in_26[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_27 = io_in_27[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_28 = io_in_28[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_29 = io_in_29[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_30 = io_in_30[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_31 = io_in_31[88]; // @[WallaceTest.scala 105:23]
  wire  c_88_32 = io_in_32[88]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_88_lo_lo = {c_88_7,c_88_6,c_88_5,c_88_4,c_88_3,c_88_2,c_88_1,c_88_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_88_lo = {c_88_15,c_88_14,c_88_13,c_88_12,c_88_11,c_88_10,c_88_9,c_88_8,io_out_88_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_88_hi_lo = {c_88_23,c_88_22,c_88_21,c_88_20,c_88_19,c_88_18,c_88_17,c_88_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_88_hi = {c_88_32,c_88_31,c_88_30,c_88_29,c_88_28,c_88_27,c_88_26,c_88_25,c_88_24,io_out_88_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_89_0 = io_in_0[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_1 = io_in_1[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_2 = io_in_2[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_3 = io_in_3[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_4 = io_in_4[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_5 = io_in_5[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_6 = io_in_6[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_7 = io_in_7[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_8 = io_in_8[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_9 = io_in_9[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_10 = io_in_10[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_11 = io_in_11[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_12 = io_in_12[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_13 = io_in_13[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_14 = io_in_14[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_15 = io_in_15[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_16 = io_in_16[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_17 = io_in_17[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_18 = io_in_18[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_19 = io_in_19[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_20 = io_in_20[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_21 = io_in_21[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_22 = io_in_22[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_23 = io_in_23[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_24 = io_in_24[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_25 = io_in_25[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_26 = io_in_26[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_27 = io_in_27[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_28 = io_in_28[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_29 = io_in_29[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_30 = io_in_30[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_31 = io_in_31[89]; // @[WallaceTest.scala 105:23]
  wire  c_89_32 = io_in_32[89]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_89_lo_lo = {c_89_7,c_89_6,c_89_5,c_89_4,c_89_3,c_89_2,c_89_1,c_89_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_89_lo = {c_89_15,c_89_14,c_89_13,c_89_12,c_89_11,c_89_10,c_89_9,c_89_8,io_out_89_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_89_hi_lo = {c_89_23,c_89_22,c_89_21,c_89_20,c_89_19,c_89_18,c_89_17,c_89_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_89_hi = {c_89_32,c_89_31,c_89_30,c_89_29,c_89_28,c_89_27,c_89_26,c_89_25,c_89_24,io_out_89_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_90_0 = io_in_0[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_1 = io_in_1[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_2 = io_in_2[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_3 = io_in_3[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_4 = io_in_4[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_5 = io_in_5[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_6 = io_in_6[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_7 = io_in_7[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_8 = io_in_8[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_9 = io_in_9[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_10 = io_in_10[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_11 = io_in_11[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_12 = io_in_12[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_13 = io_in_13[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_14 = io_in_14[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_15 = io_in_15[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_16 = io_in_16[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_17 = io_in_17[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_18 = io_in_18[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_19 = io_in_19[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_20 = io_in_20[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_21 = io_in_21[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_22 = io_in_22[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_23 = io_in_23[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_24 = io_in_24[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_25 = io_in_25[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_26 = io_in_26[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_27 = io_in_27[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_28 = io_in_28[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_29 = io_in_29[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_30 = io_in_30[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_31 = io_in_31[90]; // @[WallaceTest.scala 105:23]
  wire  c_90_32 = io_in_32[90]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_90_lo_lo = {c_90_7,c_90_6,c_90_5,c_90_4,c_90_3,c_90_2,c_90_1,c_90_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_90_lo = {c_90_15,c_90_14,c_90_13,c_90_12,c_90_11,c_90_10,c_90_9,c_90_8,io_out_90_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_90_hi_lo = {c_90_23,c_90_22,c_90_21,c_90_20,c_90_19,c_90_18,c_90_17,c_90_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_90_hi = {c_90_32,c_90_31,c_90_30,c_90_29,c_90_28,c_90_27,c_90_26,c_90_25,c_90_24,io_out_90_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_91_0 = io_in_0[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_1 = io_in_1[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_2 = io_in_2[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_3 = io_in_3[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_4 = io_in_4[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_5 = io_in_5[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_6 = io_in_6[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_7 = io_in_7[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_8 = io_in_8[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_9 = io_in_9[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_10 = io_in_10[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_11 = io_in_11[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_12 = io_in_12[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_13 = io_in_13[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_14 = io_in_14[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_15 = io_in_15[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_16 = io_in_16[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_17 = io_in_17[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_18 = io_in_18[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_19 = io_in_19[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_20 = io_in_20[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_21 = io_in_21[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_22 = io_in_22[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_23 = io_in_23[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_24 = io_in_24[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_25 = io_in_25[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_26 = io_in_26[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_27 = io_in_27[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_28 = io_in_28[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_29 = io_in_29[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_30 = io_in_30[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_31 = io_in_31[91]; // @[WallaceTest.scala 105:23]
  wire  c_91_32 = io_in_32[91]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_91_lo_lo = {c_91_7,c_91_6,c_91_5,c_91_4,c_91_3,c_91_2,c_91_1,c_91_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_91_lo = {c_91_15,c_91_14,c_91_13,c_91_12,c_91_11,c_91_10,c_91_9,c_91_8,io_out_91_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_91_hi_lo = {c_91_23,c_91_22,c_91_21,c_91_20,c_91_19,c_91_18,c_91_17,c_91_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_91_hi = {c_91_32,c_91_31,c_91_30,c_91_29,c_91_28,c_91_27,c_91_26,c_91_25,c_91_24,io_out_91_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_92_0 = io_in_0[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_1 = io_in_1[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_2 = io_in_2[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_3 = io_in_3[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_4 = io_in_4[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_5 = io_in_5[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_6 = io_in_6[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_7 = io_in_7[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_8 = io_in_8[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_9 = io_in_9[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_10 = io_in_10[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_11 = io_in_11[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_12 = io_in_12[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_13 = io_in_13[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_14 = io_in_14[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_15 = io_in_15[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_16 = io_in_16[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_17 = io_in_17[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_18 = io_in_18[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_19 = io_in_19[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_20 = io_in_20[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_21 = io_in_21[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_22 = io_in_22[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_23 = io_in_23[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_24 = io_in_24[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_25 = io_in_25[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_26 = io_in_26[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_27 = io_in_27[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_28 = io_in_28[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_29 = io_in_29[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_30 = io_in_30[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_31 = io_in_31[92]; // @[WallaceTest.scala 105:23]
  wire  c_92_32 = io_in_32[92]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_92_lo_lo = {c_92_7,c_92_6,c_92_5,c_92_4,c_92_3,c_92_2,c_92_1,c_92_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_92_lo = {c_92_15,c_92_14,c_92_13,c_92_12,c_92_11,c_92_10,c_92_9,c_92_8,io_out_92_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_92_hi_lo = {c_92_23,c_92_22,c_92_21,c_92_20,c_92_19,c_92_18,c_92_17,c_92_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_92_hi = {c_92_32,c_92_31,c_92_30,c_92_29,c_92_28,c_92_27,c_92_26,c_92_25,c_92_24,io_out_92_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_93_0 = io_in_0[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_1 = io_in_1[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_2 = io_in_2[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_3 = io_in_3[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_4 = io_in_4[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_5 = io_in_5[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_6 = io_in_6[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_7 = io_in_7[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_8 = io_in_8[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_9 = io_in_9[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_10 = io_in_10[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_11 = io_in_11[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_12 = io_in_12[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_13 = io_in_13[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_14 = io_in_14[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_15 = io_in_15[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_16 = io_in_16[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_17 = io_in_17[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_18 = io_in_18[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_19 = io_in_19[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_20 = io_in_20[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_21 = io_in_21[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_22 = io_in_22[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_23 = io_in_23[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_24 = io_in_24[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_25 = io_in_25[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_26 = io_in_26[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_27 = io_in_27[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_28 = io_in_28[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_29 = io_in_29[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_30 = io_in_30[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_31 = io_in_31[93]; // @[WallaceTest.scala 105:23]
  wire  c_93_32 = io_in_32[93]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_93_lo_lo = {c_93_7,c_93_6,c_93_5,c_93_4,c_93_3,c_93_2,c_93_1,c_93_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_93_lo = {c_93_15,c_93_14,c_93_13,c_93_12,c_93_11,c_93_10,c_93_9,c_93_8,io_out_93_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_93_hi_lo = {c_93_23,c_93_22,c_93_21,c_93_20,c_93_19,c_93_18,c_93_17,c_93_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_93_hi = {c_93_32,c_93_31,c_93_30,c_93_29,c_93_28,c_93_27,c_93_26,c_93_25,c_93_24,io_out_93_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_94_0 = io_in_0[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_1 = io_in_1[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_2 = io_in_2[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_3 = io_in_3[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_4 = io_in_4[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_5 = io_in_5[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_6 = io_in_6[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_7 = io_in_7[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_8 = io_in_8[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_9 = io_in_9[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_10 = io_in_10[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_11 = io_in_11[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_12 = io_in_12[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_13 = io_in_13[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_14 = io_in_14[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_15 = io_in_15[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_16 = io_in_16[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_17 = io_in_17[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_18 = io_in_18[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_19 = io_in_19[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_20 = io_in_20[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_21 = io_in_21[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_22 = io_in_22[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_23 = io_in_23[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_24 = io_in_24[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_25 = io_in_25[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_26 = io_in_26[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_27 = io_in_27[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_28 = io_in_28[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_29 = io_in_29[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_30 = io_in_30[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_31 = io_in_31[94]; // @[WallaceTest.scala 105:23]
  wire  c_94_32 = io_in_32[94]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_94_lo_lo = {c_94_7,c_94_6,c_94_5,c_94_4,c_94_3,c_94_2,c_94_1,c_94_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_94_lo = {c_94_15,c_94_14,c_94_13,c_94_12,c_94_11,c_94_10,c_94_9,c_94_8,io_out_94_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_94_hi_lo = {c_94_23,c_94_22,c_94_21,c_94_20,c_94_19,c_94_18,c_94_17,c_94_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_94_hi = {c_94_32,c_94_31,c_94_30,c_94_29,c_94_28,c_94_27,c_94_26,c_94_25,c_94_24,io_out_94_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_95_0 = io_in_0[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_1 = io_in_1[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_2 = io_in_2[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_3 = io_in_3[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_4 = io_in_4[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_5 = io_in_5[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_6 = io_in_6[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_7 = io_in_7[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_8 = io_in_8[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_9 = io_in_9[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_10 = io_in_10[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_11 = io_in_11[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_12 = io_in_12[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_13 = io_in_13[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_14 = io_in_14[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_15 = io_in_15[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_16 = io_in_16[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_17 = io_in_17[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_18 = io_in_18[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_19 = io_in_19[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_20 = io_in_20[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_21 = io_in_21[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_22 = io_in_22[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_23 = io_in_23[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_24 = io_in_24[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_25 = io_in_25[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_26 = io_in_26[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_27 = io_in_27[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_28 = io_in_28[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_29 = io_in_29[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_30 = io_in_30[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_31 = io_in_31[95]; // @[WallaceTest.scala 105:23]
  wire  c_95_32 = io_in_32[95]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_95_lo_lo = {c_95_7,c_95_6,c_95_5,c_95_4,c_95_3,c_95_2,c_95_1,c_95_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_95_lo = {c_95_15,c_95_14,c_95_13,c_95_12,c_95_11,c_95_10,c_95_9,c_95_8,io_out_95_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_95_hi_lo = {c_95_23,c_95_22,c_95_21,c_95_20,c_95_19,c_95_18,c_95_17,c_95_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_95_hi = {c_95_32,c_95_31,c_95_30,c_95_29,c_95_28,c_95_27,c_95_26,c_95_25,c_95_24,io_out_95_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_96_0 = io_in_0[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_1 = io_in_1[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_2 = io_in_2[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_3 = io_in_3[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_4 = io_in_4[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_5 = io_in_5[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_6 = io_in_6[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_7 = io_in_7[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_8 = io_in_8[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_9 = io_in_9[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_10 = io_in_10[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_11 = io_in_11[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_12 = io_in_12[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_13 = io_in_13[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_14 = io_in_14[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_15 = io_in_15[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_16 = io_in_16[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_17 = io_in_17[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_18 = io_in_18[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_19 = io_in_19[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_20 = io_in_20[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_21 = io_in_21[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_22 = io_in_22[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_23 = io_in_23[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_24 = io_in_24[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_25 = io_in_25[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_26 = io_in_26[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_27 = io_in_27[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_28 = io_in_28[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_29 = io_in_29[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_30 = io_in_30[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_31 = io_in_31[96]; // @[WallaceTest.scala 105:23]
  wire  c_96_32 = io_in_32[96]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_96_lo_lo = {c_96_7,c_96_6,c_96_5,c_96_4,c_96_3,c_96_2,c_96_1,c_96_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_96_lo = {c_96_15,c_96_14,c_96_13,c_96_12,c_96_11,c_96_10,c_96_9,c_96_8,io_out_96_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_96_hi_lo = {c_96_23,c_96_22,c_96_21,c_96_20,c_96_19,c_96_18,c_96_17,c_96_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_96_hi = {c_96_32,c_96_31,c_96_30,c_96_29,c_96_28,c_96_27,c_96_26,c_96_25,c_96_24,io_out_96_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_97_0 = io_in_0[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_1 = io_in_1[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_2 = io_in_2[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_3 = io_in_3[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_4 = io_in_4[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_5 = io_in_5[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_6 = io_in_6[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_7 = io_in_7[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_8 = io_in_8[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_9 = io_in_9[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_10 = io_in_10[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_11 = io_in_11[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_12 = io_in_12[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_13 = io_in_13[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_14 = io_in_14[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_15 = io_in_15[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_16 = io_in_16[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_17 = io_in_17[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_18 = io_in_18[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_19 = io_in_19[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_20 = io_in_20[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_21 = io_in_21[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_22 = io_in_22[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_23 = io_in_23[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_24 = io_in_24[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_25 = io_in_25[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_26 = io_in_26[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_27 = io_in_27[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_28 = io_in_28[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_29 = io_in_29[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_30 = io_in_30[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_31 = io_in_31[97]; // @[WallaceTest.scala 105:23]
  wire  c_97_32 = io_in_32[97]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_97_lo_lo = {c_97_7,c_97_6,c_97_5,c_97_4,c_97_3,c_97_2,c_97_1,c_97_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_97_lo = {c_97_15,c_97_14,c_97_13,c_97_12,c_97_11,c_97_10,c_97_9,c_97_8,io_out_97_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_97_hi_lo = {c_97_23,c_97_22,c_97_21,c_97_20,c_97_19,c_97_18,c_97_17,c_97_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_97_hi = {c_97_32,c_97_31,c_97_30,c_97_29,c_97_28,c_97_27,c_97_26,c_97_25,c_97_24,io_out_97_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_98_0 = io_in_0[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_1 = io_in_1[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_2 = io_in_2[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_3 = io_in_3[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_4 = io_in_4[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_5 = io_in_5[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_6 = io_in_6[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_7 = io_in_7[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_8 = io_in_8[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_9 = io_in_9[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_10 = io_in_10[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_11 = io_in_11[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_12 = io_in_12[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_13 = io_in_13[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_14 = io_in_14[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_15 = io_in_15[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_16 = io_in_16[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_17 = io_in_17[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_18 = io_in_18[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_19 = io_in_19[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_20 = io_in_20[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_21 = io_in_21[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_22 = io_in_22[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_23 = io_in_23[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_24 = io_in_24[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_25 = io_in_25[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_26 = io_in_26[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_27 = io_in_27[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_28 = io_in_28[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_29 = io_in_29[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_30 = io_in_30[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_31 = io_in_31[98]; // @[WallaceTest.scala 105:23]
  wire  c_98_32 = io_in_32[98]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_98_lo_lo = {c_98_7,c_98_6,c_98_5,c_98_4,c_98_3,c_98_2,c_98_1,c_98_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_98_lo = {c_98_15,c_98_14,c_98_13,c_98_12,c_98_11,c_98_10,c_98_9,c_98_8,io_out_98_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_98_hi_lo = {c_98_23,c_98_22,c_98_21,c_98_20,c_98_19,c_98_18,c_98_17,c_98_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_98_hi = {c_98_32,c_98_31,c_98_30,c_98_29,c_98_28,c_98_27,c_98_26,c_98_25,c_98_24,io_out_98_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_99_0 = io_in_0[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_1 = io_in_1[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_2 = io_in_2[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_3 = io_in_3[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_4 = io_in_4[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_5 = io_in_5[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_6 = io_in_6[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_7 = io_in_7[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_8 = io_in_8[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_9 = io_in_9[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_10 = io_in_10[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_11 = io_in_11[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_12 = io_in_12[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_13 = io_in_13[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_14 = io_in_14[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_15 = io_in_15[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_16 = io_in_16[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_17 = io_in_17[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_18 = io_in_18[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_19 = io_in_19[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_20 = io_in_20[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_21 = io_in_21[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_22 = io_in_22[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_23 = io_in_23[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_24 = io_in_24[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_25 = io_in_25[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_26 = io_in_26[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_27 = io_in_27[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_28 = io_in_28[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_29 = io_in_29[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_30 = io_in_30[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_31 = io_in_31[99]; // @[WallaceTest.scala 105:23]
  wire  c_99_32 = io_in_32[99]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_99_lo_lo = {c_99_7,c_99_6,c_99_5,c_99_4,c_99_3,c_99_2,c_99_1,c_99_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_99_lo = {c_99_15,c_99_14,c_99_13,c_99_12,c_99_11,c_99_10,c_99_9,c_99_8,io_out_99_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_99_hi_lo = {c_99_23,c_99_22,c_99_21,c_99_20,c_99_19,c_99_18,c_99_17,c_99_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_99_hi = {c_99_32,c_99_31,c_99_30,c_99_29,c_99_28,c_99_27,c_99_26,c_99_25,c_99_24,io_out_99_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_100_0 = io_in_0[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_1 = io_in_1[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_2 = io_in_2[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_3 = io_in_3[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_4 = io_in_4[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_5 = io_in_5[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_6 = io_in_6[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_7 = io_in_7[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_8 = io_in_8[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_9 = io_in_9[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_10 = io_in_10[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_11 = io_in_11[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_12 = io_in_12[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_13 = io_in_13[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_14 = io_in_14[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_15 = io_in_15[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_16 = io_in_16[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_17 = io_in_17[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_18 = io_in_18[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_19 = io_in_19[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_20 = io_in_20[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_21 = io_in_21[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_22 = io_in_22[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_23 = io_in_23[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_24 = io_in_24[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_25 = io_in_25[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_26 = io_in_26[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_27 = io_in_27[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_28 = io_in_28[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_29 = io_in_29[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_30 = io_in_30[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_31 = io_in_31[100]; // @[WallaceTest.scala 105:23]
  wire  c_100_32 = io_in_32[100]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_100_lo_lo = {c_100_7,c_100_6,c_100_5,c_100_4,c_100_3,c_100_2,c_100_1,c_100_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_100_lo = {c_100_15,c_100_14,c_100_13,c_100_12,c_100_11,c_100_10,c_100_9,c_100_8,io_out_100_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_100_hi_lo = {c_100_23,c_100_22,c_100_21,c_100_20,c_100_19,c_100_18,c_100_17,c_100_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_100_hi = {c_100_32,c_100_31,c_100_30,c_100_29,c_100_28,c_100_27,c_100_26,c_100_25,c_100_24,
    io_out_100_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_101_0 = io_in_0[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_1 = io_in_1[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_2 = io_in_2[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_3 = io_in_3[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_4 = io_in_4[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_5 = io_in_5[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_6 = io_in_6[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_7 = io_in_7[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_8 = io_in_8[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_9 = io_in_9[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_10 = io_in_10[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_11 = io_in_11[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_12 = io_in_12[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_13 = io_in_13[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_14 = io_in_14[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_15 = io_in_15[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_16 = io_in_16[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_17 = io_in_17[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_18 = io_in_18[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_19 = io_in_19[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_20 = io_in_20[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_21 = io_in_21[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_22 = io_in_22[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_23 = io_in_23[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_24 = io_in_24[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_25 = io_in_25[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_26 = io_in_26[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_27 = io_in_27[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_28 = io_in_28[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_29 = io_in_29[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_30 = io_in_30[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_31 = io_in_31[101]; // @[WallaceTest.scala 105:23]
  wire  c_101_32 = io_in_32[101]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_101_lo_lo = {c_101_7,c_101_6,c_101_5,c_101_4,c_101_3,c_101_2,c_101_1,c_101_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_101_lo = {c_101_15,c_101_14,c_101_13,c_101_12,c_101_11,c_101_10,c_101_9,c_101_8,io_out_101_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_101_hi_lo = {c_101_23,c_101_22,c_101_21,c_101_20,c_101_19,c_101_18,c_101_17,c_101_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_101_hi = {c_101_32,c_101_31,c_101_30,c_101_29,c_101_28,c_101_27,c_101_26,c_101_25,c_101_24,
    io_out_101_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_102_0 = io_in_0[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_1 = io_in_1[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_2 = io_in_2[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_3 = io_in_3[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_4 = io_in_4[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_5 = io_in_5[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_6 = io_in_6[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_7 = io_in_7[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_8 = io_in_8[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_9 = io_in_9[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_10 = io_in_10[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_11 = io_in_11[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_12 = io_in_12[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_13 = io_in_13[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_14 = io_in_14[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_15 = io_in_15[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_16 = io_in_16[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_17 = io_in_17[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_18 = io_in_18[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_19 = io_in_19[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_20 = io_in_20[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_21 = io_in_21[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_22 = io_in_22[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_23 = io_in_23[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_24 = io_in_24[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_25 = io_in_25[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_26 = io_in_26[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_27 = io_in_27[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_28 = io_in_28[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_29 = io_in_29[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_30 = io_in_30[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_31 = io_in_31[102]; // @[WallaceTest.scala 105:23]
  wire  c_102_32 = io_in_32[102]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_102_lo_lo = {c_102_7,c_102_6,c_102_5,c_102_4,c_102_3,c_102_2,c_102_1,c_102_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_102_lo = {c_102_15,c_102_14,c_102_13,c_102_12,c_102_11,c_102_10,c_102_9,c_102_8,io_out_102_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_102_hi_lo = {c_102_23,c_102_22,c_102_21,c_102_20,c_102_19,c_102_18,c_102_17,c_102_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_102_hi = {c_102_32,c_102_31,c_102_30,c_102_29,c_102_28,c_102_27,c_102_26,c_102_25,c_102_24,
    io_out_102_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_103_0 = io_in_0[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_1 = io_in_1[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_2 = io_in_2[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_3 = io_in_3[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_4 = io_in_4[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_5 = io_in_5[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_6 = io_in_6[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_7 = io_in_7[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_8 = io_in_8[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_9 = io_in_9[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_10 = io_in_10[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_11 = io_in_11[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_12 = io_in_12[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_13 = io_in_13[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_14 = io_in_14[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_15 = io_in_15[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_16 = io_in_16[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_17 = io_in_17[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_18 = io_in_18[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_19 = io_in_19[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_20 = io_in_20[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_21 = io_in_21[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_22 = io_in_22[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_23 = io_in_23[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_24 = io_in_24[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_25 = io_in_25[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_26 = io_in_26[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_27 = io_in_27[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_28 = io_in_28[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_29 = io_in_29[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_30 = io_in_30[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_31 = io_in_31[103]; // @[WallaceTest.scala 105:23]
  wire  c_103_32 = io_in_32[103]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_103_lo_lo = {c_103_7,c_103_6,c_103_5,c_103_4,c_103_3,c_103_2,c_103_1,c_103_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_103_lo = {c_103_15,c_103_14,c_103_13,c_103_12,c_103_11,c_103_10,c_103_9,c_103_8,io_out_103_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_103_hi_lo = {c_103_23,c_103_22,c_103_21,c_103_20,c_103_19,c_103_18,c_103_17,c_103_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_103_hi = {c_103_32,c_103_31,c_103_30,c_103_29,c_103_28,c_103_27,c_103_26,c_103_25,c_103_24,
    io_out_103_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_104_0 = io_in_0[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_1 = io_in_1[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_2 = io_in_2[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_3 = io_in_3[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_4 = io_in_4[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_5 = io_in_5[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_6 = io_in_6[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_7 = io_in_7[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_8 = io_in_8[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_9 = io_in_9[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_10 = io_in_10[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_11 = io_in_11[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_12 = io_in_12[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_13 = io_in_13[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_14 = io_in_14[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_15 = io_in_15[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_16 = io_in_16[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_17 = io_in_17[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_18 = io_in_18[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_19 = io_in_19[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_20 = io_in_20[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_21 = io_in_21[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_22 = io_in_22[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_23 = io_in_23[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_24 = io_in_24[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_25 = io_in_25[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_26 = io_in_26[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_27 = io_in_27[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_28 = io_in_28[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_29 = io_in_29[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_30 = io_in_30[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_31 = io_in_31[104]; // @[WallaceTest.scala 105:23]
  wire  c_104_32 = io_in_32[104]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_104_lo_lo = {c_104_7,c_104_6,c_104_5,c_104_4,c_104_3,c_104_2,c_104_1,c_104_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_104_lo = {c_104_15,c_104_14,c_104_13,c_104_12,c_104_11,c_104_10,c_104_9,c_104_8,io_out_104_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_104_hi_lo = {c_104_23,c_104_22,c_104_21,c_104_20,c_104_19,c_104_18,c_104_17,c_104_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_104_hi = {c_104_32,c_104_31,c_104_30,c_104_29,c_104_28,c_104_27,c_104_26,c_104_25,c_104_24,
    io_out_104_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_105_0 = io_in_0[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_1 = io_in_1[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_2 = io_in_2[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_3 = io_in_3[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_4 = io_in_4[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_5 = io_in_5[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_6 = io_in_6[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_7 = io_in_7[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_8 = io_in_8[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_9 = io_in_9[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_10 = io_in_10[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_11 = io_in_11[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_12 = io_in_12[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_13 = io_in_13[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_14 = io_in_14[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_15 = io_in_15[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_16 = io_in_16[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_17 = io_in_17[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_18 = io_in_18[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_19 = io_in_19[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_20 = io_in_20[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_21 = io_in_21[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_22 = io_in_22[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_23 = io_in_23[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_24 = io_in_24[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_25 = io_in_25[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_26 = io_in_26[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_27 = io_in_27[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_28 = io_in_28[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_29 = io_in_29[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_30 = io_in_30[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_31 = io_in_31[105]; // @[WallaceTest.scala 105:23]
  wire  c_105_32 = io_in_32[105]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_105_lo_lo = {c_105_7,c_105_6,c_105_5,c_105_4,c_105_3,c_105_2,c_105_1,c_105_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_105_lo = {c_105_15,c_105_14,c_105_13,c_105_12,c_105_11,c_105_10,c_105_9,c_105_8,io_out_105_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_105_hi_lo = {c_105_23,c_105_22,c_105_21,c_105_20,c_105_19,c_105_18,c_105_17,c_105_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_105_hi = {c_105_32,c_105_31,c_105_30,c_105_29,c_105_28,c_105_27,c_105_26,c_105_25,c_105_24,
    io_out_105_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_106_0 = io_in_0[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_1 = io_in_1[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_2 = io_in_2[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_3 = io_in_3[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_4 = io_in_4[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_5 = io_in_5[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_6 = io_in_6[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_7 = io_in_7[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_8 = io_in_8[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_9 = io_in_9[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_10 = io_in_10[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_11 = io_in_11[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_12 = io_in_12[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_13 = io_in_13[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_14 = io_in_14[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_15 = io_in_15[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_16 = io_in_16[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_17 = io_in_17[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_18 = io_in_18[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_19 = io_in_19[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_20 = io_in_20[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_21 = io_in_21[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_22 = io_in_22[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_23 = io_in_23[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_24 = io_in_24[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_25 = io_in_25[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_26 = io_in_26[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_27 = io_in_27[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_28 = io_in_28[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_29 = io_in_29[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_30 = io_in_30[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_31 = io_in_31[106]; // @[WallaceTest.scala 105:23]
  wire  c_106_32 = io_in_32[106]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_106_lo_lo = {c_106_7,c_106_6,c_106_5,c_106_4,c_106_3,c_106_2,c_106_1,c_106_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_106_lo = {c_106_15,c_106_14,c_106_13,c_106_12,c_106_11,c_106_10,c_106_9,c_106_8,io_out_106_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_106_hi_lo = {c_106_23,c_106_22,c_106_21,c_106_20,c_106_19,c_106_18,c_106_17,c_106_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_106_hi = {c_106_32,c_106_31,c_106_30,c_106_29,c_106_28,c_106_27,c_106_26,c_106_25,c_106_24,
    io_out_106_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_107_0 = io_in_0[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_1 = io_in_1[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_2 = io_in_2[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_3 = io_in_3[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_4 = io_in_4[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_5 = io_in_5[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_6 = io_in_6[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_7 = io_in_7[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_8 = io_in_8[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_9 = io_in_9[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_10 = io_in_10[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_11 = io_in_11[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_12 = io_in_12[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_13 = io_in_13[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_14 = io_in_14[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_15 = io_in_15[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_16 = io_in_16[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_17 = io_in_17[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_18 = io_in_18[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_19 = io_in_19[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_20 = io_in_20[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_21 = io_in_21[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_22 = io_in_22[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_23 = io_in_23[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_24 = io_in_24[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_25 = io_in_25[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_26 = io_in_26[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_27 = io_in_27[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_28 = io_in_28[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_29 = io_in_29[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_30 = io_in_30[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_31 = io_in_31[107]; // @[WallaceTest.scala 105:23]
  wire  c_107_32 = io_in_32[107]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_107_lo_lo = {c_107_7,c_107_6,c_107_5,c_107_4,c_107_3,c_107_2,c_107_1,c_107_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_107_lo = {c_107_15,c_107_14,c_107_13,c_107_12,c_107_11,c_107_10,c_107_9,c_107_8,io_out_107_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_107_hi_lo = {c_107_23,c_107_22,c_107_21,c_107_20,c_107_19,c_107_18,c_107_17,c_107_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_107_hi = {c_107_32,c_107_31,c_107_30,c_107_29,c_107_28,c_107_27,c_107_26,c_107_25,c_107_24,
    io_out_107_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_108_0 = io_in_0[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_1 = io_in_1[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_2 = io_in_2[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_3 = io_in_3[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_4 = io_in_4[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_5 = io_in_5[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_6 = io_in_6[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_7 = io_in_7[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_8 = io_in_8[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_9 = io_in_9[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_10 = io_in_10[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_11 = io_in_11[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_12 = io_in_12[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_13 = io_in_13[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_14 = io_in_14[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_15 = io_in_15[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_16 = io_in_16[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_17 = io_in_17[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_18 = io_in_18[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_19 = io_in_19[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_20 = io_in_20[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_21 = io_in_21[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_22 = io_in_22[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_23 = io_in_23[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_24 = io_in_24[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_25 = io_in_25[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_26 = io_in_26[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_27 = io_in_27[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_28 = io_in_28[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_29 = io_in_29[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_30 = io_in_30[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_31 = io_in_31[108]; // @[WallaceTest.scala 105:23]
  wire  c_108_32 = io_in_32[108]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_108_lo_lo = {c_108_7,c_108_6,c_108_5,c_108_4,c_108_3,c_108_2,c_108_1,c_108_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_108_lo = {c_108_15,c_108_14,c_108_13,c_108_12,c_108_11,c_108_10,c_108_9,c_108_8,io_out_108_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_108_hi_lo = {c_108_23,c_108_22,c_108_21,c_108_20,c_108_19,c_108_18,c_108_17,c_108_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_108_hi = {c_108_32,c_108_31,c_108_30,c_108_29,c_108_28,c_108_27,c_108_26,c_108_25,c_108_24,
    io_out_108_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_109_0 = io_in_0[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_1 = io_in_1[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_2 = io_in_2[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_3 = io_in_3[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_4 = io_in_4[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_5 = io_in_5[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_6 = io_in_6[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_7 = io_in_7[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_8 = io_in_8[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_9 = io_in_9[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_10 = io_in_10[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_11 = io_in_11[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_12 = io_in_12[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_13 = io_in_13[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_14 = io_in_14[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_15 = io_in_15[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_16 = io_in_16[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_17 = io_in_17[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_18 = io_in_18[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_19 = io_in_19[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_20 = io_in_20[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_21 = io_in_21[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_22 = io_in_22[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_23 = io_in_23[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_24 = io_in_24[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_25 = io_in_25[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_26 = io_in_26[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_27 = io_in_27[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_28 = io_in_28[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_29 = io_in_29[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_30 = io_in_30[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_31 = io_in_31[109]; // @[WallaceTest.scala 105:23]
  wire  c_109_32 = io_in_32[109]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_109_lo_lo = {c_109_7,c_109_6,c_109_5,c_109_4,c_109_3,c_109_2,c_109_1,c_109_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_109_lo = {c_109_15,c_109_14,c_109_13,c_109_12,c_109_11,c_109_10,c_109_9,c_109_8,io_out_109_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_109_hi_lo = {c_109_23,c_109_22,c_109_21,c_109_20,c_109_19,c_109_18,c_109_17,c_109_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_109_hi = {c_109_32,c_109_31,c_109_30,c_109_29,c_109_28,c_109_27,c_109_26,c_109_25,c_109_24,
    io_out_109_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_110_0 = io_in_0[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_1 = io_in_1[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_2 = io_in_2[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_3 = io_in_3[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_4 = io_in_4[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_5 = io_in_5[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_6 = io_in_6[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_7 = io_in_7[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_8 = io_in_8[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_9 = io_in_9[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_10 = io_in_10[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_11 = io_in_11[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_12 = io_in_12[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_13 = io_in_13[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_14 = io_in_14[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_15 = io_in_15[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_16 = io_in_16[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_17 = io_in_17[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_18 = io_in_18[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_19 = io_in_19[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_20 = io_in_20[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_21 = io_in_21[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_22 = io_in_22[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_23 = io_in_23[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_24 = io_in_24[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_25 = io_in_25[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_26 = io_in_26[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_27 = io_in_27[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_28 = io_in_28[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_29 = io_in_29[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_30 = io_in_30[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_31 = io_in_31[110]; // @[WallaceTest.scala 105:23]
  wire  c_110_32 = io_in_32[110]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_110_lo_lo = {c_110_7,c_110_6,c_110_5,c_110_4,c_110_3,c_110_2,c_110_1,c_110_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_110_lo = {c_110_15,c_110_14,c_110_13,c_110_12,c_110_11,c_110_10,c_110_9,c_110_8,io_out_110_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_110_hi_lo = {c_110_23,c_110_22,c_110_21,c_110_20,c_110_19,c_110_18,c_110_17,c_110_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_110_hi = {c_110_32,c_110_31,c_110_30,c_110_29,c_110_28,c_110_27,c_110_26,c_110_25,c_110_24,
    io_out_110_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_111_0 = io_in_0[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_1 = io_in_1[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_2 = io_in_2[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_3 = io_in_3[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_4 = io_in_4[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_5 = io_in_5[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_6 = io_in_6[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_7 = io_in_7[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_8 = io_in_8[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_9 = io_in_9[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_10 = io_in_10[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_11 = io_in_11[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_12 = io_in_12[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_13 = io_in_13[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_14 = io_in_14[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_15 = io_in_15[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_16 = io_in_16[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_17 = io_in_17[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_18 = io_in_18[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_19 = io_in_19[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_20 = io_in_20[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_21 = io_in_21[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_22 = io_in_22[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_23 = io_in_23[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_24 = io_in_24[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_25 = io_in_25[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_26 = io_in_26[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_27 = io_in_27[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_28 = io_in_28[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_29 = io_in_29[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_30 = io_in_30[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_31 = io_in_31[111]; // @[WallaceTest.scala 105:23]
  wire  c_111_32 = io_in_32[111]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_111_lo_lo = {c_111_7,c_111_6,c_111_5,c_111_4,c_111_3,c_111_2,c_111_1,c_111_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_111_lo = {c_111_15,c_111_14,c_111_13,c_111_12,c_111_11,c_111_10,c_111_9,c_111_8,io_out_111_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_111_hi_lo = {c_111_23,c_111_22,c_111_21,c_111_20,c_111_19,c_111_18,c_111_17,c_111_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_111_hi = {c_111_32,c_111_31,c_111_30,c_111_29,c_111_28,c_111_27,c_111_26,c_111_25,c_111_24,
    io_out_111_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_112_0 = io_in_0[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_1 = io_in_1[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_2 = io_in_2[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_3 = io_in_3[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_4 = io_in_4[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_5 = io_in_5[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_6 = io_in_6[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_7 = io_in_7[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_8 = io_in_8[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_9 = io_in_9[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_10 = io_in_10[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_11 = io_in_11[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_12 = io_in_12[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_13 = io_in_13[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_14 = io_in_14[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_15 = io_in_15[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_16 = io_in_16[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_17 = io_in_17[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_18 = io_in_18[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_19 = io_in_19[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_20 = io_in_20[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_21 = io_in_21[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_22 = io_in_22[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_23 = io_in_23[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_24 = io_in_24[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_25 = io_in_25[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_26 = io_in_26[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_27 = io_in_27[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_28 = io_in_28[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_29 = io_in_29[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_30 = io_in_30[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_31 = io_in_31[112]; // @[WallaceTest.scala 105:23]
  wire  c_112_32 = io_in_32[112]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_112_lo_lo = {c_112_7,c_112_6,c_112_5,c_112_4,c_112_3,c_112_2,c_112_1,c_112_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_112_lo = {c_112_15,c_112_14,c_112_13,c_112_12,c_112_11,c_112_10,c_112_9,c_112_8,io_out_112_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_112_hi_lo = {c_112_23,c_112_22,c_112_21,c_112_20,c_112_19,c_112_18,c_112_17,c_112_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_112_hi = {c_112_32,c_112_31,c_112_30,c_112_29,c_112_28,c_112_27,c_112_26,c_112_25,c_112_24,
    io_out_112_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_113_0 = io_in_0[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_1 = io_in_1[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_2 = io_in_2[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_3 = io_in_3[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_4 = io_in_4[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_5 = io_in_5[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_6 = io_in_6[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_7 = io_in_7[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_8 = io_in_8[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_9 = io_in_9[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_10 = io_in_10[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_11 = io_in_11[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_12 = io_in_12[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_13 = io_in_13[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_14 = io_in_14[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_15 = io_in_15[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_16 = io_in_16[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_17 = io_in_17[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_18 = io_in_18[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_19 = io_in_19[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_20 = io_in_20[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_21 = io_in_21[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_22 = io_in_22[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_23 = io_in_23[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_24 = io_in_24[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_25 = io_in_25[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_26 = io_in_26[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_27 = io_in_27[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_28 = io_in_28[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_29 = io_in_29[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_30 = io_in_30[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_31 = io_in_31[113]; // @[WallaceTest.scala 105:23]
  wire  c_113_32 = io_in_32[113]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_113_lo_lo = {c_113_7,c_113_6,c_113_5,c_113_4,c_113_3,c_113_2,c_113_1,c_113_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_113_lo = {c_113_15,c_113_14,c_113_13,c_113_12,c_113_11,c_113_10,c_113_9,c_113_8,io_out_113_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_113_hi_lo = {c_113_23,c_113_22,c_113_21,c_113_20,c_113_19,c_113_18,c_113_17,c_113_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_113_hi = {c_113_32,c_113_31,c_113_30,c_113_29,c_113_28,c_113_27,c_113_26,c_113_25,c_113_24,
    io_out_113_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_114_0 = io_in_0[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_1 = io_in_1[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_2 = io_in_2[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_3 = io_in_3[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_4 = io_in_4[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_5 = io_in_5[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_6 = io_in_6[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_7 = io_in_7[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_8 = io_in_8[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_9 = io_in_9[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_10 = io_in_10[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_11 = io_in_11[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_12 = io_in_12[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_13 = io_in_13[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_14 = io_in_14[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_15 = io_in_15[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_16 = io_in_16[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_17 = io_in_17[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_18 = io_in_18[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_19 = io_in_19[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_20 = io_in_20[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_21 = io_in_21[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_22 = io_in_22[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_23 = io_in_23[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_24 = io_in_24[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_25 = io_in_25[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_26 = io_in_26[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_27 = io_in_27[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_28 = io_in_28[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_29 = io_in_29[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_30 = io_in_30[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_31 = io_in_31[114]; // @[WallaceTest.scala 105:23]
  wire  c_114_32 = io_in_32[114]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_114_lo_lo = {c_114_7,c_114_6,c_114_5,c_114_4,c_114_3,c_114_2,c_114_1,c_114_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_114_lo = {c_114_15,c_114_14,c_114_13,c_114_12,c_114_11,c_114_10,c_114_9,c_114_8,io_out_114_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_114_hi_lo = {c_114_23,c_114_22,c_114_21,c_114_20,c_114_19,c_114_18,c_114_17,c_114_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_114_hi = {c_114_32,c_114_31,c_114_30,c_114_29,c_114_28,c_114_27,c_114_26,c_114_25,c_114_24,
    io_out_114_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_115_0 = io_in_0[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_1 = io_in_1[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_2 = io_in_2[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_3 = io_in_3[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_4 = io_in_4[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_5 = io_in_5[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_6 = io_in_6[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_7 = io_in_7[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_8 = io_in_8[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_9 = io_in_9[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_10 = io_in_10[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_11 = io_in_11[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_12 = io_in_12[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_13 = io_in_13[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_14 = io_in_14[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_15 = io_in_15[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_16 = io_in_16[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_17 = io_in_17[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_18 = io_in_18[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_19 = io_in_19[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_20 = io_in_20[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_21 = io_in_21[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_22 = io_in_22[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_23 = io_in_23[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_24 = io_in_24[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_25 = io_in_25[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_26 = io_in_26[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_27 = io_in_27[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_28 = io_in_28[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_29 = io_in_29[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_30 = io_in_30[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_31 = io_in_31[115]; // @[WallaceTest.scala 105:23]
  wire  c_115_32 = io_in_32[115]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_115_lo_lo = {c_115_7,c_115_6,c_115_5,c_115_4,c_115_3,c_115_2,c_115_1,c_115_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_115_lo = {c_115_15,c_115_14,c_115_13,c_115_12,c_115_11,c_115_10,c_115_9,c_115_8,io_out_115_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_115_hi_lo = {c_115_23,c_115_22,c_115_21,c_115_20,c_115_19,c_115_18,c_115_17,c_115_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_115_hi = {c_115_32,c_115_31,c_115_30,c_115_29,c_115_28,c_115_27,c_115_26,c_115_25,c_115_24,
    io_out_115_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_116_0 = io_in_0[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_1 = io_in_1[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_2 = io_in_2[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_3 = io_in_3[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_4 = io_in_4[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_5 = io_in_5[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_6 = io_in_6[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_7 = io_in_7[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_8 = io_in_8[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_9 = io_in_9[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_10 = io_in_10[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_11 = io_in_11[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_12 = io_in_12[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_13 = io_in_13[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_14 = io_in_14[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_15 = io_in_15[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_16 = io_in_16[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_17 = io_in_17[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_18 = io_in_18[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_19 = io_in_19[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_20 = io_in_20[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_21 = io_in_21[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_22 = io_in_22[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_23 = io_in_23[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_24 = io_in_24[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_25 = io_in_25[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_26 = io_in_26[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_27 = io_in_27[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_28 = io_in_28[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_29 = io_in_29[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_30 = io_in_30[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_31 = io_in_31[116]; // @[WallaceTest.scala 105:23]
  wire  c_116_32 = io_in_32[116]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_116_lo_lo = {c_116_7,c_116_6,c_116_5,c_116_4,c_116_3,c_116_2,c_116_1,c_116_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_116_lo = {c_116_15,c_116_14,c_116_13,c_116_12,c_116_11,c_116_10,c_116_9,c_116_8,io_out_116_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_116_hi_lo = {c_116_23,c_116_22,c_116_21,c_116_20,c_116_19,c_116_18,c_116_17,c_116_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_116_hi = {c_116_32,c_116_31,c_116_30,c_116_29,c_116_28,c_116_27,c_116_26,c_116_25,c_116_24,
    io_out_116_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_117_0 = io_in_0[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_1 = io_in_1[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_2 = io_in_2[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_3 = io_in_3[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_4 = io_in_4[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_5 = io_in_5[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_6 = io_in_6[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_7 = io_in_7[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_8 = io_in_8[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_9 = io_in_9[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_10 = io_in_10[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_11 = io_in_11[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_12 = io_in_12[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_13 = io_in_13[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_14 = io_in_14[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_15 = io_in_15[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_16 = io_in_16[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_17 = io_in_17[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_18 = io_in_18[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_19 = io_in_19[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_20 = io_in_20[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_21 = io_in_21[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_22 = io_in_22[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_23 = io_in_23[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_24 = io_in_24[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_25 = io_in_25[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_26 = io_in_26[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_27 = io_in_27[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_28 = io_in_28[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_29 = io_in_29[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_30 = io_in_30[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_31 = io_in_31[117]; // @[WallaceTest.scala 105:23]
  wire  c_117_32 = io_in_32[117]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_117_lo_lo = {c_117_7,c_117_6,c_117_5,c_117_4,c_117_3,c_117_2,c_117_1,c_117_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_117_lo = {c_117_15,c_117_14,c_117_13,c_117_12,c_117_11,c_117_10,c_117_9,c_117_8,io_out_117_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_117_hi_lo = {c_117_23,c_117_22,c_117_21,c_117_20,c_117_19,c_117_18,c_117_17,c_117_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_117_hi = {c_117_32,c_117_31,c_117_30,c_117_29,c_117_28,c_117_27,c_117_26,c_117_25,c_117_24,
    io_out_117_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_118_0 = io_in_0[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_1 = io_in_1[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_2 = io_in_2[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_3 = io_in_3[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_4 = io_in_4[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_5 = io_in_5[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_6 = io_in_6[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_7 = io_in_7[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_8 = io_in_8[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_9 = io_in_9[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_10 = io_in_10[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_11 = io_in_11[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_12 = io_in_12[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_13 = io_in_13[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_14 = io_in_14[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_15 = io_in_15[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_16 = io_in_16[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_17 = io_in_17[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_18 = io_in_18[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_19 = io_in_19[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_20 = io_in_20[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_21 = io_in_21[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_22 = io_in_22[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_23 = io_in_23[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_24 = io_in_24[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_25 = io_in_25[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_26 = io_in_26[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_27 = io_in_27[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_28 = io_in_28[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_29 = io_in_29[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_30 = io_in_30[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_31 = io_in_31[118]; // @[WallaceTest.scala 105:23]
  wire  c_118_32 = io_in_32[118]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_118_lo_lo = {c_118_7,c_118_6,c_118_5,c_118_4,c_118_3,c_118_2,c_118_1,c_118_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_118_lo = {c_118_15,c_118_14,c_118_13,c_118_12,c_118_11,c_118_10,c_118_9,c_118_8,io_out_118_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_118_hi_lo = {c_118_23,c_118_22,c_118_21,c_118_20,c_118_19,c_118_18,c_118_17,c_118_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_118_hi = {c_118_32,c_118_31,c_118_30,c_118_29,c_118_28,c_118_27,c_118_26,c_118_25,c_118_24,
    io_out_118_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_119_0 = io_in_0[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_1 = io_in_1[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_2 = io_in_2[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_3 = io_in_3[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_4 = io_in_4[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_5 = io_in_5[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_6 = io_in_6[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_7 = io_in_7[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_8 = io_in_8[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_9 = io_in_9[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_10 = io_in_10[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_11 = io_in_11[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_12 = io_in_12[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_13 = io_in_13[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_14 = io_in_14[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_15 = io_in_15[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_16 = io_in_16[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_17 = io_in_17[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_18 = io_in_18[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_19 = io_in_19[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_20 = io_in_20[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_21 = io_in_21[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_22 = io_in_22[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_23 = io_in_23[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_24 = io_in_24[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_25 = io_in_25[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_26 = io_in_26[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_27 = io_in_27[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_28 = io_in_28[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_29 = io_in_29[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_30 = io_in_30[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_31 = io_in_31[119]; // @[WallaceTest.scala 105:23]
  wire  c_119_32 = io_in_32[119]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_119_lo_lo = {c_119_7,c_119_6,c_119_5,c_119_4,c_119_3,c_119_2,c_119_1,c_119_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_119_lo = {c_119_15,c_119_14,c_119_13,c_119_12,c_119_11,c_119_10,c_119_9,c_119_8,io_out_119_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_119_hi_lo = {c_119_23,c_119_22,c_119_21,c_119_20,c_119_19,c_119_18,c_119_17,c_119_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_119_hi = {c_119_32,c_119_31,c_119_30,c_119_29,c_119_28,c_119_27,c_119_26,c_119_25,c_119_24,
    io_out_119_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_120_0 = io_in_0[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_1 = io_in_1[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_2 = io_in_2[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_3 = io_in_3[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_4 = io_in_4[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_5 = io_in_5[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_6 = io_in_6[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_7 = io_in_7[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_8 = io_in_8[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_9 = io_in_9[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_10 = io_in_10[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_11 = io_in_11[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_12 = io_in_12[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_13 = io_in_13[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_14 = io_in_14[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_15 = io_in_15[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_16 = io_in_16[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_17 = io_in_17[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_18 = io_in_18[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_19 = io_in_19[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_20 = io_in_20[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_21 = io_in_21[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_22 = io_in_22[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_23 = io_in_23[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_24 = io_in_24[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_25 = io_in_25[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_26 = io_in_26[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_27 = io_in_27[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_28 = io_in_28[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_29 = io_in_29[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_30 = io_in_30[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_31 = io_in_31[120]; // @[WallaceTest.scala 105:23]
  wire  c_120_32 = io_in_32[120]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_120_lo_lo = {c_120_7,c_120_6,c_120_5,c_120_4,c_120_3,c_120_2,c_120_1,c_120_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_120_lo = {c_120_15,c_120_14,c_120_13,c_120_12,c_120_11,c_120_10,c_120_9,c_120_8,io_out_120_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_120_hi_lo = {c_120_23,c_120_22,c_120_21,c_120_20,c_120_19,c_120_18,c_120_17,c_120_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_120_hi = {c_120_32,c_120_31,c_120_30,c_120_29,c_120_28,c_120_27,c_120_26,c_120_25,c_120_24,
    io_out_120_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_121_0 = io_in_0[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_1 = io_in_1[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_2 = io_in_2[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_3 = io_in_3[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_4 = io_in_4[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_5 = io_in_5[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_6 = io_in_6[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_7 = io_in_7[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_8 = io_in_8[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_9 = io_in_9[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_10 = io_in_10[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_11 = io_in_11[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_12 = io_in_12[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_13 = io_in_13[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_14 = io_in_14[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_15 = io_in_15[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_16 = io_in_16[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_17 = io_in_17[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_18 = io_in_18[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_19 = io_in_19[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_20 = io_in_20[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_21 = io_in_21[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_22 = io_in_22[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_23 = io_in_23[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_24 = io_in_24[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_25 = io_in_25[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_26 = io_in_26[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_27 = io_in_27[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_28 = io_in_28[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_29 = io_in_29[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_30 = io_in_30[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_31 = io_in_31[121]; // @[WallaceTest.scala 105:23]
  wire  c_121_32 = io_in_32[121]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_121_lo_lo = {c_121_7,c_121_6,c_121_5,c_121_4,c_121_3,c_121_2,c_121_1,c_121_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_121_lo = {c_121_15,c_121_14,c_121_13,c_121_12,c_121_11,c_121_10,c_121_9,c_121_8,io_out_121_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_121_hi_lo = {c_121_23,c_121_22,c_121_21,c_121_20,c_121_19,c_121_18,c_121_17,c_121_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_121_hi = {c_121_32,c_121_31,c_121_30,c_121_29,c_121_28,c_121_27,c_121_26,c_121_25,c_121_24,
    io_out_121_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_122_0 = io_in_0[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_1 = io_in_1[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_2 = io_in_2[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_3 = io_in_3[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_4 = io_in_4[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_5 = io_in_5[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_6 = io_in_6[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_7 = io_in_7[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_8 = io_in_8[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_9 = io_in_9[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_10 = io_in_10[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_11 = io_in_11[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_12 = io_in_12[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_13 = io_in_13[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_14 = io_in_14[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_15 = io_in_15[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_16 = io_in_16[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_17 = io_in_17[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_18 = io_in_18[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_19 = io_in_19[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_20 = io_in_20[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_21 = io_in_21[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_22 = io_in_22[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_23 = io_in_23[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_24 = io_in_24[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_25 = io_in_25[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_26 = io_in_26[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_27 = io_in_27[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_28 = io_in_28[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_29 = io_in_29[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_30 = io_in_30[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_31 = io_in_31[122]; // @[WallaceTest.scala 105:23]
  wire  c_122_32 = io_in_32[122]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_122_lo_lo = {c_122_7,c_122_6,c_122_5,c_122_4,c_122_3,c_122_2,c_122_1,c_122_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_122_lo = {c_122_15,c_122_14,c_122_13,c_122_12,c_122_11,c_122_10,c_122_9,c_122_8,io_out_122_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_122_hi_lo = {c_122_23,c_122_22,c_122_21,c_122_20,c_122_19,c_122_18,c_122_17,c_122_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_122_hi = {c_122_32,c_122_31,c_122_30,c_122_29,c_122_28,c_122_27,c_122_26,c_122_25,c_122_24,
    io_out_122_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_123_0 = io_in_0[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_1 = io_in_1[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_2 = io_in_2[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_3 = io_in_3[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_4 = io_in_4[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_5 = io_in_5[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_6 = io_in_6[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_7 = io_in_7[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_8 = io_in_8[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_9 = io_in_9[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_10 = io_in_10[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_11 = io_in_11[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_12 = io_in_12[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_13 = io_in_13[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_14 = io_in_14[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_15 = io_in_15[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_16 = io_in_16[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_17 = io_in_17[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_18 = io_in_18[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_19 = io_in_19[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_20 = io_in_20[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_21 = io_in_21[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_22 = io_in_22[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_23 = io_in_23[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_24 = io_in_24[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_25 = io_in_25[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_26 = io_in_26[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_27 = io_in_27[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_28 = io_in_28[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_29 = io_in_29[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_30 = io_in_30[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_31 = io_in_31[123]; // @[WallaceTest.scala 105:23]
  wire  c_123_32 = io_in_32[123]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_123_lo_lo = {c_123_7,c_123_6,c_123_5,c_123_4,c_123_3,c_123_2,c_123_1,c_123_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_123_lo = {c_123_15,c_123_14,c_123_13,c_123_12,c_123_11,c_123_10,c_123_9,c_123_8,io_out_123_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_123_hi_lo = {c_123_23,c_123_22,c_123_21,c_123_20,c_123_19,c_123_18,c_123_17,c_123_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_123_hi = {c_123_32,c_123_31,c_123_30,c_123_29,c_123_28,c_123_27,c_123_26,c_123_25,c_123_24,
    io_out_123_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_124_0 = io_in_0[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_1 = io_in_1[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_2 = io_in_2[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_3 = io_in_3[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_4 = io_in_4[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_5 = io_in_5[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_6 = io_in_6[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_7 = io_in_7[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_8 = io_in_8[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_9 = io_in_9[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_10 = io_in_10[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_11 = io_in_11[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_12 = io_in_12[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_13 = io_in_13[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_14 = io_in_14[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_15 = io_in_15[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_16 = io_in_16[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_17 = io_in_17[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_18 = io_in_18[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_19 = io_in_19[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_20 = io_in_20[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_21 = io_in_21[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_22 = io_in_22[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_23 = io_in_23[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_24 = io_in_24[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_25 = io_in_25[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_26 = io_in_26[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_27 = io_in_27[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_28 = io_in_28[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_29 = io_in_29[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_30 = io_in_30[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_31 = io_in_31[124]; // @[WallaceTest.scala 105:23]
  wire  c_124_32 = io_in_32[124]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_124_lo_lo = {c_124_7,c_124_6,c_124_5,c_124_4,c_124_3,c_124_2,c_124_1,c_124_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_124_lo = {c_124_15,c_124_14,c_124_13,c_124_12,c_124_11,c_124_10,c_124_9,c_124_8,io_out_124_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_124_hi_lo = {c_124_23,c_124_22,c_124_21,c_124_20,c_124_19,c_124_18,c_124_17,c_124_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_124_hi = {c_124_32,c_124_31,c_124_30,c_124_29,c_124_28,c_124_27,c_124_26,c_124_25,c_124_24,
    io_out_124_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_125_0 = io_in_0[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_1 = io_in_1[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_2 = io_in_2[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_3 = io_in_3[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_4 = io_in_4[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_5 = io_in_5[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_6 = io_in_6[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_7 = io_in_7[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_8 = io_in_8[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_9 = io_in_9[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_10 = io_in_10[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_11 = io_in_11[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_12 = io_in_12[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_13 = io_in_13[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_14 = io_in_14[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_15 = io_in_15[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_16 = io_in_16[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_17 = io_in_17[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_18 = io_in_18[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_19 = io_in_19[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_20 = io_in_20[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_21 = io_in_21[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_22 = io_in_22[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_23 = io_in_23[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_24 = io_in_24[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_25 = io_in_25[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_26 = io_in_26[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_27 = io_in_27[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_28 = io_in_28[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_29 = io_in_29[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_30 = io_in_30[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_31 = io_in_31[125]; // @[WallaceTest.scala 105:23]
  wire  c_125_32 = io_in_32[125]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_125_lo_lo = {c_125_7,c_125_6,c_125_5,c_125_4,c_125_3,c_125_2,c_125_1,c_125_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_125_lo = {c_125_15,c_125_14,c_125_13,c_125_12,c_125_11,c_125_10,c_125_9,c_125_8,io_out_125_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_125_hi_lo = {c_125_23,c_125_22,c_125_21,c_125_20,c_125_19,c_125_18,c_125_17,c_125_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_125_hi = {c_125_32,c_125_31,c_125_30,c_125_29,c_125_28,c_125_27,c_125_26,c_125_25,c_125_24,
    io_out_125_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_126_0 = io_in_0[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_1 = io_in_1[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_2 = io_in_2[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_3 = io_in_3[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_4 = io_in_4[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_5 = io_in_5[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_6 = io_in_6[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_7 = io_in_7[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_8 = io_in_8[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_9 = io_in_9[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_10 = io_in_10[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_11 = io_in_11[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_12 = io_in_12[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_13 = io_in_13[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_14 = io_in_14[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_15 = io_in_15[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_16 = io_in_16[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_17 = io_in_17[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_18 = io_in_18[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_19 = io_in_19[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_20 = io_in_20[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_21 = io_in_21[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_22 = io_in_22[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_23 = io_in_23[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_24 = io_in_24[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_25 = io_in_25[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_26 = io_in_26[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_27 = io_in_27[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_28 = io_in_28[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_29 = io_in_29[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_30 = io_in_30[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_31 = io_in_31[126]; // @[WallaceTest.scala 105:23]
  wire  c_126_32 = io_in_32[126]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_126_lo_lo = {c_126_7,c_126_6,c_126_5,c_126_4,c_126_3,c_126_2,c_126_1,c_126_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_126_lo = {c_126_15,c_126_14,c_126_13,c_126_12,c_126_11,c_126_10,c_126_9,c_126_8,io_out_126_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_126_hi_lo = {c_126_23,c_126_22,c_126_21,c_126_20,c_126_19,c_126_18,c_126_17,c_126_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_126_hi = {c_126_32,c_126_31,c_126_30,c_126_29,c_126_28,c_126_27,c_126_26,c_126_25,c_126_24,
    io_out_126_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_127_0 = io_in_0[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_1 = io_in_1[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_2 = io_in_2[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_3 = io_in_3[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_4 = io_in_4[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_5 = io_in_5[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_6 = io_in_6[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_7 = io_in_7[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_8 = io_in_8[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_9 = io_in_9[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_10 = io_in_10[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_11 = io_in_11[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_12 = io_in_12[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_13 = io_in_13[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_14 = io_in_14[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_15 = io_in_15[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_16 = io_in_16[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_17 = io_in_17[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_18 = io_in_18[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_19 = io_in_19[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_20 = io_in_20[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_21 = io_in_21[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_22 = io_in_22[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_23 = io_in_23[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_24 = io_in_24[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_25 = io_in_25[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_26 = io_in_26[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_27 = io_in_27[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_28 = io_in_28[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_29 = io_in_29[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_30 = io_in_30[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_31 = io_in_31[127]; // @[WallaceTest.scala 105:23]
  wire  c_127_32 = io_in_32[127]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_127_lo_lo = {c_127_7,c_127_6,c_127_5,c_127_4,c_127_3,c_127_2,c_127_1,c_127_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_127_lo = {c_127_15,c_127_14,c_127_13,c_127_12,c_127_11,c_127_10,c_127_9,c_127_8,io_out_127_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_127_hi_lo = {c_127_23,c_127_22,c_127_21,c_127_20,c_127_19,c_127_18,c_127_17,c_127_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_127_hi = {c_127_32,c_127_31,c_127_30,c_127_29,c_127_28,c_127_27,c_127_26,c_127_25,c_127_24,
    io_out_127_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_128_0 = io_in_0[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_1 = io_in_1[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_2 = io_in_2[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_3 = io_in_3[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_4 = io_in_4[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_5 = io_in_5[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_6 = io_in_6[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_7 = io_in_7[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_8 = io_in_8[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_9 = io_in_9[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_10 = io_in_10[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_11 = io_in_11[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_12 = io_in_12[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_13 = io_in_13[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_14 = io_in_14[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_15 = io_in_15[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_16 = io_in_16[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_17 = io_in_17[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_18 = io_in_18[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_19 = io_in_19[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_20 = io_in_20[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_21 = io_in_21[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_22 = io_in_22[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_23 = io_in_23[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_24 = io_in_24[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_25 = io_in_25[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_26 = io_in_26[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_27 = io_in_27[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_28 = io_in_28[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_29 = io_in_29[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_30 = io_in_30[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_31 = io_in_31[128]; // @[WallaceTest.scala 105:23]
  wire  c_128_32 = io_in_32[128]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_128_lo_lo = {c_128_7,c_128_6,c_128_5,c_128_4,c_128_3,c_128_2,c_128_1,c_128_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_128_lo = {c_128_15,c_128_14,c_128_13,c_128_12,c_128_11,c_128_10,c_128_9,c_128_8,io_out_128_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_128_hi_lo = {c_128_23,c_128_22,c_128_21,c_128_20,c_128_19,c_128_18,c_128_17,c_128_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_128_hi = {c_128_32,c_128_31,c_128_30,c_128_29,c_128_28,c_128_27,c_128_26,c_128_25,c_128_24,
    io_out_128_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_129_0 = io_in_0[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_1 = io_in_1[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_2 = io_in_2[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_3 = io_in_3[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_4 = io_in_4[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_5 = io_in_5[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_6 = io_in_6[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_7 = io_in_7[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_8 = io_in_8[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_9 = io_in_9[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_10 = io_in_10[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_11 = io_in_11[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_12 = io_in_12[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_13 = io_in_13[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_14 = io_in_14[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_15 = io_in_15[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_16 = io_in_16[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_17 = io_in_17[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_18 = io_in_18[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_19 = io_in_19[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_20 = io_in_20[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_21 = io_in_21[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_22 = io_in_22[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_23 = io_in_23[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_24 = io_in_24[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_25 = io_in_25[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_26 = io_in_26[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_27 = io_in_27[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_28 = io_in_28[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_29 = io_in_29[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_30 = io_in_30[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_31 = io_in_31[129]; // @[WallaceTest.scala 105:23]
  wire  c_129_32 = io_in_32[129]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_129_lo_lo = {c_129_7,c_129_6,c_129_5,c_129_4,c_129_3,c_129_2,c_129_1,c_129_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_129_lo = {c_129_15,c_129_14,c_129_13,c_129_12,c_129_11,c_129_10,c_129_9,c_129_8,io_out_129_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_129_hi_lo = {c_129_23,c_129_22,c_129_21,c_129_20,c_129_19,c_129_18,c_129_17,c_129_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_129_hi = {c_129_32,c_129_31,c_129_30,c_129_29,c_129_28,c_129_27,c_129_26,c_129_25,c_129_24,
    io_out_129_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_130_0 = io_in_0[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_1 = io_in_1[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_2 = io_in_2[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_3 = io_in_3[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_4 = io_in_4[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_5 = io_in_5[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_6 = io_in_6[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_7 = io_in_7[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_8 = io_in_8[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_9 = io_in_9[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_10 = io_in_10[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_11 = io_in_11[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_12 = io_in_12[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_13 = io_in_13[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_14 = io_in_14[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_15 = io_in_15[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_16 = io_in_16[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_17 = io_in_17[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_18 = io_in_18[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_19 = io_in_19[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_20 = io_in_20[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_21 = io_in_21[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_22 = io_in_22[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_23 = io_in_23[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_24 = io_in_24[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_25 = io_in_25[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_26 = io_in_26[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_27 = io_in_27[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_28 = io_in_28[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_29 = io_in_29[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_30 = io_in_30[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_31 = io_in_31[130]; // @[WallaceTest.scala 105:23]
  wire  c_130_32 = io_in_32[130]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_130_lo_lo = {c_130_7,c_130_6,c_130_5,c_130_4,c_130_3,c_130_2,c_130_1,c_130_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_130_lo = {c_130_15,c_130_14,c_130_13,c_130_12,c_130_11,c_130_10,c_130_9,c_130_8,io_out_130_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_130_hi_lo = {c_130_23,c_130_22,c_130_21,c_130_20,c_130_19,c_130_18,c_130_17,c_130_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_130_hi = {c_130_32,c_130_31,c_130_30,c_130_29,c_130_28,c_130_27,c_130_26,c_130_25,c_130_24,
    io_out_130_hi_lo}; // @[WallaceTest.scala 107:20]
  wire  c_131_0 = io_in_0[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_1 = io_in_1[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_2 = io_in_2[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_3 = io_in_3[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_4 = io_in_4[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_5 = io_in_5[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_6 = io_in_6[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_7 = io_in_7[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_8 = io_in_8[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_9 = io_in_9[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_10 = io_in_10[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_11 = io_in_11[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_12 = io_in_12[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_13 = io_in_13[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_14 = io_in_14[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_15 = io_in_15[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_16 = io_in_16[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_17 = io_in_17[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_18 = io_in_18[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_19 = io_in_19[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_20 = io_in_20[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_21 = io_in_21[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_22 = io_in_22[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_23 = io_in_23[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_24 = io_in_24[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_25 = io_in_25[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_26 = io_in_26[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_27 = io_in_27[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_28 = io_in_28[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_29 = io_in_29[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_30 = io_in_30[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_31 = io_in_31[131]; // @[WallaceTest.scala 105:23]
  wire  c_131_32 = io_in_32[131]; // @[WallaceTest.scala 105:23]
  wire [7:0] io_out_131_lo_lo = {c_131_7,c_131_6,c_131_5,c_131_4,c_131_3,c_131_2,c_131_1,c_131_0}; // @[WallaceTest.scala 107:20]
  wire [15:0] io_out_131_lo = {c_131_15,c_131_14,c_131_13,c_131_12,c_131_11,c_131_10,c_131_9,c_131_8,io_out_131_lo_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_out_131_hi_lo = {c_131_23,c_131_22,c_131_21,c_131_20,c_131_19,c_131_18,c_131_17,c_131_16}; // @[WallaceTest.scala 107:20]
  wire [16:0] io_out_131_hi = {c_131_32,c_131_31,c_131_30,c_131_29,c_131_28,c_131_27,c_131_26,c_131_25,c_131_24,
    io_out_131_hi_lo}; // @[WallaceTest.scala 107:20]
  wire [7:0] io_cout_lo_lo = {io_cin_7,io_cin_6,io_cin_5,io_cin_4,io_cin_3,io_cin_2,io_cin_1,io_cin_0}; // @[WallaceTest.scala 115:19]
  wire [7:0] io_cout_hi_lo = {io_cin_23,io_cin_22,io_cin_21,io_cin_20,io_cin_19,io_cin_18,io_cin_17,io_cin_16}; // @[WallaceTest.scala 115:19]
  wire [16:0] io_cout_hi = {io_cin_32,io_cin_31,io_cin_30,io_cin_29,io_cin_28,io_cin_27,io_cin_26,io_cin_25,io_cin_24,
    io_cout_hi_lo}; // @[WallaceTest.scala 115:19]
  wire [32:0] _io_cout_T = {io_cout_hi,io_cin_15,io_cin_14,io_cin_13,io_cin_12,io_cin_11,io_cin_10,io_cin_9,io_cin_8,
    io_cout_lo_lo}; // @[WallaceTest.scala 115:19]
  assign io_out_0 = {io_out_0_hi,io_out_0_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_1 = {io_out_1_hi,io_out_1_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_2 = {io_out_2_hi,io_out_2_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_3 = {io_out_3_hi,io_out_3_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_4 = {io_out_4_hi,io_out_4_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_5 = {io_out_5_hi,io_out_5_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_6 = {io_out_6_hi,io_out_6_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_7 = {io_out_7_hi,io_out_7_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_8 = {io_out_8_hi,io_out_8_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_9 = {io_out_9_hi,io_out_9_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_10 = {io_out_10_hi,io_out_10_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_11 = {io_out_11_hi,io_out_11_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_12 = {io_out_12_hi,io_out_12_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_13 = {io_out_13_hi,io_out_13_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_14 = {io_out_14_hi,io_out_14_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_15 = {io_out_15_hi,io_out_15_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_16 = {io_out_16_hi,io_out_16_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_17 = {io_out_17_hi,io_out_17_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_18 = {io_out_18_hi,io_out_18_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_19 = {io_out_19_hi,io_out_19_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_20 = {io_out_20_hi,io_out_20_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_21 = {io_out_21_hi,io_out_21_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_22 = {io_out_22_hi,io_out_22_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_23 = {io_out_23_hi,io_out_23_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_24 = {io_out_24_hi,io_out_24_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_25 = {io_out_25_hi,io_out_25_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_26 = {io_out_26_hi,io_out_26_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_27 = {io_out_27_hi,io_out_27_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_28 = {io_out_28_hi,io_out_28_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_29 = {io_out_29_hi,io_out_29_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_30 = {io_out_30_hi,io_out_30_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_31 = {io_out_31_hi,io_out_31_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_32 = {io_out_32_hi,io_out_32_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_33 = {io_out_33_hi,io_out_33_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_34 = {io_out_34_hi,io_out_34_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_35 = {io_out_35_hi,io_out_35_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_36 = {io_out_36_hi,io_out_36_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_37 = {io_out_37_hi,io_out_37_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_38 = {io_out_38_hi,io_out_38_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_39 = {io_out_39_hi,io_out_39_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_40 = {io_out_40_hi,io_out_40_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_41 = {io_out_41_hi,io_out_41_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_42 = {io_out_42_hi,io_out_42_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_43 = {io_out_43_hi,io_out_43_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_44 = {io_out_44_hi,io_out_44_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_45 = {io_out_45_hi,io_out_45_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_46 = {io_out_46_hi,io_out_46_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_47 = {io_out_47_hi,io_out_47_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_48 = {io_out_48_hi,io_out_48_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_49 = {io_out_49_hi,io_out_49_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_50 = {io_out_50_hi,io_out_50_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_51 = {io_out_51_hi,io_out_51_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_52 = {io_out_52_hi,io_out_52_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_53 = {io_out_53_hi,io_out_53_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_54 = {io_out_54_hi,io_out_54_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_55 = {io_out_55_hi,io_out_55_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_56 = {io_out_56_hi,io_out_56_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_57 = {io_out_57_hi,io_out_57_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_58 = {io_out_58_hi,io_out_58_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_59 = {io_out_59_hi,io_out_59_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_60 = {io_out_60_hi,io_out_60_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_61 = {io_out_61_hi,io_out_61_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_62 = {io_out_62_hi,io_out_62_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_63 = {io_out_63_hi,io_out_63_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_64 = {io_out_64_hi,io_out_64_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_65 = {io_out_65_hi,io_out_65_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_66 = {io_out_66_hi,io_out_66_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_67 = {io_out_67_hi,io_out_67_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_68 = {io_out_68_hi,io_out_68_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_69 = {io_out_69_hi,io_out_69_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_70 = {io_out_70_hi,io_out_70_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_71 = {io_out_71_hi,io_out_71_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_72 = {io_out_72_hi,io_out_72_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_73 = {io_out_73_hi,io_out_73_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_74 = {io_out_74_hi,io_out_74_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_75 = {io_out_75_hi,io_out_75_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_76 = {io_out_76_hi,io_out_76_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_77 = {io_out_77_hi,io_out_77_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_78 = {io_out_78_hi,io_out_78_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_79 = {io_out_79_hi,io_out_79_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_80 = {io_out_80_hi,io_out_80_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_81 = {io_out_81_hi,io_out_81_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_82 = {io_out_82_hi,io_out_82_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_83 = {io_out_83_hi,io_out_83_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_84 = {io_out_84_hi,io_out_84_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_85 = {io_out_85_hi,io_out_85_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_86 = {io_out_86_hi,io_out_86_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_87 = {io_out_87_hi,io_out_87_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_88 = {io_out_88_hi,io_out_88_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_89 = {io_out_89_hi,io_out_89_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_90 = {io_out_90_hi,io_out_90_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_91 = {io_out_91_hi,io_out_91_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_92 = {io_out_92_hi,io_out_92_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_93 = {io_out_93_hi,io_out_93_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_94 = {io_out_94_hi,io_out_94_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_95 = {io_out_95_hi,io_out_95_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_96 = {io_out_96_hi,io_out_96_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_97 = {io_out_97_hi,io_out_97_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_98 = {io_out_98_hi,io_out_98_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_99 = {io_out_99_hi,io_out_99_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_100 = {io_out_100_hi,io_out_100_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_101 = {io_out_101_hi,io_out_101_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_102 = {io_out_102_hi,io_out_102_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_103 = {io_out_103_hi,io_out_103_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_104 = {io_out_104_hi,io_out_104_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_105 = {io_out_105_hi,io_out_105_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_106 = {io_out_106_hi,io_out_106_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_107 = {io_out_107_hi,io_out_107_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_108 = {io_out_108_hi,io_out_108_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_109 = {io_out_109_hi,io_out_109_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_110 = {io_out_110_hi,io_out_110_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_111 = {io_out_111_hi,io_out_111_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_112 = {io_out_112_hi,io_out_112_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_113 = {io_out_113_hi,io_out_113_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_114 = {io_out_114_hi,io_out_114_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_115 = {io_out_115_hi,io_out_115_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_116 = {io_out_116_hi,io_out_116_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_117 = {io_out_117_hi,io_out_117_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_118 = {io_out_118_hi,io_out_118_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_119 = {io_out_119_hi,io_out_119_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_120 = {io_out_120_hi,io_out_120_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_121 = {io_out_121_hi,io_out_121_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_122 = {io_out_122_hi,io_out_122_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_123 = {io_out_123_hi,io_out_123_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_124 = {io_out_124_hi,io_out_124_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_125 = {io_out_125_hi,io_out_125_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_126 = {io_out_126_hi,io_out_126_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_127 = {io_out_127_hi,io_out_127_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_128 = {io_out_128_hi,io_out_128_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_129 = {io_out_129_hi,io_out_129_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_130 = {io_out_130_hi,io_out_130_lo}; // @[WallaceTest.scala 107:20]
  assign io_out_131 = {io_out_131_hi,io_out_131_lo}; // @[WallaceTest.scala 107:20]
  assign io_cout = _io_cout_T[31:0]; // @[WallaceTest.scala 115:25]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[0] == c__0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[0] == c__0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[1] == c__1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[1] == c__1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[2] == c__2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[2] == c__2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[3] == c__3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[3] == c__3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[4] == c__4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[4] == c__4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[5] == c__5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[5] == c__5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[6] == c__6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[6] == c__6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[7] == c__7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[7] == c__7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[8] == c__8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[8] == c__8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[9] == c__9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[9] == c__9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[10] == c__10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[10] == c__10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[11] == c__11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[11] == c__11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[12] == c__12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[12] == c__12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[13] == c__13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[13] == c__13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[14] == c__14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[14] == c__14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[15] == c__15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[15] == c__15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[16] == c__16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[16] == c__16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[17] == c__17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[17] == c__17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[18] == c__18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[18] == c__18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[19] == c__19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[19] == c__19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[20] == c__20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[20] == c__20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[21] == c__21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[21] == c__21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[22] == c__22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[22] == c__22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[23] == c__23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[23] == c__23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[24] == c__24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[24] == c__24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[25] == c__25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[25] == c__25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[26] == c__26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[26] == c__26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[27] == c__27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[27] == c__27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[28] == c__28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[28] == c__28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[29] == c__29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[29] == c__29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[30] == c__30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[30] == c__30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[31] == c__31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[31] == c__31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_0[32] == c__32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_0[32] == c__32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[0] == c_1_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[0] == c_1_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[1] == c_1_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[1] == c_1_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[2] == c_1_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[2] == c_1_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[3] == c_1_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[3] == c_1_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[4] == c_1_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[4] == c_1_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[5] == c_1_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[5] == c_1_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[6] == c_1_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[6] == c_1_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[7] == c_1_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[7] == c_1_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[8] == c_1_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[8] == c_1_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[9] == c_1_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[9] == c_1_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[10] == c_1_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[10] == c_1_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[11] == c_1_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[11] == c_1_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[12] == c_1_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[12] == c_1_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[13] == c_1_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[13] == c_1_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[14] == c_1_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[14] == c_1_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[15] == c_1_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[15] == c_1_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[16] == c_1_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[16] == c_1_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[17] == c_1_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[17] == c_1_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[18] == c_1_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[18] == c_1_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[19] == c_1_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[19] == c_1_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[20] == c_1_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[20] == c_1_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[21] == c_1_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[21] == c_1_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[22] == c_1_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[22] == c_1_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[23] == c_1_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[23] == c_1_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[24] == c_1_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[24] == c_1_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[25] == c_1_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[25] == c_1_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[26] == c_1_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[26] == c_1_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[27] == c_1_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[27] == c_1_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[28] == c_1_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[28] == c_1_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[29] == c_1_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[29] == c_1_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[30] == c_1_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[30] == c_1_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[31] == c_1_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[31] == c_1_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_1[32] == c_1_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_1[32] == c_1_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[0] == c_2_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[0] == c_2_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[1] == c_2_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[1] == c_2_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[2] == c_2_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[2] == c_2_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[3] == c_2_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[3] == c_2_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[4] == c_2_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[4] == c_2_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[5] == c_2_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[5] == c_2_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[6] == c_2_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[6] == c_2_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[7] == c_2_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[7] == c_2_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[8] == c_2_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[8] == c_2_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[9] == c_2_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[9] == c_2_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[10] == c_2_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[10] == c_2_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[11] == c_2_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[11] == c_2_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[12] == c_2_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[12] == c_2_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[13] == c_2_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[13] == c_2_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[14] == c_2_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[14] == c_2_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[15] == c_2_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[15] == c_2_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[16] == c_2_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[16] == c_2_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[17] == c_2_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[17] == c_2_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[18] == c_2_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[18] == c_2_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[19] == c_2_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[19] == c_2_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[20] == c_2_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[20] == c_2_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[21] == c_2_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[21] == c_2_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[22] == c_2_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[22] == c_2_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[23] == c_2_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[23] == c_2_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[24] == c_2_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[24] == c_2_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[25] == c_2_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[25] == c_2_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[26] == c_2_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[26] == c_2_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[27] == c_2_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[27] == c_2_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[28] == c_2_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[28] == c_2_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[29] == c_2_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[29] == c_2_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[30] == c_2_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[30] == c_2_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[31] == c_2_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[31] == c_2_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_2[32] == c_2_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_2[32] == c_2_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[0] == c_3_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[0] == c_3_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[1] == c_3_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[1] == c_3_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[2] == c_3_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[2] == c_3_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[3] == c_3_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[3] == c_3_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[4] == c_3_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[4] == c_3_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[5] == c_3_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[5] == c_3_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[6] == c_3_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[6] == c_3_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[7] == c_3_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[7] == c_3_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[8] == c_3_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[8] == c_3_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[9] == c_3_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[9] == c_3_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[10] == c_3_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[10] == c_3_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[11] == c_3_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[11] == c_3_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[12] == c_3_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[12] == c_3_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[13] == c_3_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[13] == c_3_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[14] == c_3_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[14] == c_3_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[15] == c_3_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[15] == c_3_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[16] == c_3_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[16] == c_3_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[17] == c_3_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[17] == c_3_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[18] == c_3_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[18] == c_3_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[19] == c_3_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[19] == c_3_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[20] == c_3_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[20] == c_3_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[21] == c_3_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[21] == c_3_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[22] == c_3_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[22] == c_3_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[23] == c_3_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[23] == c_3_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[24] == c_3_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[24] == c_3_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[25] == c_3_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[25] == c_3_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[26] == c_3_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[26] == c_3_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[27] == c_3_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[27] == c_3_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[28] == c_3_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[28] == c_3_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[29] == c_3_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[29] == c_3_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[30] == c_3_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[30] == c_3_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[31] == c_3_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[31] == c_3_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_3[32] == c_3_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_3[32] == c_3_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[0] == c_4_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[0] == c_4_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[1] == c_4_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[1] == c_4_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[2] == c_4_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[2] == c_4_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[3] == c_4_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[3] == c_4_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[4] == c_4_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[4] == c_4_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[5] == c_4_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[5] == c_4_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[6] == c_4_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[6] == c_4_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[7] == c_4_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[7] == c_4_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[8] == c_4_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[8] == c_4_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[9] == c_4_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[9] == c_4_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[10] == c_4_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[10] == c_4_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[11] == c_4_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[11] == c_4_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[12] == c_4_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[12] == c_4_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[13] == c_4_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[13] == c_4_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[14] == c_4_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[14] == c_4_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[15] == c_4_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[15] == c_4_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[16] == c_4_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[16] == c_4_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[17] == c_4_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[17] == c_4_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[18] == c_4_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[18] == c_4_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[19] == c_4_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[19] == c_4_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[20] == c_4_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[20] == c_4_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[21] == c_4_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[21] == c_4_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[22] == c_4_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[22] == c_4_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[23] == c_4_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[23] == c_4_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[24] == c_4_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[24] == c_4_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[25] == c_4_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[25] == c_4_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[26] == c_4_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[26] == c_4_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[27] == c_4_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[27] == c_4_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[28] == c_4_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[28] == c_4_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[29] == c_4_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[29] == c_4_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[30] == c_4_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[30] == c_4_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[31] == c_4_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[31] == c_4_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_4[32] == c_4_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_4[32] == c_4_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[0] == c_5_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[0] == c_5_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[1] == c_5_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[1] == c_5_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[2] == c_5_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[2] == c_5_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[3] == c_5_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[3] == c_5_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[4] == c_5_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[4] == c_5_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[5] == c_5_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[5] == c_5_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[6] == c_5_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[6] == c_5_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[7] == c_5_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[7] == c_5_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[8] == c_5_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[8] == c_5_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[9] == c_5_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[9] == c_5_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[10] == c_5_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[10] == c_5_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[11] == c_5_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[11] == c_5_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[12] == c_5_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[12] == c_5_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[13] == c_5_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[13] == c_5_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[14] == c_5_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[14] == c_5_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[15] == c_5_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[15] == c_5_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[16] == c_5_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[16] == c_5_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[17] == c_5_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[17] == c_5_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[18] == c_5_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[18] == c_5_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[19] == c_5_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[19] == c_5_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[20] == c_5_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[20] == c_5_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[21] == c_5_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[21] == c_5_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[22] == c_5_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[22] == c_5_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[23] == c_5_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[23] == c_5_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[24] == c_5_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[24] == c_5_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[25] == c_5_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[25] == c_5_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[26] == c_5_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[26] == c_5_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[27] == c_5_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[27] == c_5_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[28] == c_5_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[28] == c_5_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[29] == c_5_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[29] == c_5_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[30] == c_5_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[30] == c_5_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[31] == c_5_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[31] == c_5_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_5[32] == c_5_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_5[32] == c_5_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[0] == c_6_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[0] == c_6_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[1] == c_6_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[1] == c_6_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[2] == c_6_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[2] == c_6_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[3] == c_6_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[3] == c_6_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[4] == c_6_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[4] == c_6_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[5] == c_6_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[5] == c_6_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[6] == c_6_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[6] == c_6_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[7] == c_6_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[7] == c_6_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[8] == c_6_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[8] == c_6_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[9] == c_6_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[9] == c_6_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[10] == c_6_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[10] == c_6_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[11] == c_6_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[11] == c_6_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[12] == c_6_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[12] == c_6_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[13] == c_6_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[13] == c_6_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[14] == c_6_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[14] == c_6_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[15] == c_6_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[15] == c_6_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[16] == c_6_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[16] == c_6_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[17] == c_6_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[17] == c_6_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[18] == c_6_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[18] == c_6_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[19] == c_6_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[19] == c_6_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[20] == c_6_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[20] == c_6_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[21] == c_6_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[21] == c_6_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[22] == c_6_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[22] == c_6_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[23] == c_6_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[23] == c_6_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[24] == c_6_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[24] == c_6_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[25] == c_6_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[25] == c_6_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[26] == c_6_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[26] == c_6_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[27] == c_6_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[27] == c_6_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[28] == c_6_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[28] == c_6_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[29] == c_6_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[29] == c_6_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[30] == c_6_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[30] == c_6_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[31] == c_6_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[31] == c_6_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_6[32] == c_6_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_6[32] == c_6_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[0] == c_7_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[0] == c_7_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[1] == c_7_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[1] == c_7_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[2] == c_7_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[2] == c_7_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[3] == c_7_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[3] == c_7_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[4] == c_7_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[4] == c_7_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[5] == c_7_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[5] == c_7_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[6] == c_7_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[6] == c_7_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[7] == c_7_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[7] == c_7_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[8] == c_7_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[8] == c_7_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[9] == c_7_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[9] == c_7_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[10] == c_7_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[10] == c_7_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[11] == c_7_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[11] == c_7_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[12] == c_7_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[12] == c_7_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[13] == c_7_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[13] == c_7_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[14] == c_7_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[14] == c_7_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[15] == c_7_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[15] == c_7_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[16] == c_7_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[16] == c_7_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[17] == c_7_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[17] == c_7_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[18] == c_7_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[18] == c_7_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[19] == c_7_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[19] == c_7_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[20] == c_7_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[20] == c_7_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[21] == c_7_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[21] == c_7_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[22] == c_7_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[22] == c_7_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[23] == c_7_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[23] == c_7_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[24] == c_7_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[24] == c_7_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[25] == c_7_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[25] == c_7_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[26] == c_7_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[26] == c_7_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[27] == c_7_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[27] == c_7_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[28] == c_7_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[28] == c_7_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[29] == c_7_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[29] == c_7_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[30] == c_7_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[30] == c_7_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[31] == c_7_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[31] == c_7_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_7[32] == c_7_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_7[32] == c_7_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[0] == c_8_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[0] == c_8_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[1] == c_8_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[1] == c_8_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[2] == c_8_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[2] == c_8_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[3] == c_8_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[3] == c_8_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[4] == c_8_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[4] == c_8_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[5] == c_8_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[5] == c_8_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[6] == c_8_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[6] == c_8_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[7] == c_8_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[7] == c_8_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[8] == c_8_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[8] == c_8_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[9] == c_8_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[9] == c_8_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[10] == c_8_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[10] == c_8_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[11] == c_8_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[11] == c_8_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[12] == c_8_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[12] == c_8_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[13] == c_8_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[13] == c_8_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[14] == c_8_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[14] == c_8_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[15] == c_8_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[15] == c_8_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[16] == c_8_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[16] == c_8_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[17] == c_8_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[17] == c_8_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[18] == c_8_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[18] == c_8_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[19] == c_8_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[19] == c_8_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[20] == c_8_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[20] == c_8_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[21] == c_8_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[21] == c_8_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[22] == c_8_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[22] == c_8_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[23] == c_8_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[23] == c_8_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[24] == c_8_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[24] == c_8_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[25] == c_8_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[25] == c_8_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[26] == c_8_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[26] == c_8_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[27] == c_8_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[27] == c_8_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[28] == c_8_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[28] == c_8_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[29] == c_8_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[29] == c_8_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[30] == c_8_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[30] == c_8_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[31] == c_8_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[31] == c_8_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_8[32] == c_8_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_8[32] == c_8_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[0] == c_9_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[0] == c_9_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[1] == c_9_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[1] == c_9_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[2] == c_9_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[2] == c_9_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[3] == c_9_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[3] == c_9_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[4] == c_9_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[4] == c_9_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[5] == c_9_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[5] == c_9_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[6] == c_9_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[6] == c_9_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[7] == c_9_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[7] == c_9_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[8] == c_9_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[8] == c_9_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[9] == c_9_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[9] == c_9_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[10] == c_9_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[10] == c_9_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[11] == c_9_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[11] == c_9_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[12] == c_9_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[12] == c_9_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[13] == c_9_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[13] == c_9_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[14] == c_9_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[14] == c_9_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[15] == c_9_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[15] == c_9_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[16] == c_9_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[16] == c_9_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[17] == c_9_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[17] == c_9_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[18] == c_9_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[18] == c_9_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[19] == c_9_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[19] == c_9_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[20] == c_9_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[20] == c_9_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[21] == c_9_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[21] == c_9_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[22] == c_9_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[22] == c_9_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[23] == c_9_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[23] == c_9_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[24] == c_9_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[24] == c_9_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[25] == c_9_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[25] == c_9_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[26] == c_9_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[26] == c_9_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[27] == c_9_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[27] == c_9_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[28] == c_9_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[28] == c_9_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[29] == c_9_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[29] == c_9_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[30] == c_9_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[30] == c_9_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[31] == c_9_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[31] == c_9_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_9[32] == c_9_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_9[32] == c_9_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[0] == c_10_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[0] == c_10_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[1] == c_10_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[1] == c_10_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[2] == c_10_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[2] == c_10_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[3] == c_10_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[3] == c_10_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[4] == c_10_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[4] == c_10_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[5] == c_10_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[5] == c_10_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[6] == c_10_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[6] == c_10_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[7] == c_10_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[7] == c_10_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[8] == c_10_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[8] == c_10_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[9] == c_10_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[9] == c_10_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[10] == c_10_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[10] == c_10_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[11] == c_10_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[11] == c_10_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[12] == c_10_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[12] == c_10_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[13] == c_10_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[13] == c_10_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[14] == c_10_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[14] == c_10_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[15] == c_10_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[15] == c_10_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[16] == c_10_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[16] == c_10_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[17] == c_10_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[17] == c_10_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[18] == c_10_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[18] == c_10_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[19] == c_10_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[19] == c_10_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[20] == c_10_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[20] == c_10_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[21] == c_10_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[21] == c_10_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[22] == c_10_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[22] == c_10_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[23] == c_10_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[23] == c_10_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[24] == c_10_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[24] == c_10_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[25] == c_10_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[25] == c_10_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[26] == c_10_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[26] == c_10_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[27] == c_10_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[27] == c_10_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[28] == c_10_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[28] == c_10_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[29] == c_10_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[29] == c_10_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[30] == c_10_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[30] == c_10_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[31] == c_10_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[31] == c_10_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_10[32] == c_10_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_10[32] == c_10_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[0] == c_11_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[0] == c_11_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[1] == c_11_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[1] == c_11_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[2] == c_11_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[2] == c_11_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[3] == c_11_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[3] == c_11_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[4] == c_11_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[4] == c_11_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[5] == c_11_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[5] == c_11_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[6] == c_11_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[6] == c_11_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[7] == c_11_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[7] == c_11_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[8] == c_11_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[8] == c_11_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[9] == c_11_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[9] == c_11_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[10] == c_11_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[10] == c_11_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[11] == c_11_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[11] == c_11_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[12] == c_11_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[12] == c_11_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[13] == c_11_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[13] == c_11_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[14] == c_11_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[14] == c_11_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[15] == c_11_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[15] == c_11_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[16] == c_11_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[16] == c_11_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[17] == c_11_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[17] == c_11_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[18] == c_11_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[18] == c_11_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[19] == c_11_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[19] == c_11_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[20] == c_11_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[20] == c_11_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[21] == c_11_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[21] == c_11_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[22] == c_11_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[22] == c_11_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[23] == c_11_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[23] == c_11_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[24] == c_11_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[24] == c_11_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[25] == c_11_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[25] == c_11_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[26] == c_11_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[26] == c_11_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[27] == c_11_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[27] == c_11_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[28] == c_11_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[28] == c_11_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[29] == c_11_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[29] == c_11_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[30] == c_11_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[30] == c_11_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[31] == c_11_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[31] == c_11_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_11[32] == c_11_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_11[32] == c_11_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[0] == c_12_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[0] == c_12_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[1] == c_12_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[1] == c_12_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[2] == c_12_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[2] == c_12_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[3] == c_12_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[3] == c_12_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[4] == c_12_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[4] == c_12_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[5] == c_12_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[5] == c_12_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[6] == c_12_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[6] == c_12_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[7] == c_12_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[7] == c_12_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[8] == c_12_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[8] == c_12_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[9] == c_12_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[9] == c_12_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[10] == c_12_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[10] == c_12_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[11] == c_12_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[11] == c_12_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[12] == c_12_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[12] == c_12_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[13] == c_12_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[13] == c_12_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[14] == c_12_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[14] == c_12_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[15] == c_12_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[15] == c_12_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[16] == c_12_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[16] == c_12_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[17] == c_12_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[17] == c_12_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[18] == c_12_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[18] == c_12_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[19] == c_12_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[19] == c_12_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[20] == c_12_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[20] == c_12_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[21] == c_12_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[21] == c_12_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[22] == c_12_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[22] == c_12_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[23] == c_12_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[23] == c_12_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[24] == c_12_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[24] == c_12_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[25] == c_12_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[25] == c_12_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[26] == c_12_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[26] == c_12_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[27] == c_12_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[27] == c_12_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[28] == c_12_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[28] == c_12_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[29] == c_12_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[29] == c_12_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[30] == c_12_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[30] == c_12_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[31] == c_12_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[31] == c_12_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_12[32] == c_12_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_12[32] == c_12_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[0] == c_13_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[0] == c_13_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[1] == c_13_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[1] == c_13_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[2] == c_13_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[2] == c_13_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[3] == c_13_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[3] == c_13_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[4] == c_13_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[4] == c_13_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[5] == c_13_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[5] == c_13_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[6] == c_13_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[6] == c_13_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[7] == c_13_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[7] == c_13_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[8] == c_13_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[8] == c_13_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[9] == c_13_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[9] == c_13_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[10] == c_13_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[10] == c_13_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[11] == c_13_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[11] == c_13_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[12] == c_13_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[12] == c_13_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[13] == c_13_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[13] == c_13_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[14] == c_13_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[14] == c_13_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[15] == c_13_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[15] == c_13_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[16] == c_13_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[16] == c_13_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[17] == c_13_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[17] == c_13_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[18] == c_13_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[18] == c_13_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[19] == c_13_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[19] == c_13_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[20] == c_13_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[20] == c_13_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[21] == c_13_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[21] == c_13_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[22] == c_13_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[22] == c_13_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[23] == c_13_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[23] == c_13_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[24] == c_13_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[24] == c_13_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[25] == c_13_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[25] == c_13_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[26] == c_13_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[26] == c_13_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[27] == c_13_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[27] == c_13_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[28] == c_13_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[28] == c_13_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[29] == c_13_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[29] == c_13_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[30] == c_13_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[30] == c_13_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[31] == c_13_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[31] == c_13_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_13[32] == c_13_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_13[32] == c_13_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[0] == c_14_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[0] == c_14_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[1] == c_14_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[1] == c_14_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[2] == c_14_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[2] == c_14_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[3] == c_14_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[3] == c_14_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[4] == c_14_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[4] == c_14_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[5] == c_14_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[5] == c_14_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[6] == c_14_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[6] == c_14_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[7] == c_14_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[7] == c_14_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[8] == c_14_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[8] == c_14_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[9] == c_14_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[9] == c_14_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[10] == c_14_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[10] == c_14_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[11] == c_14_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[11] == c_14_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[12] == c_14_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[12] == c_14_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[13] == c_14_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[13] == c_14_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[14] == c_14_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[14] == c_14_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[15] == c_14_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[15] == c_14_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[16] == c_14_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[16] == c_14_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[17] == c_14_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[17] == c_14_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[18] == c_14_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[18] == c_14_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[19] == c_14_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[19] == c_14_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[20] == c_14_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[20] == c_14_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[21] == c_14_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[21] == c_14_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[22] == c_14_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[22] == c_14_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[23] == c_14_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[23] == c_14_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[24] == c_14_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[24] == c_14_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[25] == c_14_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[25] == c_14_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[26] == c_14_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[26] == c_14_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[27] == c_14_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[27] == c_14_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[28] == c_14_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[28] == c_14_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[29] == c_14_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[29] == c_14_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[30] == c_14_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[30] == c_14_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[31] == c_14_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[31] == c_14_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_14[32] == c_14_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_14[32] == c_14_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[0] == c_15_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[0] == c_15_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[1] == c_15_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[1] == c_15_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[2] == c_15_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[2] == c_15_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[3] == c_15_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[3] == c_15_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[4] == c_15_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[4] == c_15_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[5] == c_15_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[5] == c_15_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[6] == c_15_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[6] == c_15_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[7] == c_15_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[7] == c_15_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[8] == c_15_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[8] == c_15_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[9] == c_15_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[9] == c_15_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[10] == c_15_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[10] == c_15_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[11] == c_15_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[11] == c_15_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[12] == c_15_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[12] == c_15_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[13] == c_15_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[13] == c_15_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[14] == c_15_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[14] == c_15_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[15] == c_15_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[15] == c_15_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[16] == c_15_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[16] == c_15_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[17] == c_15_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[17] == c_15_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[18] == c_15_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[18] == c_15_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[19] == c_15_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[19] == c_15_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[20] == c_15_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[20] == c_15_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[21] == c_15_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[21] == c_15_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[22] == c_15_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[22] == c_15_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[23] == c_15_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[23] == c_15_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[24] == c_15_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[24] == c_15_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[25] == c_15_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[25] == c_15_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[26] == c_15_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[26] == c_15_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[27] == c_15_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[27] == c_15_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[28] == c_15_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[28] == c_15_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[29] == c_15_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[29] == c_15_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[30] == c_15_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[30] == c_15_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[31] == c_15_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[31] == c_15_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_15[32] == c_15_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_15[32] == c_15_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[0] == c_16_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[0] == c_16_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[1] == c_16_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[1] == c_16_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[2] == c_16_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[2] == c_16_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[3] == c_16_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[3] == c_16_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[4] == c_16_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[4] == c_16_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[5] == c_16_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[5] == c_16_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[6] == c_16_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[6] == c_16_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[7] == c_16_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[7] == c_16_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[8] == c_16_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[8] == c_16_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[9] == c_16_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[9] == c_16_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[10] == c_16_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[10] == c_16_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[11] == c_16_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[11] == c_16_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[12] == c_16_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[12] == c_16_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[13] == c_16_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[13] == c_16_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[14] == c_16_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[14] == c_16_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[15] == c_16_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[15] == c_16_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[16] == c_16_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[16] == c_16_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[17] == c_16_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[17] == c_16_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[18] == c_16_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[18] == c_16_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[19] == c_16_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[19] == c_16_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[20] == c_16_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[20] == c_16_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[21] == c_16_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[21] == c_16_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[22] == c_16_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[22] == c_16_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[23] == c_16_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[23] == c_16_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[24] == c_16_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[24] == c_16_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[25] == c_16_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[25] == c_16_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[26] == c_16_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[26] == c_16_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[27] == c_16_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[27] == c_16_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[28] == c_16_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[28] == c_16_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[29] == c_16_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[29] == c_16_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[30] == c_16_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[30] == c_16_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[31] == c_16_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[31] == c_16_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_16[32] == c_16_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_16[32] == c_16_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[0] == c_17_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[0] == c_17_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[1] == c_17_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[1] == c_17_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[2] == c_17_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[2] == c_17_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[3] == c_17_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[3] == c_17_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[4] == c_17_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[4] == c_17_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[5] == c_17_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[5] == c_17_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[6] == c_17_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[6] == c_17_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[7] == c_17_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[7] == c_17_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[8] == c_17_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[8] == c_17_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[9] == c_17_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[9] == c_17_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[10] == c_17_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[10] == c_17_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[11] == c_17_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[11] == c_17_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[12] == c_17_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[12] == c_17_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[13] == c_17_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[13] == c_17_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[14] == c_17_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[14] == c_17_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[15] == c_17_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[15] == c_17_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[16] == c_17_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[16] == c_17_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[17] == c_17_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[17] == c_17_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[18] == c_17_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[18] == c_17_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[19] == c_17_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[19] == c_17_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[20] == c_17_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[20] == c_17_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[21] == c_17_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[21] == c_17_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[22] == c_17_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[22] == c_17_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[23] == c_17_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[23] == c_17_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[24] == c_17_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[24] == c_17_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[25] == c_17_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[25] == c_17_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[26] == c_17_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[26] == c_17_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[27] == c_17_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[27] == c_17_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[28] == c_17_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[28] == c_17_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[29] == c_17_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[29] == c_17_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[30] == c_17_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[30] == c_17_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[31] == c_17_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[31] == c_17_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_17[32] == c_17_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_17[32] == c_17_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[0] == c_18_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[0] == c_18_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[1] == c_18_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[1] == c_18_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[2] == c_18_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[2] == c_18_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[3] == c_18_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[3] == c_18_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[4] == c_18_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[4] == c_18_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[5] == c_18_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[5] == c_18_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[6] == c_18_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[6] == c_18_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[7] == c_18_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[7] == c_18_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[8] == c_18_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[8] == c_18_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[9] == c_18_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[9] == c_18_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[10] == c_18_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[10] == c_18_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[11] == c_18_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[11] == c_18_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[12] == c_18_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[12] == c_18_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[13] == c_18_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[13] == c_18_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[14] == c_18_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[14] == c_18_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[15] == c_18_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[15] == c_18_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[16] == c_18_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[16] == c_18_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[17] == c_18_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[17] == c_18_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[18] == c_18_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[18] == c_18_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[19] == c_18_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[19] == c_18_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[20] == c_18_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[20] == c_18_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[21] == c_18_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[21] == c_18_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[22] == c_18_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[22] == c_18_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[23] == c_18_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[23] == c_18_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[24] == c_18_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[24] == c_18_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[25] == c_18_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[25] == c_18_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[26] == c_18_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[26] == c_18_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[27] == c_18_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[27] == c_18_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[28] == c_18_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[28] == c_18_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[29] == c_18_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[29] == c_18_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[30] == c_18_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[30] == c_18_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[31] == c_18_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[31] == c_18_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_18[32] == c_18_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_18[32] == c_18_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[0] == c_19_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[0] == c_19_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[1] == c_19_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[1] == c_19_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[2] == c_19_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[2] == c_19_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[3] == c_19_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[3] == c_19_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[4] == c_19_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[4] == c_19_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[5] == c_19_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[5] == c_19_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[6] == c_19_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[6] == c_19_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[7] == c_19_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[7] == c_19_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[8] == c_19_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[8] == c_19_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[9] == c_19_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[9] == c_19_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[10] == c_19_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[10] == c_19_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[11] == c_19_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[11] == c_19_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[12] == c_19_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[12] == c_19_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[13] == c_19_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[13] == c_19_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[14] == c_19_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[14] == c_19_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[15] == c_19_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[15] == c_19_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[16] == c_19_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[16] == c_19_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[17] == c_19_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[17] == c_19_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[18] == c_19_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[18] == c_19_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[19] == c_19_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[19] == c_19_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[20] == c_19_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[20] == c_19_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[21] == c_19_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[21] == c_19_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[22] == c_19_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[22] == c_19_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[23] == c_19_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[23] == c_19_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[24] == c_19_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[24] == c_19_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[25] == c_19_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[25] == c_19_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[26] == c_19_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[26] == c_19_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[27] == c_19_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[27] == c_19_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[28] == c_19_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[28] == c_19_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[29] == c_19_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[29] == c_19_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[30] == c_19_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[30] == c_19_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[31] == c_19_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[31] == c_19_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_19[32] == c_19_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_19[32] == c_19_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[0] == c_20_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[0] == c_20_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[1] == c_20_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[1] == c_20_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[2] == c_20_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[2] == c_20_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[3] == c_20_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[3] == c_20_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[4] == c_20_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[4] == c_20_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[5] == c_20_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[5] == c_20_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[6] == c_20_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[6] == c_20_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[7] == c_20_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[7] == c_20_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[8] == c_20_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[8] == c_20_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[9] == c_20_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[9] == c_20_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[10] == c_20_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[10] == c_20_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[11] == c_20_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[11] == c_20_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[12] == c_20_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[12] == c_20_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[13] == c_20_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[13] == c_20_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[14] == c_20_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[14] == c_20_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[15] == c_20_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[15] == c_20_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[16] == c_20_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[16] == c_20_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[17] == c_20_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[17] == c_20_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[18] == c_20_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[18] == c_20_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[19] == c_20_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[19] == c_20_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[20] == c_20_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[20] == c_20_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[21] == c_20_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[21] == c_20_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[22] == c_20_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[22] == c_20_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[23] == c_20_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[23] == c_20_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[24] == c_20_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[24] == c_20_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[25] == c_20_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[25] == c_20_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[26] == c_20_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[26] == c_20_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[27] == c_20_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[27] == c_20_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[28] == c_20_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[28] == c_20_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[29] == c_20_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[29] == c_20_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[30] == c_20_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[30] == c_20_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[31] == c_20_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[31] == c_20_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_20[32] == c_20_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_20[32] == c_20_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[0] == c_21_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[0] == c_21_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[1] == c_21_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[1] == c_21_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[2] == c_21_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[2] == c_21_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[3] == c_21_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[3] == c_21_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[4] == c_21_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[4] == c_21_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[5] == c_21_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[5] == c_21_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[6] == c_21_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[6] == c_21_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[7] == c_21_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[7] == c_21_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[8] == c_21_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[8] == c_21_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[9] == c_21_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[9] == c_21_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[10] == c_21_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[10] == c_21_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[11] == c_21_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[11] == c_21_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[12] == c_21_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[12] == c_21_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[13] == c_21_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[13] == c_21_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[14] == c_21_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[14] == c_21_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[15] == c_21_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[15] == c_21_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[16] == c_21_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[16] == c_21_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[17] == c_21_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[17] == c_21_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[18] == c_21_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[18] == c_21_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[19] == c_21_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[19] == c_21_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[20] == c_21_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[20] == c_21_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[21] == c_21_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[21] == c_21_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[22] == c_21_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[22] == c_21_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[23] == c_21_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[23] == c_21_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[24] == c_21_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[24] == c_21_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[25] == c_21_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[25] == c_21_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[26] == c_21_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[26] == c_21_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[27] == c_21_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[27] == c_21_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[28] == c_21_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[28] == c_21_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[29] == c_21_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[29] == c_21_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[30] == c_21_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[30] == c_21_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[31] == c_21_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[31] == c_21_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_21[32] == c_21_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_21[32] == c_21_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[0] == c_22_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[0] == c_22_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[1] == c_22_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[1] == c_22_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[2] == c_22_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[2] == c_22_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[3] == c_22_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[3] == c_22_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[4] == c_22_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[4] == c_22_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[5] == c_22_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[5] == c_22_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[6] == c_22_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[6] == c_22_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[7] == c_22_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[7] == c_22_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[8] == c_22_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[8] == c_22_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[9] == c_22_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[9] == c_22_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[10] == c_22_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[10] == c_22_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[11] == c_22_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[11] == c_22_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[12] == c_22_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[12] == c_22_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[13] == c_22_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[13] == c_22_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[14] == c_22_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[14] == c_22_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[15] == c_22_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[15] == c_22_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[16] == c_22_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[16] == c_22_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[17] == c_22_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[17] == c_22_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[18] == c_22_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[18] == c_22_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[19] == c_22_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[19] == c_22_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[20] == c_22_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[20] == c_22_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[21] == c_22_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[21] == c_22_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[22] == c_22_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[22] == c_22_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[23] == c_22_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[23] == c_22_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[24] == c_22_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[24] == c_22_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[25] == c_22_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[25] == c_22_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[26] == c_22_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[26] == c_22_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[27] == c_22_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[27] == c_22_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[28] == c_22_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[28] == c_22_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[29] == c_22_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[29] == c_22_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[30] == c_22_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[30] == c_22_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[31] == c_22_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[31] == c_22_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_22[32] == c_22_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_22[32] == c_22_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[0] == c_23_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[0] == c_23_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[1] == c_23_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[1] == c_23_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[2] == c_23_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[2] == c_23_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[3] == c_23_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[3] == c_23_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[4] == c_23_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[4] == c_23_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[5] == c_23_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[5] == c_23_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[6] == c_23_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[6] == c_23_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[7] == c_23_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[7] == c_23_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[8] == c_23_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[8] == c_23_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[9] == c_23_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[9] == c_23_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[10] == c_23_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[10] == c_23_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[11] == c_23_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[11] == c_23_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[12] == c_23_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[12] == c_23_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[13] == c_23_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[13] == c_23_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[14] == c_23_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[14] == c_23_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[15] == c_23_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[15] == c_23_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[16] == c_23_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[16] == c_23_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[17] == c_23_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[17] == c_23_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[18] == c_23_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[18] == c_23_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[19] == c_23_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[19] == c_23_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[20] == c_23_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[20] == c_23_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[21] == c_23_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[21] == c_23_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[22] == c_23_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[22] == c_23_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[23] == c_23_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[23] == c_23_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[24] == c_23_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[24] == c_23_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[25] == c_23_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[25] == c_23_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[26] == c_23_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[26] == c_23_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[27] == c_23_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[27] == c_23_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[28] == c_23_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[28] == c_23_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[29] == c_23_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[29] == c_23_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[30] == c_23_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[30] == c_23_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[31] == c_23_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[31] == c_23_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_23[32] == c_23_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_23[32] == c_23_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[0] == c_24_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[0] == c_24_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[1] == c_24_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[1] == c_24_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[2] == c_24_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[2] == c_24_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[3] == c_24_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[3] == c_24_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[4] == c_24_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[4] == c_24_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[5] == c_24_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[5] == c_24_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[6] == c_24_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[6] == c_24_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[7] == c_24_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[7] == c_24_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[8] == c_24_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[8] == c_24_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[9] == c_24_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[9] == c_24_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[10] == c_24_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[10] == c_24_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[11] == c_24_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[11] == c_24_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[12] == c_24_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[12] == c_24_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[13] == c_24_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[13] == c_24_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[14] == c_24_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[14] == c_24_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[15] == c_24_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[15] == c_24_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[16] == c_24_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[16] == c_24_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[17] == c_24_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[17] == c_24_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[18] == c_24_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[18] == c_24_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[19] == c_24_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[19] == c_24_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[20] == c_24_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[20] == c_24_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[21] == c_24_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[21] == c_24_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[22] == c_24_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[22] == c_24_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[23] == c_24_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[23] == c_24_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[24] == c_24_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[24] == c_24_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[25] == c_24_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[25] == c_24_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[26] == c_24_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[26] == c_24_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[27] == c_24_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[27] == c_24_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[28] == c_24_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[28] == c_24_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[29] == c_24_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[29] == c_24_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[30] == c_24_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[30] == c_24_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[31] == c_24_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[31] == c_24_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_24[32] == c_24_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_24[32] == c_24_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[0] == c_25_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[0] == c_25_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[1] == c_25_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[1] == c_25_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[2] == c_25_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[2] == c_25_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[3] == c_25_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[3] == c_25_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[4] == c_25_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[4] == c_25_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[5] == c_25_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[5] == c_25_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[6] == c_25_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[6] == c_25_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[7] == c_25_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[7] == c_25_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[8] == c_25_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[8] == c_25_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[9] == c_25_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[9] == c_25_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[10] == c_25_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[10] == c_25_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[11] == c_25_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[11] == c_25_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[12] == c_25_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[12] == c_25_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[13] == c_25_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[13] == c_25_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[14] == c_25_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[14] == c_25_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[15] == c_25_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[15] == c_25_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[16] == c_25_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[16] == c_25_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[17] == c_25_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[17] == c_25_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[18] == c_25_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[18] == c_25_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[19] == c_25_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[19] == c_25_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[20] == c_25_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[20] == c_25_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[21] == c_25_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[21] == c_25_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[22] == c_25_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[22] == c_25_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[23] == c_25_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[23] == c_25_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[24] == c_25_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[24] == c_25_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[25] == c_25_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[25] == c_25_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[26] == c_25_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[26] == c_25_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[27] == c_25_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[27] == c_25_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[28] == c_25_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[28] == c_25_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[29] == c_25_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[29] == c_25_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[30] == c_25_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[30] == c_25_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[31] == c_25_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[31] == c_25_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_25[32] == c_25_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_25[32] == c_25_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[0] == c_26_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[0] == c_26_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[1] == c_26_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[1] == c_26_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[2] == c_26_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[2] == c_26_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[3] == c_26_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[3] == c_26_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[4] == c_26_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[4] == c_26_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[5] == c_26_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[5] == c_26_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[6] == c_26_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[6] == c_26_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[7] == c_26_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[7] == c_26_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[8] == c_26_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[8] == c_26_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[9] == c_26_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[9] == c_26_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[10] == c_26_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[10] == c_26_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[11] == c_26_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[11] == c_26_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[12] == c_26_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[12] == c_26_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[13] == c_26_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[13] == c_26_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[14] == c_26_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[14] == c_26_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[15] == c_26_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[15] == c_26_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[16] == c_26_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[16] == c_26_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[17] == c_26_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[17] == c_26_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[18] == c_26_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[18] == c_26_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[19] == c_26_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[19] == c_26_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[20] == c_26_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[20] == c_26_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[21] == c_26_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[21] == c_26_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[22] == c_26_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[22] == c_26_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[23] == c_26_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[23] == c_26_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[24] == c_26_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[24] == c_26_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[25] == c_26_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[25] == c_26_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[26] == c_26_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[26] == c_26_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[27] == c_26_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[27] == c_26_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[28] == c_26_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[28] == c_26_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[29] == c_26_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[29] == c_26_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[30] == c_26_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[30] == c_26_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[31] == c_26_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[31] == c_26_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_26[32] == c_26_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_26[32] == c_26_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[0] == c_27_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[0] == c_27_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[1] == c_27_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[1] == c_27_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[2] == c_27_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[2] == c_27_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[3] == c_27_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[3] == c_27_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[4] == c_27_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[4] == c_27_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[5] == c_27_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[5] == c_27_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[6] == c_27_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[6] == c_27_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[7] == c_27_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[7] == c_27_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[8] == c_27_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[8] == c_27_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[9] == c_27_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[9] == c_27_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[10] == c_27_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[10] == c_27_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[11] == c_27_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[11] == c_27_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[12] == c_27_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[12] == c_27_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[13] == c_27_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[13] == c_27_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[14] == c_27_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[14] == c_27_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[15] == c_27_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[15] == c_27_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[16] == c_27_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[16] == c_27_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[17] == c_27_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[17] == c_27_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[18] == c_27_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[18] == c_27_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[19] == c_27_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[19] == c_27_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[20] == c_27_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[20] == c_27_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[21] == c_27_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[21] == c_27_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[22] == c_27_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[22] == c_27_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[23] == c_27_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[23] == c_27_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[24] == c_27_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[24] == c_27_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[25] == c_27_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[25] == c_27_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[26] == c_27_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[26] == c_27_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[27] == c_27_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[27] == c_27_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[28] == c_27_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[28] == c_27_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[29] == c_27_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[29] == c_27_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[30] == c_27_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[30] == c_27_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[31] == c_27_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[31] == c_27_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_27[32] == c_27_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_27[32] == c_27_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[0] == c_28_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[0] == c_28_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[1] == c_28_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[1] == c_28_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[2] == c_28_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[2] == c_28_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[3] == c_28_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[3] == c_28_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[4] == c_28_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[4] == c_28_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[5] == c_28_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[5] == c_28_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[6] == c_28_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[6] == c_28_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[7] == c_28_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[7] == c_28_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[8] == c_28_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[8] == c_28_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[9] == c_28_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[9] == c_28_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[10] == c_28_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[10] == c_28_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[11] == c_28_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[11] == c_28_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[12] == c_28_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[12] == c_28_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[13] == c_28_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[13] == c_28_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[14] == c_28_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[14] == c_28_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[15] == c_28_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[15] == c_28_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[16] == c_28_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[16] == c_28_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[17] == c_28_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[17] == c_28_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[18] == c_28_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[18] == c_28_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[19] == c_28_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[19] == c_28_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[20] == c_28_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[20] == c_28_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[21] == c_28_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[21] == c_28_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[22] == c_28_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[22] == c_28_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[23] == c_28_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[23] == c_28_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[24] == c_28_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[24] == c_28_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[25] == c_28_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[25] == c_28_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[26] == c_28_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[26] == c_28_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[27] == c_28_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[27] == c_28_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[28] == c_28_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[28] == c_28_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[29] == c_28_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[29] == c_28_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[30] == c_28_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[30] == c_28_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[31] == c_28_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[31] == c_28_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_28[32] == c_28_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_28[32] == c_28_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[0] == c_29_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[0] == c_29_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[1] == c_29_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[1] == c_29_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[2] == c_29_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[2] == c_29_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[3] == c_29_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[3] == c_29_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[4] == c_29_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[4] == c_29_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[5] == c_29_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[5] == c_29_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[6] == c_29_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[6] == c_29_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[7] == c_29_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[7] == c_29_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[8] == c_29_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[8] == c_29_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[9] == c_29_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[9] == c_29_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[10] == c_29_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[10] == c_29_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[11] == c_29_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[11] == c_29_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[12] == c_29_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[12] == c_29_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[13] == c_29_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[13] == c_29_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[14] == c_29_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[14] == c_29_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[15] == c_29_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[15] == c_29_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[16] == c_29_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[16] == c_29_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[17] == c_29_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[17] == c_29_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[18] == c_29_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[18] == c_29_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[19] == c_29_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[19] == c_29_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[20] == c_29_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[20] == c_29_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[21] == c_29_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[21] == c_29_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[22] == c_29_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[22] == c_29_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[23] == c_29_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[23] == c_29_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[24] == c_29_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[24] == c_29_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[25] == c_29_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[25] == c_29_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[26] == c_29_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[26] == c_29_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[27] == c_29_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[27] == c_29_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[28] == c_29_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[28] == c_29_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[29] == c_29_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[29] == c_29_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[30] == c_29_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[30] == c_29_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[31] == c_29_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[31] == c_29_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_29[32] == c_29_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_29[32] == c_29_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[0] == c_30_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[0] == c_30_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[1] == c_30_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[1] == c_30_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[2] == c_30_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[2] == c_30_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[3] == c_30_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[3] == c_30_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[4] == c_30_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[4] == c_30_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[5] == c_30_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[5] == c_30_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[6] == c_30_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[6] == c_30_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[7] == c_30_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[7] == c_30_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[8] == c_30_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[8] == c_30_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[9] == c_30_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[9] == c_30_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[10] == c_30_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[10] == c_30_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[11] == c_30_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[11] == c_30_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[12] == c_30_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[12] == c_30_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[13] == c_30_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[13] == c_30_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[14] == c_30_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[14] == c_30_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[15] == c_30_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[15] == c_30_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[16] == c_30_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[16] == c_30_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[17] == c_30_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[17] == c_30_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[18] == c_30_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[18] == c_30_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[19] == c_30_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[19] == c_30_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[20] == c_30_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[20] == c_30_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[21] == c_30_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[21] == c_30_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[22] == c_30_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[22] == c_30_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[23] == c_30_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[23] == c_30_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[24] == c_30_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[24] == c_30_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[25] == c_30_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[25] == c_30_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[26] == c_30_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[26] == c_30_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[27] == c_30_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[27] == c_30_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[28] == c_30_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[28] == c_30_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[29] == c_30_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[29] == c_30_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[30] == c_30_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[30] == c_30_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[31] == c_30_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[31] == c_30_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_30[32] == c_30_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_30[32] == c_30_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[0] == c_31_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[0] == c_31_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[1] == c_31_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[1] == c_31_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[2] == c_31_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[2] == c_31_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[3] == c_31_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[3] == c_31_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[4] == c_31_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[4] == c_31_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[5] == c_31_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[5] == c_31_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[6] == c_31_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[6] == c_31_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[7] == c_31_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[7] == c_31_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[8] == c_31_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[8] == c_31_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[9] == c_31_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[9] == c_31_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[10] == c_31_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[10] == c_31_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[11] == c_31_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[11] == c_31_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[12] == c_31_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[12] == c_31_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[13] == c_31_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[13] == c_31_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[14] == c_31_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[14] == c_31_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[15] == c_31_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[15] == c_31_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[16] == c_31_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[16] == c_31_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[17] == c_31_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[17] == c_31_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[18] == c_31_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[18] == c_31_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[19] == c_31_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[19] == c_31_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[20] == c_31_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[20] == c_31_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[21] == c_31_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[21] == c_31_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[22] == c_31_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[22] == c_31_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[23] == c_31_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[23] == c_31_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[24] == c_31_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[24] == c_31_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[25] == c_31_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[25] == c_31_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[26] == c_31_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[26] == c_31_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[27] == c_31_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[27] == c_31_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[28] == c_31_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[28] == c_31_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[29] == c_31_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[29] == c_31_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[30] == c_31_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[30] == c_31_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[31] == c_31_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[31] == c_31_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_31[32] == c_31_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_31[32] == c_31_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[0] == c_32_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[0] == c_32_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[1] == c_32_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[1] == c_32_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[2] == c_32_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[2] == c_32_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[3] == c_32_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[3] == c_32_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[4] == c_32_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[4] == c_32_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[5] == c_32_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[5] == c_32_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[6] == c_32_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[6] == c_32_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[7] == c_32_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[7] == c_32_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[8] == c_32_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[8] == c_32_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[9] == c_32_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[9] == c_32_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[10] == c_32_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[10] == c_32_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[11] == c_32_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[11] == c_32_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[12] == c_32_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[12] == c_32_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[13] == c_32_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[13] == c_32_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[14] == c_32_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[14] == c_32_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[15] == c_32_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[15] == c_32_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[16] == c_32_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[16] == c_32_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[17] == c_32_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[17] == c_32_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[18] == c_32_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[18] == c_32_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[19] == c_32_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[19] == c_32_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[20] == c_32_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[20] == c_32_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[21] == c_32_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[21] == c_32_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[22] == c_32_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[22] == c_32_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[23] == c_32_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[23] == c_32_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[24] == c_32_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[24] == c_32_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[25] == c_32_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[25] == c_32_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[26] == c_32_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[26] == c_32_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[27] == c_32_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[27] == c_32_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[28] == c_32_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[28] == c_32_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[29] == c_32_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[29] == c_32_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[30] == c_32_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[30] == c_32_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[31] == c_32_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[31] == c_32_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_32[32] == c_32_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_32[32] == c_32_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[0] == c_33_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[0] == c_33_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[1] == c_33_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[1] == c_33_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[2] == c_33_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[2] == c_33_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[3] == c_33_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[3] == c_33_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[4] == c_33_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[4] == c_33_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[5] == c_33_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[5] == c_33_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[6] == c_33_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[6] == c_33_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[7] == c_33_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[7] == c_33_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[8] == c_33_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[8] == c_33_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[9] == c_33_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[9] == c_33_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[10] == c_33_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[10] == c_33_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[11] == c_33_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[11] == c_33_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[12] == c_33_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[12] == c_33_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[13] == c_33_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[13] == c_33_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[14] == c_33_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[14] == c_33_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[15] == c_33_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[15] == c_33_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[16] == c_33_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[16] == c_33_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[17] == c_33_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[17] == c_33_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[18] == c_33_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[18] == c_33_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[19] == c_33_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[19] == c_33_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[20] == c_33_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[20] == c_33_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[21] == c_33_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[21] == c_33_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[22] == c_33_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[22] == c_33_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[23] == c_33_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[23] == c_33_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[24] == c_33_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[24] == c_33_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[25] == c_33_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[25] == c_33_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[26] == c_33_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[26] == c_33_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[27] == c_33_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[27] == c_33_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[28] == c_33_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[28] == c_33_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[29] == c_33_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[29] == c_33_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[30] == c_33_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[30] == c_33_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[31] == c_33_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[31] == c_33_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_33[32] == c_33_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_33[32] == c_33_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[0] == c_34_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[0] == c_34_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[1] == c_34_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[1] == c_34_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[2] == c_34_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[2] == c_34_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[3] == c_34_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[3] == c_34_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[4] == c_34_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[4] == c_34_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[5] == c_34_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[5] == c_34_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[6] == c_34_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[6] == c_34_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[7] == c_34_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[7] == c_34_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[8] == c_34_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[8] == c_34_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[9] == c_34_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[9] == c_34_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[10] == c_34_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[10] == c_34_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[11] == c_34_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[11] == c_34_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[12] == c_34_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[12] == c_34_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[13] == c_34_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[13] == c_34_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[14] == c_34_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[14] == c_34_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[15] == c_34_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[15] == c_34_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[16] == c_34_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[16] == c_34_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[17] == c_34_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[17] == c_34_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[18] == c_34_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[18] == c_34_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[19] == c_34_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[19] == c_34_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[20] == c_34_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[20] == c_34_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[21] == c_34_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[21] == c_34_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[22] == c_34_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[22] == c_34_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[23] == c_34_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[23] == c_34_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[24] == c_34_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[24] == c_34_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[25] == c_34_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[25] == c_34_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[26] == c_34_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[26] == c_34_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[27] == c_34_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[27] == c_34_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[28] == c_34_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[28] == c_34_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[29] == c_34_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[29] == c_34_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[30] == c_34_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[30] == c_34_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[31] == c_34_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[31] == c_34_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_34[32] == c_34_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_34[32] == c_34_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[0] == c_35_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[0] == c_35_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[1] == c_35_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[1] == c_35_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[2] == c_35_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[2] == c_35_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[3] == c_35_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[3] == c_35_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[4] == c_35_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[4] == c_35_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[5] == c_35_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[5] == c_35_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[6] == c_35_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[6] == c_35_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[7] == c_35_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[7] == c_35_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[8] == c_35_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[8] == c_35_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[9] == c_35_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[9] == c_35_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[10] == c_35_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[10] == c_35_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[11] == c_35_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[11] == c_35_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[12] == c_35_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[12] == c_35_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[13] == c_35_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[13] == c_35_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[14] == c_35_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[14] == c_35_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[15] == c_35_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[15] == c_35_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[16] == c_35_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[16] == c_35_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[17] == c_35_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[17] == c_35_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[18] == c_35_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[18] == c_35_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[19] == c_35_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[19] == c_35_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[20] == c_35_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[20] == c_35_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[21] == c_35_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[21] == c_35_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[22] == c_35_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[22] == c_35_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[23] == c_35_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[23] == c_35_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[24] == c_35_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[24] == c_35_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[25] == c_35_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[25] == c_35_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[26] == c_35_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[26] == c_35_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[27] == c_35_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[27] == c_35_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[28] == c_35_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[28] == c_35_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[29] == c_35_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[29] == c_35_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[30] == c_35_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[30] == c_35_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[31] == c_35_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[31] == c_35_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_35[32] == c_35_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_35[32] == c_35_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[0] == c_36_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[0] == c_36_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[1] == c_36_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[1] == c_36_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[2] == c_36_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[2] == c_36_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[3] == c_36_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[3] == c_36_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[4] == c_36_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[4] == c_36_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[5] == c_36_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[5] == c_36_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[6] == c_36_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[6] == c_36_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[7] == c_36_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[7] == c_36_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[8] == c_36_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[8] == c_36_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[9] == c_36_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[9] == c_36_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[10] == c_36_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[10] == c_36_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[11] == c_36_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[11] == c_36_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[12] == c_36_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[12] == c_36_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[13] == c_36_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[13] == c_36_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[14] == c_36_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[14] == c_36_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[15] == c_36_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[15] == c_36_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[16] == c_36_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[16] == c_36_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[17] == c_36_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[17] == c_36_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[18] == c_36_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[18] == c_36_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[19] == c_36_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[19] == c_36_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[20] == c_36_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[20] == c_36_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[21] == c_36_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[21] == c_36_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[22] == c_36_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[22] == c_36_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[23] == c_36_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[23] == c_36_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[24] == c_36_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[24] == c_36_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[25] == c_36_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[25] == c_36_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[26] == c_36_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[26] == c_36_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[27] == c_36_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[27] == c_36_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[28] == c_36_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[28] == c_36_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[29] == c_36_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[29] == c_36_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[30] == c_36_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[30] == c_36_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[31] == c_36_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[31] == c_36_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_36[32] == c_36_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_36[32] == c_36_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[0] == c_37_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[0] == c_37_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[1] == c_37_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[1] == c_37_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[2] == c_37_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[2] == c_37_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[3] == c_37_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[3] == c_37_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[4] == c_37_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[4] == c_37_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[5] == c_37_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[5] == c_37_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[6] == c_37_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[6] == c_37_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[7] == c_37_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[7] == c_37_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[8] == c_37_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[8] == c_37_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[9] == c_37_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[9] == c_37_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[10] == c_37_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[10] == c_37_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[11] == c_37_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[11] == c_37_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[12] == c_37_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[12] == c_37_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[13] == c_37_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[13] == c_37_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[14] == c_37_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[14] == c_37_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[15] == c_37_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[15] == c_37_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[16] == c_37_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[16] == c_37_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[17] == c_37_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[17] == c_37_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[18] == c_37_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[18] == c_37_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[19] == c_37_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[19] == c_37_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[20] == c_37_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[20] == c_37_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[21] == c_37_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[21] == c_37_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[22] == c_37_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[22] == c_37_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[23] == c_37_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[23] == c_37_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[24] == c_37_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[24] == c_37_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[25] == c_37_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[25] == c_37_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[26] == c_37_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[26] == c_37_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[27] == c_37_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[27] == c_37_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[28] == c_37_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[28] == c_37_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[29] == c_37_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[29] == c_37_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[30] == c_37_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[30] == c_37_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[31] == c_37_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[31] == c_37_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_37[32] == c_37_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_37[32] == c_37_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[0] == c_38_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[0] == c_38_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[1] == c_38_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[1] == c_38_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[2] == c_38_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[2] == c_38_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[3] == c_38_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[3] == c_38_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[4] == c_38_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[4] == c_38_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[5] == c_38_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[5] == c_38_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[6] == c_38_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[6] == c_38_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[7] == c_38_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[7] == c_38_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[8] == c_38_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[8] == c_38_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[9] == c_38_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[9] == c_38_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[10] == c_38_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[10] == c_38_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[11] == c_38_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[11] == c_38_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[12] == c_38_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[12] == c_38_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[13] == c_38_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[13] == c_38_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[14] == c_38_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[14] == c_38_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[15] == c_38_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[15] == c_38_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[16] == c_38_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[16] == c_38_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[17] == c_38_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[17] == c_38_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[18] == c_38_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[18] == c_38_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[19] == c_38_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[19] == c_38_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[20] == c_38_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[20] == c_38_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[21] == c_38_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[21] == c_38_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[22] == c_38_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[22] == c_38_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[23] == c_38_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[23] == c_38_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[24] == c_38_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[24] == c_38_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[25] == c_38_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[25] == c_38_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[26] == c_38_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[26] == c_38_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[27] == c_38_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[27] == c_38_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[28] == c_38_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[28] == c_38_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[29] == c_38_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[29] == c_38_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[30] == c_38_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[30] == c_38_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[31] == c_38_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[31] == c_38_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_38[32] == c_38_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_38[32] == c_38_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[0] == c_39_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[0] == c_39_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[1] == c_39_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[1] == c_39_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[2] == c_39_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[2] == c_39_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[3] == c_39_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[3] == c_39_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[4] == c_39_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[4] == c_39_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[5] == c_39_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[5] == c_39_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[6] == c_39_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[6] == c_39_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[7] == c_39_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[7] == c_39_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[8] == c_39_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[8] == c_39_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[9] == c_39_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[9] == c_39_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[10] == c_39_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[10] == c_39_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[11] == c_39_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[11] == c_39_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[12] == c_39_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[12] == c_39_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[13] == c_39_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[13] == c_39_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[14] == c_39_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[14] == c_39_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[15] == c_39_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[15] == c_39_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[16] == c_39_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[16] == c_39_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[17] == c_39_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[17] == c_39_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[18] == c_39_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[18] == c_39_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[19] == c_39_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[19] == c_39_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[20] == c_39_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[20] == c_39_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[21] == c_39_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[21] == c_39_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[22] == c_39_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[22] == c_39_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[23] == c_39_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[23] == c_39_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[24] == c_39_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[24] == c_39_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[25] == c_39_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[25] == c_39_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[26] == c_39_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[26] == c_39_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[27] == c_39_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[27] == c_39_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[28] == c_39_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[28] == c_39_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[29] == c_39_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[29] == c_39_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[30] == c_39_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[30] == c_39_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[31] == c_39_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[31] == c_39_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_39[32] == c_39_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_39[32] == c_39_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[0] == c_40_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[0] == c_40_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[1] == c_40_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[1] == c_40_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[2] == c_40_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[2] == c_40_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[3] == c_40_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[3] == c_40_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[4] == c_40_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[4] == c_40_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[5] == c_40_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[5] == c_40_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[6] == c_40_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[6] == c_40_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[7] == c_40_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[7] == c_40_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[8] == c_40_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[8] == c_40_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[9] == c_40_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[9] == c_40_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[10] == c_40_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[10] == c_40_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[11] == c_40_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[11] == c_40_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[12] == c_40_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[12] == c_40_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[13] == c_40_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[13] == c_40_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[14] == c_40_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[14] == c_40_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[15] == c_40_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[15] == c_40_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[16] == c_40_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[16] == c_40_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[17] == c_40_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[17] == c_40_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[18] == c_40_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[18] == c_40_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[19] == c_40_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[19] == c_40_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[20] == c_40_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[20] == c_40_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[21] == c_40_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[21] == c_40_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[22] == c_40_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[22] == c_40_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[23] == c_40_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[23] == c_40_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[24] == c_40_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[24] == c_40_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[25] == c_40_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[25] == c_40_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[26] == c_40_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[26] == c_40_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[27] == c_40_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[27] == c_40_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[28] == c_40_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[28] == c_40_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[29] == c_40_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[29] == c_40_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[30] == c_40_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[30] == c_40_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[31] == c_40_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[31] == c_40_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_40[32] == c_40_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_40[32] == c_40_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[0] == c_41_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[0] == c_41_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[1] == c_41_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[1] == c_41_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[2] == c_41_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[2] == c_41_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[3] == c_41_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[3] == c_41_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[4] == c_41_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[4] == c_41_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[5] == c_41_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[5] == c_41_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[6] == c_41_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[6] == c_41_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[7] == c_41_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[7] == c_41_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[8] == c_41_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[8] == c_41_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[9] == c_41_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[9] == c_41_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[10] == c_41_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[10] == c_41_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[11] == c_41_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[11] == c_41_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[12] == c_41_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[12] == c_41_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[13] == c_41_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[13] == c_41_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[14] == c_41_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[14] == c_41_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[15] == c_41_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[15] == c_41_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[16] == c_41_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[16] == c_41_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[17] == c_41_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[17] == c_41_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[18] == c_41_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[18] == c_41_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[19] == c_41_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[19] == c_41_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[20] == c_41_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[20] == c_41_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[21] == c_41_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[21] == c_41_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[22] == c_41_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[22] == c_41_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[23] == c_41_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[23] == c_41_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[24] == c_41_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[24] == c_41_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[25] == c_41_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[25] == c_41_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[26] == c_41_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[26] == c_41_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[27] == c_41_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[27] == c_41_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[28] == c_41_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[28] == c_41_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[29] == c_41_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[29] == c_41_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[30] == c_41_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[30] == c_41_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[31] == c_41_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[31] == c_41_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_41[32] == c_41_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_41[32] == c_41_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[0] == c_42_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[0] == c_42_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[1] == c_42_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[1] == c_42_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[2] == c_42_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[2] == c_42_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[3] == c_42_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[3] == c_42_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[4] == c_42_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[4] == c_42_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[5] == c_42_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[5] == c_42_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[6] == c_42_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[6] == c_42_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[7] == c_42_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[7] == c_42_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[8] == c_42_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[8] == c_42_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[9] == c_42_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[9] == c_42_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[10] == c_42_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[10] == c_42_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[11] == c_42_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[11] == c_42_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[12] == c_42_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[12] == c_42_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[13] == c_42_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[13] == c_42_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[14] == c_42_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[14] == c_42_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[15] == c_42_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[15] == c_42_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[16] == c_42_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[16] == c_42_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[17] == c_42_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[17] == c_42_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[18] == c_42_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[18] == c_42_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[19] == c_42_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[19] == c_42_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[20] == c_42_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[20] == c_42_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[21] == c_42_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[21] == c_42_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[22] == c_42_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[22] == c_42_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[23] == c_42_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[23] == c_42_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[24] == c_42_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[24] == c_42_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[25] == c_42_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[25] == c_42_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[26] == c_42_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[26] == c_42_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[27] == c_42_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[27] == c_42_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[28] == c_42_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[28] == c_42_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[29] == c_42_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[29] == c_42_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[30] == c_42_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[30] == c_42_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[31] == c_42_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[31] == c_42_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_42[32] == c_42_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_42[32] == c_42_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[0] == c_43_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[0] == c_43_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[1] == c_43_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[1] == c_43_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[2] == c_43_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[2] == c_43_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[3] == c_43_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[3] == c_43_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[4] == c_43_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[4] == c_43_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[5] == c_43_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[5] == c_43_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[6] == c_43_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[6] == c_43_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[7] == c_43_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[7] == c_43_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[8] == c_43_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[8] == c_43_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[9] == c_43_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[9] == c_43_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[10] == c_43_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[10] == c_43_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[11] == c_43_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[11] == c_43_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[12] == c_43_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[12] == c_43_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[13] == c_43_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[13] == c_43_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[14] == c_43_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[14] == c_43_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[15] == c_43_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[15] == c_43_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[16] == c_43_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[16] == c_43_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[17] == c_43_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[17] == c_43_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[18] == c_43_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[18] == c_43_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[19] == c_43_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[19] == c_43_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[20] == c_43_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[20] == c_43_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[21] == c_43_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[21] == c_43_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[22] == c_43_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[22] == c_43_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[23] == c_43_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[23] == c_43_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[24] == c_43_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[24] == c_43_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[25] == c_43_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[25] == c_43_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[26] == c_43_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[26] == c_43_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[27] == c_43_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[27] == c_43_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[28] == c_43_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[28] == c_43_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[29] == c_43_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[29] == c_43_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[30] == c_43_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[30] == c_43_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[31] == c_43_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[31] == c_43_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_43[32] == c_43_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_43[32] == c_43_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[0] == c_44_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[0] == c_44_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[1] == c_44_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[1] == c_44_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[2] == c_44_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[2] == c_44_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[3] == c_44_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[3] == c_44_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[4] == c_44_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[4] == c_44_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[5] == c_44_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[5] == c_44_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[6] == c_44_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[6] == c_44_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[7] == c_44_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[7] == c_44_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[8] == c_44_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[8] == c_44_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[9] == c_44_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[9] == c_44_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[10] == c_44_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[10] == c_44_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[11] == c_44_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[11] == c_44_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[12] == c_44_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[12] == c_44_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[13] == c_44_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[13] == c_44_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[14] == c_44_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[14] == c_44_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[15] == c_44_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[15] == c_44_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[16] == c_44_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[16] == c_44_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[17] == c_44_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[17] == c_44_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[18] == c_44_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[18] == c_44_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[19] == c_44_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[19] == c_44_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[20] == c_44_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[20] == c_44_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[21] == c_44_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[21] == c_44_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[22] == c_44_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[22] == c_44_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[23] == c_44_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[23] == c_44_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[24] == c_44_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[24] == c_44_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[25] == c_44_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[25] == c_44_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[26] == c_44_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[26] == c_44_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[27] == c_44_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[27] == c_44_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[28] == c_44_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[28] == c_44_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[29] == c_44_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[29] == c_44_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[30] == c_44_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[30] == c_44_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[31] == c_44_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[31] == c_44_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_44[32] == c_44_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_44[32] == c_44_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[0] == c_45_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[0] == c_45_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[1] == c_45_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[1] == c_45_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[2] == c_45_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[2] == c_45_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[3] == c_45_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[3] == c_45_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[4] == c_45_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[4] == c_45_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[5] == c_45_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[5] == c_45_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[6] == c_45_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[6] == c_45_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[7] == c_45_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[7] == c_45_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[8] == c_45_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[8] == c_45_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[9] == c_45_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[9] == c_45_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[10] == c_45_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[10] == c_45_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[11] == c_45_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[11] == c_45_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[12] == c_45_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[12] == c_45_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[13] == c_45_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[13] == c_45_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[14] == c_45_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[14] == c_45_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[15] == c_45_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[15] == c_45_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[16] == c_45_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[16] == c_45_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[17] == c_45_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[17] == c_45_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[18] == c_45_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[18] == c_45_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[19] == c_45_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[19] == c_45_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[20] == c_45_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[20] == c_45_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[21] == c_45_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[21] == c_45_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[22] == c_45_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[22] == c_45_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[23] == c_45_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[23] == c_45_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[24] == c_45_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[24] == c_45_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[25] == c_45_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[25] == c_45_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[26] == c_45_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[26] == c_45_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[27] == c_45_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[27] == c_45_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[28] == c_45_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[28] == c_45_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[29] == c_45_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[29] == c_45_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[30] == c_45_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[30] == c_45_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[31] == c_45_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[31] == c_45_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_45[32] == c_45_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_45[32] == c_45_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[0] == c_46_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[0] == c_46_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[1] == c_46_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[1] == c_46_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[2] == c_46_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[2] == c_46_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[3] == c_46_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[3] == c_46_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[4] == c_46_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[4] == c_46_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[5] == c_46_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[5] == c_46_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[6] == c_46_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[6] == c_46_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[7] == c_46_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[7] == c_46_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[8] == c_46_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[8] == c_46_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[9] == c_46_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[9] == c_46_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[10] == c_46_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[10] == c_46_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[11] == c_46_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[11] == c_46_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[12] == c_46_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[12] == c_46_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[13] == c_46_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[13] == c_46_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[14] == c_46_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[14] == c_46_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[15] == c_46_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[15] == c_46_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[16] == c_46_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[16] == c_46_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[17] == c_46_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[17] == c_46_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[18] == c_46_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[18] == c_46_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[19] == c_46_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[19] == c_46_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[20] == c_46_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[20] == c_46_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[21] == c_46_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[21] == c_46_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[22] == c_46_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[22] == c_46_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[23] == c_46_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[23] == c_46_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[24] == c_46_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[24] == c_46_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[25] == c_46_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[25] == c_46_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[26] == c_46_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[26] == c_46_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[27] == c_46_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[27] == c_46_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[28] == c_46_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[28] == c_46_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[29] == c_46_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[29] == c_46_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[30] == c_46_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[30] == c_46_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[31] == c_46_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[31] == c_46_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_46[32] == c_46_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_46[32] == c_46_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[0] == c_47_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[0] == c_47_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[1] == c_47_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[1] == c_47_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[2] == c_47_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[2] == c_47_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[3] == c_47_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[3] == c_47_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[4] == c_47_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[4] == c_47_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[5] == c_47_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[5] == c_47_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[6] == c_47_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[6] == c_47_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[7] == c_47_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[7] == c_47_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[8] == c_47_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[8] == c_47_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[9] == c_47_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[9] == c_47_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[10] == c_47_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[10] == c_47_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[11] == c_47_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[11] == c_47_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[12] == c_47_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[12] == c_47_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[13] == c_47_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[13] == c_47_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[14] == c_47_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[14] == c_47_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[15] == c_47_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[15] == c_47_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[16] == c_47_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[16] == c_47_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[17] == c_47_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[17] == c_47_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[18] == c_47_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[18] == c_47_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[19] == c_47_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[19] == c_47_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[20] == c_47_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[20] == c_47_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[21] == c_47_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[21] == c_47_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[22] == c_47_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[22] == c_47_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[23] == c_47_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[23] == c_47_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[24] == c_47_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[24] == c_47_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[25] == c_47_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[25] == c_47_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[26] == c_47_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[26] == c_47_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[27] == c_47_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[27] == c_47_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[28] == c_47_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[28] == c_47_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[29] == c_47_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[29] == c_47_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[30] == c_47_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[30] == c_47_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[31] == c_47_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[31] == c_47_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_47[32] == c_47_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_47[32] == c_47_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[0] == c_48_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[0] == c_48_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[1] == c_48_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[1] == c_48_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[2] == c_48_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[2] == c_48_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[3] == c_48_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[3] == c_48_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[4] == c_48_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[4] == c_48_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[5] == c_48_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[5] == c_48_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[6] == c_48_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[6] == c_48_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[7] == c_48_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[7] == c_48_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[8] == c_48_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[8] == c_48_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[9] == c_48_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[9] == c_48_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[10] == c_48_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[10] == c_48_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[11] == c_48_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[11] == c_48_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[12] == c_48_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[12] == c_48_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[13] == c_48_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[13] == c_48_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[14] == c_48_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[14] == c_48_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[15] == c_48_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[15] == c_48_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[16] == c_48_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[16] == c_48_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[17] == c_48_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[17] == c_48_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[18] == c_48_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[18] == c_48_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[19] == c_48_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[19] == c_48_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[20] == c_48_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[20] == c_48_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[21] == c_48_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[21] == c_48_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[22] == c_48_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[22] == c_48_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[23] == c_48_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[23] == c_48_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[24] == c_48_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[24] == c_48_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[25] == c_48_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[25] == c_48_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[26] == c_48_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[26] == c_48_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[27] == c_48_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[27] == c_48_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[28] == c_48_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[28] == c_48_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[29] == c_48_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[29] == c_48_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[30] == c_48_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[30] == c_48_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[31] == c_48_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[31] == c_48_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_48[32] == c_48_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_48[32] == c_48_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[0] == c_49_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[0] == c_49_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[1] == c_49_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[1] == c_49_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[2] == c_49_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[2] == c_49_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[3] == c_49_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[3] == c_49_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[4] == c_49_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[4] == c_49_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[5] == c_49_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[5] == c_49_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[6] == c_49_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[6] == c_49_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[7] == c_49_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[7] == c_49_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[8] == c_49_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[8] == c_49_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[9] == c_49_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[9] == c_49_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[10] == c_49_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[10] == c_49_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[11] == c_49_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[11] == c_49_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[12] == c_49_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[12] == c_49_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[13] == c_49_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[13] == c_49_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[14] == c_49_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[14] == c_49_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[15] == c_49_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[15] == c_49_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[16] == c_49_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[16] == c_49_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[17] == c_49_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[17] == c_49_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[18] == c_49_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[18] == c_49_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[19] == c_49_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[19] == c_49_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[20] == c_49_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[20] == c_49_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[21] == c_49_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[21] == c_49_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[22] == c_49_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[22] == c_49_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[23] == c_49_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[23] == c_49_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[24] == c_49_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[24] == c_49_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[25] == c_49_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[25] == c_49_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[26] == c_49_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[26] == c_49_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[27] == c_49_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[27] == c_49_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[28] == c_49_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[28] == c_49_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[29] == c_49_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[29] == c_49_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[30] == c_49_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[30] == c_49_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[31] == c_49_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[31] == c_49_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_49[32] == c_49_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_49[32] == c_49_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[0] == c_50_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[0] == c_50_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[1] == c_50_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[1] == c_50_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[2] == c_50_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[2] == c_50_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[3] == c_50_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[3] == c_50_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[4] == c_50_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[4] == c_50_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[5] == c_50_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[5] == c_50_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[6] == c_50_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[6] == c_50_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[7] == c_50_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[7] == c_50_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[8] == c_50_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[8] == c_50_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[9] == c_50_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[9] == c_50_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[10] == c_50_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[10] == c_50_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[11] == c_50_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[11] == c_50_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[12] == c_50_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[12] == c_50_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[13] == c_50_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[13] == c_50_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[14] == c_50_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[14] == c_50_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[15] == c_50_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[15] == c_50_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[16] == c_50_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[16] == c_50_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[17] == c_50_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[17] == c_50_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[18] == c_50_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[18] == c_50_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[19] == c_50_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[19] == c_50_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[20] == c_50_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[20] == c_50_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[21] == c_50_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[21] == c_50_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[22] == c_50_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[22] == c_50_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[23] == c_50_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[23] == c_50_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[24] == c_50_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[24] == c_50_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[25] == c_50_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[25] == c_50_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[26] == c_50_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[26] == c_50_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[27] == c_50_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[27] == c_50_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[28] == c_50_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[28] == c_50_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[29] == c_50_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[29] == c_50_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[30] == c_50_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[30] == c_50_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[31] == c_50_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[31] == c_50_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_50[32] == c_50_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_50[32] == c_50_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[0] == c_51_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[0] == c_51_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[1] == c_51_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[1] == c_51_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[2] == c_51_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[2] == c_51_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[3] == c_51_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[3] == c_51_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[4] == c_51_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[4] == c_51_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[5] == c_51_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[5] == c_51_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[6] == c_51_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[6] == c_51_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[7] == c_51_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[7] == c_51_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[8] == c_51_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[8] == c_51_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[9] == c_51_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[9] == c_51_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[10] == c_51_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[10] == c_51_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[11] == c_51_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[11] == c_51_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[12] == c_51_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[12] == c_51_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[13] == c_51_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[13] == c_51_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[14] == c_51_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[14] == c_51_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[15] == c_51_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[15] == c_51_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[16] == c_51_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[16] == c_51_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[17] == c_51_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[17] == c_51_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[18] == c_51_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[18] == c_51_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[19] == c_51_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[19] == c_51_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[20] == c_51_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[20] == c_51_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[21] == c_51_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[21] == c_51_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[22] == c_51_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[22] == c_51_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[23] == c_51_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[23] == c_51_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[24] == c_51_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[24] == c_51_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[25] == c_51_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[25] == c_51_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[26] == c_51_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[26] == c_51_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[27] == c_51_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[27] == c_51_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[28] == c_51_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[28] == c_51_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[29] == c_51_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[29] == c_51_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[30] == c_51_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[30] == c_51_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[31] == c_51_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[31] == c_51_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_51[32] == c_51_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_51[32] == c_51_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[0] == c_52_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[0] == c_52_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[1] == c_52_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[1] == c_52_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[2] == c_52_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[2] == c_52_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[3] == c_52_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[3] == c_52_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[4] == c_52_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[4] == c_52_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[5] == c_52_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[5] == c_52_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[6] == c_52_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[6] == c_52_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[7] == c_52_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[7] == c_52_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[8] == c_52_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[8] == c_52_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[9] == c_52_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[9] == c_52_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[10] == c_52_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[10] == c_52_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[11] == c_52_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[11] == c_52_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[12] == c_52_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[12] == c_52_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[13] == c_52_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[13] == c_52_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[14] == c_52_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[14] == c_52_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[15] == c_52_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[15] == c_52_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[16] == c_52_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[16] == c_52_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[17] == c_52_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[17] == c_52_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[18] == c_52_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[18] == c_52_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[19] == c_52_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[19] == c_52_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[20] == c_52_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[20] == c_52_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[21] == c_52_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[21] == c_52_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[22] == c_52_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[22] == c_52_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[23] == c_52_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[23] == c_52_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[24] == c_52_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[24] == c_52_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[25] == c_52_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[25] == c_52_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[26] == c_52_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[26] == c_52_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[27] == c_52_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[27] == c_52_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[28] == c_52_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[28] == c_52_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[29] == c_52_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[29] == c_52_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[30] == c_52_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[30] == c_52_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[31] == c_52_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[31] == c_52_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_52[32] == c_52_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_52[32] == c_52_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[0] == c_53_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[0] == c_53_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[1] == c_53_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[1] == c_53_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[2] == c_53_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[2] == c_53_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[3] == c_53_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[3] == c_53_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[4] == c_53_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[4] == c_53_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[5] == c_53_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[5] == c_53_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[6] == c_53_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[6] == c_53_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[7] == c_53_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[7] == c_53_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[8] == c_53_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[8] == c_53_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[9] == c_53_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[9] == c_53_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[10] == c_53_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[10] == c_53_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[11] == c_53_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[11] == c_53_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[12] == c_53_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[12] == c_53_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[13] == c_53_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[13] == c_53_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[14] == c_53_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[14] == c_53_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[15] == c_53_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[15] == c_53_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[16] == c_53_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[16] == c_53_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[17] == c_53_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[17] == c_53_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[18] == c_53_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[18] == c_53_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[19] == c_53_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[19] == c_53_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[20] == c_53_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[20] == c_53_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[21] == c_53_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[21] == c_53_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[22] == c_53_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[22] == c_53_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[23] == c_53_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[23] == c_53_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[24] == c_53_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[24] == c_53_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[25] == c_53_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[25] == c_53_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[26] == c_53_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[26] == c_53_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[27] == c_53_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[27] == c_53_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[28] == c_53_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[28] == c_53_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[29] == c_53_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[29] == c_53_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[30] == c_53_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[30] == c_53_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[31] == c_53_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[31] == c_53_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_53[32] == c_53_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_53[32] == c_53_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[0] == c_54_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[0] == c_54_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[1] == c_54_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[1] == c_54_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[2] == c_54_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[2] == c_54_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[3] == c_54_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[3] == c_54_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[4] == c_54_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[4] == c_54_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[5] == c_54_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[5] == c_54_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[6] == c_54_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[6] == c_54_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[7] == c_54_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[7] == c_54_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[8] == c_54_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[8] == c_54_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[9] == c_54_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[9] == c_54_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[10] == c_54_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[10] == c_54_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[11] == c_54_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[11] == c_54_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[12] == c_54_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[12] == c_54_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[13] == c_54_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[13] == c_54_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[14] == c_54_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[14] == c_54_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[15] == c_54_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[15] == c_54_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[16] == c_54_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[16] == c_54_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[17] == c_54_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[17] == c_54_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[18] == c_54_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[18] == c_54_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[19] == c_54_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[19] == c_54_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[20] == c_54_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[20] == c_54_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[21] == c_54_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[21] == c_54_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[22] == c_54_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[22] == c_54_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[23] == c_54_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[23] == c_54_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[24] == c_54_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[24] == c_54_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[25] == c_54_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[25] == c_54_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[26] == c_54_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[26] == c_54_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[27] == c_54_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[27] == c_54_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[28] == c_54_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[28] == c_54_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[29] == c_54_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[29] == c_54_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[30] == c_54_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[30] == c_54_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[31] == c_54_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[31] == c_54_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_54[32] == c_54_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_54[32] == c_54_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[0] == c_55_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[0] == c_55_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[1] == c_55_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[1] == c_55_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[2] == c_55_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[2] == c_55_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[3] == c_55_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[3] == c_55_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[4] == c_55_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[4] == c_55_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[5] == c_55_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[5] == c_55_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[6] == c_55_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[6] == c_55_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[7] == c_55_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[7] == c_55_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[8] == c_55_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[8] == c_55_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[9] == c_55_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[9] == c_55_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[10] == c_55_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[10] == c_55_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[11] == c_55_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[11] == c_55_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[12] == c_55_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[12] == c_55_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[13] == c_55_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[13] == c_55_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[14] == c_55_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[14] == c_55_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[15] == c_55_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[15] == c_55_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[16] == c_55_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[16] == c_55_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[17] == c_55_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[17] == c_55_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[18] == c_55_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[18] == c_55_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[19] == c_55_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[19] == c_55_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[20] == c_55_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[20] == c_55_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[21] == c_55_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[21] == c_55_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[22] == c_55_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[22] == c_55_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[23] == c_55_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[23] == c_55_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[24] == c_55_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[24] == c_55_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[25] == c_55_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[25] == c_55_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[26] == c_55_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[26] == c_55_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[27] == c_55_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[27] == c_55_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[28] == c_55_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[28] == c_55_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[29] == c_55_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[29] == c_55_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[30] == c_55_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[30] == c_55_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[31] == c_55_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[31] == c_55_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_55[32] == c_55_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_55[32] == c_55_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[0] == c_56_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[0] == c_56_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[1] == c_56_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[1] == c_56_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[2] == c_56_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[2] == c_56_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[3] == c_56_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[3] == c_56_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[4] == c_56_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[4] == c_56_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[5] == c_56_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[5] == c_56_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[6] == c_56_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[6] == c_56_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[7] == c_56_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[7] == c_56_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[8] == c_56_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[8] == c_56_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[9] == c_56_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[9] == c_56_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[10] == c_56_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[10] == c_56_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[11] == c_56_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[11] == c_56_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[12] == c_56_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[12] == c_56_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[13] == c_56_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[13] == c_56_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[14] == c_56_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[14] == c_56_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[15] == c_56_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[15] == c_56_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[16] == c_56_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[16] == c_56_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[17] == c_56_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[17] == c_56_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[18] == c_56_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[18] == c_56_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[19] == c_56_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[19] == c_56_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[20] == c_56_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[20] == c_56_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[21] == c_56_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[21] == c_56_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[22] == c_56_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[22] == c_56_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[23] == c_56_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[23] == c_56_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[24] == c_56_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[24] == c_56_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[25] == c_56_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[25] == c_56_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[26] == c_56_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[26] == c_56_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[27] == c_56_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[27] == c_56_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[28] == c_56_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[28] == c_56_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[29] == c_56_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[29] == c_56_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[30] == c_56_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[30] == c_56_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[31] == c_56_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[31] == c_56_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_56[32] == c_56_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_56[32] == c_56_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[0] == c_57_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[0] == c_57_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[1] == c_57_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[1] == c_57_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[2] == c_57_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[2] == c_57_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[3] == c_57_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[3] == c_57_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[4] == c_57_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[4] == c_57_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[5] == c_57_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[5] == c_57_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[6] == c_57_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[6] == c_57_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[7] == c_57_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[7] == c_57_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[8] == c_57_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[8] == c_57_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[9] == c_57_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[9] == c_57_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[10] == c_57_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[10] == c_57_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[11] == c_57_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[11] == c_57_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[12] == c_57_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[12] == c_57_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[13] == c_57_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[13] == c_57_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[14] == c_57_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[14] == c_57_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[15] == c_57_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[15] == c_57_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[16] == c_57_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[16] == c_57_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[17] == c_57_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[17] == c_57_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[18] == c_57_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[18] == c_57_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[19] == c_57_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[19] == c_57_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[20] == c_57_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[20] == c_57_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[21] == c_57_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[21] == c_57_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[22] == c_57_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[22] == c_57_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[23] == c_57_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[23] == c_57_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[24] == c_57_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[24] == c_57_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[25] == c_57_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[25] == c_57_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[26] == c_57_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[26] == c_57_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[27] == c_57_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[27] == c_57_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[28] == c_57_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[28] == c_57_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[29] == c_57_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[29] == c_57_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[30] == c_57_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[30] == c_57_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[31] == c_57_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[31] == c_57_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_57[32] == c_57_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_57[32] == c_57_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[0] == c_58_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[0] == c_58_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[1] == c_58_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[1] == c_58_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[2] == c_58_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[2] == c_58_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[3] == c_58_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[3] == c_58_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[4] == c_58_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[4] == c_58_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[5] == c_58_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[5] == c_58_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[6] == c_58_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[6] == c_58_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[7] == c_58_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[7] == c_58_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[8] == c_58_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[8] == c_58_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[9] == c_58_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[9] == c_58_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[10] == c_58_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[10] == c_58_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[11] == c_58_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[11] == c_58_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[12] == c_58_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[12] == c_58_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[13] == c_58_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[13] == c_58_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[14] == c_58_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[14] == c_58_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[15] == c_58_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[15] == c_58_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[16] == c_58_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[16] == c_58_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[17] == c_58_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[17] == c_58_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[18] == c_58_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[18] == c_58_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[19] == c_58_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[19] == c_58_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[20] == c_58_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[20] == c_58_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[21] == c_58_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[21] == c_58_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[22] == c_58_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[22] == c_58_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[23] == c_58_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[23] == c_58_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[24] == c_58_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[24] == c_58_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[25] == c_58_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[25] == c_58_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[26] == c_58_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[26] == c_58_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[27] == c_58_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[27] == c_58_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[28] == c_58_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[28] == c_58_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[29] == c_58_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[29] == c_58_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[30] == c_58_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[30] == c_58_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[31] == c_58_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[31] == c_58_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_58[32] == c_58_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_58[32] == c_58_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[0] == c_59_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[0] == c_59_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[1] == c_59_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[1] == c_59_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[2] == c_59_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[2] == c_59_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[3] == c_59_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[3] == c_59_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[4] == c_59_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[4] == c_59_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[5] == c_59_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[5] == c_59_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[6] == c_59_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[6] == c_59_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[7] == c_59_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[7] == c_59_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[8] == c_59_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[8] == c_59_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[9] == c_59_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[9] == c_59_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[10] == c_59_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[10] == c_59_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[11] == c_59_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[11] == c_59_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[12] == c_59_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[12] == c_59_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[13] == c_59_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[13] == c_59_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[14] == c_59_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[14] == c_59_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[15] == c_59_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[15] == c_59_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[16] == c_59_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[16] == c_59_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[17] == c_59_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[17] == c_59_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[18] == c_59_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[18] == c_59_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[19] == c_59_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[19] == c_59_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[20] == c_59_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[20] == c_59_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[21] == c_59_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[21] == c_59_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[22] == c_59_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[22] == c_59_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[23] == c_59_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[23] == c_59_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[24] == c_59_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[24] == c_59_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[25] == c_59_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[25] == c_59_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[26] == c_59_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[26] == c_59_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[27] == c_59_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[27] == c_59_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[28] == c_59_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[28] == c_59_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[29] == c_59_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[29] == c_59_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[30] == c_59_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[30] == c_59_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[31] == c_59_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[31] == c_59_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_59[32] == c_59_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_59[32] == c_59_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[0] == c_60_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[0] == c_60_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[1] == c_60_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[1] == c_60_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[2] == c_60_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[2] == c_60_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[3] == c_60_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[3] == c_60_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[4] == c_60_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[4] == c_60_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[5] == c_60_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[5] == c_60_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[6] == c_60_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[6] == c_60_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[7] == c_60_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[7] == c_60_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[8] == c_60_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[8] == c_60_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[9] == c_60_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[9] == c_60_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[10] == c_60_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[10] == c_60_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[11] == c_60_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[11] == c_60_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[12] == c_60_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[12] == c_60_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[13] == c_60_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[13] == c_60_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[14] == c_60_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[14] == c_60_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[15] == c_60_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[15] == c_60_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[16] == c_60_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[16] == c_60_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[17] == c_60_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[17] == c_60_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[18] == c_60_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[18] == c_60_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[19] == c_60_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[19] == c_60_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[20] == c_60_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[20] == c_60_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[21] == c_60_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[21] == c_60_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[22] == c_60_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[22] == c_60_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[23] == c_60_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[23] == c_60_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[24] == c_60_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[24] == c_60_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[25] == c_60_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[25] == c_60_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[26] == c_60_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[26] == c_60_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[27] == c_60_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[27] == c_60_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[28] == c_60_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[28] == c_60_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[29] == c_60_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[29] == c_60_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[30] == c_60_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[30] == c_60_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[31] == c_60_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[31] == c_60_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_60[32] == c_60_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_60[32] == c_60_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[0] == c_61_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[0] == c_61_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[1] == c_61_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[1] == c_61_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[2] == c_61_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[2] == c_61_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[3] == c_61_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[3] == c_61_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[4] == c_61_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[4] == c_61_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[5] == c_61_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[5] == c_61_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[6] == c_61_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[6] == c_61_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[7] == c_61_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[7] == c_61_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[8] == c_61_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[8] == c_61_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[9] == c_61_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[9] == c_61_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[10] == c_61_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[10] == c_61_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[11] == c_61_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[11] == c_61_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[12] == c_61_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[12] == c_61_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[13] == c_61_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[13] == c_61_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[14] == c_61_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[14] == c_61_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[15] == c_61_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[15] == c_61_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[16] == c_61_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[16] == c_61_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[17] == c_61_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[17] == c_61_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[18] == c_61_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[18] == c_61_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[19] == c_61_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[19] == c_61_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[20] == c_61_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[20] == c_61_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[21] == c_61_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[21] == c_61_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[22] == c_61_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[22] == c_61_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[23] == c_61_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[23] == c_61_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[24] == c_61_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[24] == c_61_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[25] == c_61_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[25] == c_61_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[26] == c_61_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[26] == c_61_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[27] == c_61_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[27] == c_61_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[28] == c_61_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[28] == c_61_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[29] == c_61_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[29] == c_61_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[30] == c_61_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[30] == c_61_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[31] == c_61_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[31] == c_61_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_61[32] == c_61_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_61[32] == c_61_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[0] == c_62_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[0] == c_62_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[1] == c_62_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[1] == c_62_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[2] == c_62_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[2] == c_62_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[3] == c_62_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[3] == c_62_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[4] == c_62_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[4] == c_62_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[5] == c_62_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[5] == c_62_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[6] == c_62_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[6] == c_62_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[7] == c_62_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[7] == c_62_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[8] == c_62_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[8] == c_62_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[9] == c_62_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[9] == c_62_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[10] == c_62_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[10] == c_62_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[11] == c_62_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[11] == c_62_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[12] == c_62_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[12] == c_62_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[13] == c_62_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[13] == c_62_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[14] == c_62_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[14] == c_62_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[15] == c_62_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[15] == c_62_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[16] == c_62_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[16] == c_62_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[17] == c_62_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[17] == c_62_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[18] == c_62_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[18] == c_62_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[19] == c_62_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[19] == c_62_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[20] == c_62_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[20] == c_62_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[21] == c_62_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[21] == c_62_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[22] == c_62_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[22] == c_62_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[23] == c_62_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[23] == c_62_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[24] == c_62_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[24] == c_62_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[25] == c_62_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[25] == c_62_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[26] == c_62_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[26] == c_62_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[27] == c_62_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[27] == c_62_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[28] == c_62_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[28] == c_62_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[29] == c_62_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[29] == c_62_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[30] == c_62_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[30] == c_62_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[31] == c_62_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[31] == c_62_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_62[32] == c_62_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_62[32] == c_62_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[0] == c_63_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[0] == c_63_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[1] == c_63_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[1] == c_63_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[2] == c_63_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[2] == c_63_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[3] == c_63_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[3] == c_63_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[4] == c_63_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[4] == c_63_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[5] == c_63_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[5] == c_63_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[6] == c_63_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[6] == c_63_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[7] == c_63_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[7] == c_63_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[8] == c_63_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[8] == c_63_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[9] == c_63_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[9] == c_63_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[10] == c_63_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[10] == c_63_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[11] == c_63_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[11] == c_63_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[12] == c_63_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[12] == c_63_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[13] == c_63_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[13] == c_63_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[14] == c_63_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[14] == c_63_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[15] == c_63_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[15] == c_63_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[16] == c_63_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[16] == c_63_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[17] == c_63_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[17] == c_63_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[18] == c_63_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[18] == c_63_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[19] == c_63_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[19] == c_63_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[20] == c_63_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[20] == c_63_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[21] == c_63_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[21] == c_63_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[22] == c_63_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[22] == c_63_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[23] == c_63_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[23] == c_63_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[24] == c_63_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[24] == c_63_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[25] == c_63_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[25] == c_63_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[26] == c_63_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[26] == c_63_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[27] == c_63_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[27] == c_63_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[28] == c_63_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[28] == c_63_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[29] == c_63_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[29] == c_63_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[30] == c_63_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[30] == c_63_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[31] == c_63_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[31] == c_63_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_63[32] == c_63_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_63[32] == c_63_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[0] == c_64_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[0] == c_64_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[1] == c_64_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[1] == c_64_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[2] == c_64_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[2] == c_64_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[3] == c_64_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[3] == c_64_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[4] == c_64_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[4] == c_64_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[5] == c_64_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[5] == c_64_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[6] == c_64_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[6] == c_64_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[7] == c_64_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[7] == c_64_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[8] == c_64_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[8] == c_64_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[9] == c_64_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[9] == c_64_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[10] == c_64_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[10] == c_64_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[11] == c_64_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[11] == c_64_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[12] == c_64_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[12] == c_64_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[13] == c_64_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[13] == c_64_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[14] == c_64_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[14] == c_64_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[15] == c_64_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[15] == c_64_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[16] == c_64_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[16] == c_64_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[17] == c_64_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[17] == c_64_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[18] == c_64_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[18] == c_64_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[19] == c_64_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[19] == c_64_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[20] == c_64_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[20] == c_64_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[21] == c_64_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[21] == c_64_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[22] == c_64_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[22] == c_64_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[23] == c_64_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[23] == c_64_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[24] == c_64_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[24] == c_64_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[25] == c_64_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[25] == c_64_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[26] == c_64_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[26] == c_64_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[27] == c_64_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[27] == c_64_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[28] == c_64_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[28] == c_64_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[29] == c_64_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[29] == c_64_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[30] == c_64_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[30] == c_64_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[31] == c_64_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[31] == c_64_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_64[32] == c_64_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_64[32] == c_64_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[0] == c_65_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[0] == c_65_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[1] == c_65_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[1] == c_65_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[2] == c_65_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[2] == c_65_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[3] == c_65_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[3] == c_65_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[4] == c_65_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[4] == c_65_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[5] == c_65_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[5] == c_65_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[6] == c_65_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[6] == c_65_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[7] == c_65_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[7] == c_65_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[8] == c_65_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[8] == c_65_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[9] == c_65_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[9] == c_65_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[10] == c_65_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[10] == c_65_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[11] == c_65_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[11] == c_65_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[12] == c_65_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[12] == c_65_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[13] == c_65_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[13] == c_65_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[14] == c_65_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[14] == c_65_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[15] == c_65_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[15] == c_65_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[16] == c_65_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[16] == c_65_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[17] == c_65_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[17] == c_65_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[18] == c_65_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[18] == c_65_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[19] == c_65_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[19] == c_65_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[20] == c_65_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[20] == c_65_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[21] == c_65_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[21] == c_65_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[22] == c_65_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[22] == c_65_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[23] == c_65_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[23] == c_65_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[24] == c_65_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[24] == c_65_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[25] == c_65_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[25] == c_65_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[26] == c_65_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[26] == c_65_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[27] == c_65_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[27] == c_65_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[28] == c_65_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[28] == c_65_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[29] == c_65_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[29] == c_65_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[30] == c_65_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[30] == c_65_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[31] == c_65_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[31] == c_65_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_65[32] == c_65_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_65[32] == c_65_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[0] == c_66_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[0] == c_66_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[1] == c_66_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[1] == c_66_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[2] == c_66_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[2] == c_66_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[3] == c_66_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[3] == c_66_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[4] == c_66_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[4] == c_66_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[5] == c_66_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[5] == c_66_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[6] == c_66_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[6] == c_66_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[7] == c_66_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[7] == c_66_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[8] == c_66_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[8] == c_66_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[9] == c_66_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[9] == c_66_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[10] == c_66_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[10] == c_66_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[11] == c_66_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[11] == c_66_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[12] == c_66_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[12] == c_66_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[13] == c_66_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[13] == c_66_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[14] == c_66_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[14] == c_66_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[15] == c_66_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[15] == c_66_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[16] == c_66_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[16] == c_66_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[17] == c_66_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[17] == c_66_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[18] == c_66_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[18] == c_66_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[19] == c_66_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[19] == c_66_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[20] == c_66_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[20] == c_66_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[21] == c_66_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[21] == c_66_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[22] == c_66_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[22] == c_66_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[23] == c_66_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[23] == c_66_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[24] == c_66_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[24] == c_66_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[25] == c_66_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[25] == c_66_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[26] == c_66_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[26] == c_66_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[27] == c_66_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[27] == c_66_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[28] == c_66_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[28] == c_66_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[29] == c_66_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[29] == c_66_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[30] == c_66_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[30] == c_66_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[31] == c_66_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[31] == c_66_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_66[32] == c_66_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_66[32] == c_66_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[0] == c_67_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[0] == c_67_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[1] == c_67_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[1] == c_67_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[2] == c_67_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[2] == c_67_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[3] == c_67_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[3] == c_67_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[4] == c_67_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[4] == c_67_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[5] == c_67_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[5] == c_67_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[6] == c_67_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[6] == c_67_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[7] == c_67_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[7] == c_67_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[8] == c_67_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[8] == c_67_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[9] == c_67_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[9] == c_67_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[10] == c_67_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[10] == c_67_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[11] == c_67_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[11] == c_67_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[12] == c_67_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[12] == c_67_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[13] == c_67_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[13] == c_67_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[14] == c_67_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[14] == c_67_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[15] == c_67_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[15] == c_67_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[16] == c_67_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[16] == c_67_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[17] == c_67_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[17] == c_67_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[18] == c_67_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[18] == c_67_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[19] == c_67_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[19] == c_67_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[20] == c_67_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[20] == c_67_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[21] == c_67_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[21] == c_67_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[22] == c_67_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[22] == c_67_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[23] == c_67_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[23] == c_67_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[24] == c_67_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[24] == c_67_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[25] == c_67_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[25] == c_67_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[26] == c_67_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[26] == c_67_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[27] == c_67_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[27] == c_67_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[28] == c_67_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[28] == c_67_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[29] == c_67_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[29] == c_67_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[30] == c_67_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[30] == c_67_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[31] == c_67_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[31] == c_67_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_67[32] == c_67_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_67[32] == c_67_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[0] == c_68_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[0] == c_68_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[1] == c_68_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[1] == c_68_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[2] == c_68_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[2] == c_68_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[3] == c_68_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[3] == c_68_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[4] == c_68_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[4] == c_68_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[5] == c_68_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[5] == c_68_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[6] == c_68_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[6] == c_68_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[7] == c_68_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[7] == c_68_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[8] == c_68_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[8] == c_68_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[9] == c_68_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[9] == c_68_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[10] == c_68_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[10] == c_68_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[11] == c_68_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[11] == c_68_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[12] == c_68_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[12] == c_68_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[13] == c_68_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[13] == c_68_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[14] == c_68_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[14] == c_68_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[15] == c_68_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[15] == c_68_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[16] == c_68_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[16] == c_68_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[17] == c_68_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[17] == c_68_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[18] == c_68_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[18] == c_68_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[19] == c_68_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[19] == c_68_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[20] == c_68_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[20] == c_68_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[21] == c_68_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[21] == c_68_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[22] == c_68_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[22] == c_68_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[23] == c_68_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[23] == c_68_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[24] == c_68_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[24] == c_68_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[25] == c_68_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[25] == c_68_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[26] == c_68_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[26] == c_68_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[27] == c_68_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[27] == c_68_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[28] == c_68_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[28] == c_68_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[29] == c_68_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[29] == c_68_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[30] == c_68_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[30] == c_68_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[31] == c_68_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[31] == c_68_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_68[32] == c_68_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_68[32] == c_68_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[0] == c_69_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[0] == c_69_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[1] == c_69_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[1] == c_69_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[2] == c_69_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[2] == c_69_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[3] == c_69_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[3] == c_69_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[4] == c_69_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[4] == c_69_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[5] == c_69_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[5] == c_69_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[6] == c_69_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[6] == c_69_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[7] == c_69_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[7] == c_69_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[8] == c_69_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[8] == c_69_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[9] == c_69_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[9] == c_69_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[10] == c_69_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[10] == c_69_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[11] == c_69_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[11] == c_69_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[12] == c_69_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[12] == c_69_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[13] == c_69_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[13] == c_69_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[14] == c_69_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[14] == c_69_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[15] == c_69_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[15] == c_69_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[16] == c_69_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[16] == c_69_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[17] == c_69_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[17] == c_69_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[18] == c_69_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[18] == c_69_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[19] == c_69_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[19] == c_69_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[20] == c_69_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[20] == c_69_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[21] == c_69_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[21] == c_69_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[22] == c_69_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[22] == c_69_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[23] == c_69_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[23] == c_69_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[24] == c_69_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[24] == c_69_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[25] == c_69_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[25] == c_69_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[26] == c_69_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[26] == c_69_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[27] == c_69_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[27] == c_69_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[28] == c_69_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[28] == c_69_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[29] == c_69_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[29] == c_69_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[30] == c_69_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[30] == c_69_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[31] == c_69_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[31] == c_69_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_69[32] == c_69_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_69[32] == c_69_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[0] == c_70_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[0] == c_70_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[1] == c_70_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[1] == c_70_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[2] == c_70_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[2] == c_70_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[3] == c_70_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[3] == c_70_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[4] == c_70_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[4] == c_70_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[5] == c_70_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[5] == c_70_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[6] == c_70_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[6] == c_70_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[7] == c_70_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[7] == c_70_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[8] == c_70_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[8] == c_70_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[9] == c_70_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[9] == c_70_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[10] == c_70_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[10] == c_70_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[11] == c_70_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[11] == c_70_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[12] == c_70_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[12] == c_70_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[13] == c_70_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[13] == c_70_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[14] == c_70_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[14] == c_70_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[15] == c_70_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[15] == c_70_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[16] == c_70_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[16] == c_70_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[17] == c_70_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[17] == c_70_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[18] == c_70_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[18] == c_70_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[19] == c_70_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[19] == c_70_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[20] == c_70_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[20] == c_70_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[21] == c_70_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[21] == c_70_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[22] == c_70_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[22] == c_70_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[23] == c_70_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[23] == c_70_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[24] == c_70_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[24] == c_70_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[25] == c_70_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[25] == c_70_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[26] == c_70_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[26] == c_70_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[27] == c_70_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[27] == c_70_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[28] == c_70_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[28] == c_70_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[29] == c_70_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[29] == c_70_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[30] == c_70_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[30] == c_70_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[31] == c_70_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[31] == c_70_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_70[32] == c_70_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_70[32] == c_70_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[0] == c_71_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[0] == c_71_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[1] == c_71_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[1] == c_71_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[2] == c_71_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[2] == c_71_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[3] == c_71_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[3] == c_71_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[4] == c_71_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[4] == c_71_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[5] == c_71_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[5] == c_71_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[6] == c_71_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[6] == c_71_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[7] == c_71_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[7] == c_71_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[8] == c_71_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[8] == c_71_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[9] == c_71_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[9] == c_71_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[10] == c_71_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[10] == c_71_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[11] == c_71_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[11] == c_71_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[12] == c_71_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[12] == c_71_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[13] == c_71_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[13] == c_71_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[14] == c_71_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[14] == c_71_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[15] == c_71_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[15] == c_71_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[16] == c_71_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[16] == c_71_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[17] == c_71_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[17] == c_71_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[18] == c_71_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[18] == c_71_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[19] == c_71_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[19] == c_71_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[20] == c_71_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[20] == c_71_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[21] == c_71_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[21] == c_71_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[22] == c_71_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[22] == c_71_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[23] == c_71_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[23] == c_71_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[24] == c_71_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[24] == c_71_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[25] == c_71_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[25] == c_71_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[26] == c_71_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[26] == c_71_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[27] == c_71_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[27] == c_71_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[28] == c_71_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[28] == c_71_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[29] == c_71_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[29] == c_71_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[30] == c_71_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[30] == c_71_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[31] == c_71_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[31] == c_71_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_71[32] == c_71_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_71[32] == c_71_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[0] == c_72_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[0] == c_72_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[1] == c_72_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[1] == c_72_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[2] == c_72_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[2] == c_72_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[3] == c_72_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[3] == c_72_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[4] == c_72_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[4] == c_72_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[5] == c_72_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[5] == c_72_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[6] == c_72_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[6] == c_72_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[7] == c_72_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[7] == c_72_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[8] == c_72_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[8] == c_72_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[9] == c_72_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[9] == c_72_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[10] == c_72_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[10] == c_72_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[11] == c_72_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[11] == c_72_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[12] == c_72_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[12] == c_72_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[13] == c_72_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[13] == c_72_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[14] == c_72_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[14] == c_72_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[15] == c_72_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[15] == c_72_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[16] == c_72_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[16] == c_72_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[17] == c_72_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[17] == c_72_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[18] == c_72_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[18] == c_72_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[19] == c_72_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[19] == c_72_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[20] == c_72_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[20] == c_72_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[21] == c_72_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[21] == c_72_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[22] == c_72_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[22] == c_72_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[23] == c_72_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[23] == c_72_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[24] == c_72_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[24] == c_72_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[25] == c_72_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[25] == c_72_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[26] == c_72_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[26] == c_72_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[27] == c_72_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[27] == c_72_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[28] == c_72_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[28] == c_72_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[29] == c_72_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[29] == c_72_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[30] == c_72_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[30] == c_72_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[31] == c_72_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[31] == c_72_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_72[32] == c_72_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_72[32] == c_72_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[0] == c_73_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[0] == c_73_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[1] == c_73_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[1] == c_73_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[2] == c_73_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[2] == c_73_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[3] == c_73_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[3] == c_73_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[4] == c_73_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[4] == c_73_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[5] == c_73_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[5] == c_73_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[6] == c_73_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[6] == c_73_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[7] == c_73_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[7] == c_73_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[8] == c_73_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[8] == c_73_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[9] == c_73_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[9] == c_73_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[10] == c_73_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[10] == c_73_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[11] == c_73_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[11] == c_73_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[12] == c_73_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[12] == c_73_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[13] == c_73_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[13] == c_73_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[14] == c_73_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[14] == c_73_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[15] == c_73_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[15] == c_73_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[16] == c_73_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[16] == c_73_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[17] == c_73_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[17] == c_73_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[18] == c_73_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[18] == c_73_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[19] == c_73_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[19] == c_73_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[20] == c_73_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[20] == c_73_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[21] == c_73_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[21] == c_73_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[22] == c_73_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[22] == c_73_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[23] == c_73_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[23] == c_73_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[24] == c_73_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[24] == c_73_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[25] == c_73_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[25] == c_73_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[26] == c_73_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[26] == c_73_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[27] == c_73_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[27] == c_73_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[28] == c_73_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[28] == c_73_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[29] == c_73_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[29] == c_73_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[30] == c_73_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[30] == c_73_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[31] == c_73_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[31] == c_73_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_73[32] == c_73_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_73[32] == c_73_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[0] == c_74_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[0] == c_74_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[1] == c_74_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[1] == c_74_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[2] == c_74_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[2] == c_74_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[3] == c_74_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[3] == c_74_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[4] == c_74_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[4] == c_74_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[5] == c_74_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[5] == c_74_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[6] == c_74_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[6] == c_74_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[7] == c_74_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[7] == c_74_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[8] == c_74_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[8] == c_74_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[9] == c_74_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[9] == c_74_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[10] == c_74_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[10] == c_74_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[11] == c_74_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[11] == c_74_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[12] == c_74_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[12] == c_74_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[13] == c_74_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[13] == c_74_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[14] == c_74_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[14] == c_74_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[15] == c_74_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[15] == c_74_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[16] == c_74_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[16] == c_74_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[17] == c_74_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[17] == c_74_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[18] == c_74_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[18] == c_74_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[19] == c_74_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[19] == c_74_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[20] == c_74_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[20] == c_74_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[21] == c_74_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[21] == c_74_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[22] == c_74_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[22] == c_74_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[23] == c_74_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[23] == c_74_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[24] == c_74_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[24] == c_74_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[25] == c_74_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[25] == c_74_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[26] == c_74_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[26] == c_74_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[27] == c_74_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[27] == c_74_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[28] == c_74_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[28] == c_74_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[29] == c_74_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[29] == c_74_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[30] == c_74_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[30] == c_74_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[31] == c_74_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[31] == c_74_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_74[32] == c_74_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_74[32] == c_74_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[0] == c_75_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[0] == c_75_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[1] == c_75_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[1] == c_75_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[2] == c_75_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[2] == c_75_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[3] == c_75_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[3] == c_75_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[4] == c_75_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[4] == c_75_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[5] == c_75_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[5] == c_75_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[6] == c_75_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[6] == c_75_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[7] == c_75_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[7] == c_75_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[8] == c_75_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[8] == c_75_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[9] == c_75_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[9] == c_75_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[10] == c_75_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[10] == c_75_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[11] == c_75_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[11] == c_75_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[12] == c_75_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[12] == c_75_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[13] == c_75_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[13] == c_75_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[14] == c_75_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[14] == c_75_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[15] == c_75_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[15] == c_75_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[16] == c_75_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[16] == c_75_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[17] == c_75_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[17] == c_75_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[18] == c_75_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[18] == c_75_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[19] == c_75_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[19] == c_75_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[20] == c_75_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[20] == c_75_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[21] == c_75_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[21] == c_75_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[22] == c_75_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[22] == c_75_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[23] == c_75_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[23] == c_75_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[24] == c_75_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[24] == c_75_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[25] == c_75_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[25] == c_75_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[26] == c_75_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[26] == c_75_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[27] == c_75_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[27] == c_75_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[28] == c_75_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[28] == c_75_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[29] == c_75_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[29] == c_75_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[30] == c_75_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[30] == c_75_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[31] == c_75_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[31] == c_75_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_75[32] == c_75_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_75[32] == c_75_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[0] == c_76_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[0] == c_76_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[1] == c_76_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[1] == c_76_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[2] == c_76_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[2] == c_76_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[3] == c_76_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[3] == c_76_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[4] == c_76_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[4] == c_76_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[5] == c_76_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[5] == c_76_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[6] == c_76_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[6] == c_76_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[7] == c_76_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[7] == c_76_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[8] == c_76_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[8] == c_76_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[9] == c_76_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[9] == c_76_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[10] == c_76_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[10] == c_76_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[11] == c_76_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[11] == c_76_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[12] == c_76_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[12] == c_76_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[13] == c_76_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[13] == c_76_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[14] == c_76_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[14] == c_76_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[15] == c_76_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[15] == c_76_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[16] == c_76_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[16] == c_76_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[17] == c_76_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[17] == c_76_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[18] == c_76_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[18] == c_76_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[19] == c_76_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[19] == c_76_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[20] == c_76_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[20] == c_76_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[21] == c_76_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[21] == c_76_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[22] == c_76_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[22] == c_76_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[23] == c_76_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[23] == c_76_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[24] == c_76_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[24] == c_76_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[25] == c_76_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[25] == c_76_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[26] == c_76_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[26] == c_76_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[27] == c_76_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[27] == c_76_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[28] == c_76_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[28] == c_76_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[29] == c_76_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[29] == c_76_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[30] == c_76_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[30] == c_76_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[31] == c_76_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[31] == c_76_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_76[32] == c_76_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_76[32] == c_76_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[0] == c_77_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[0] == c_77_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[1] == c_77_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[1] == c_77_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[2] == c_77_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[2] == c_77_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[3] == c_77_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[3] == c_77_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[4] == c_77_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[4] == c_77_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[5] == c_77_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[5] == c_77_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[6] == c_77_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[6] == c_77_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[7] == c_77_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[7] == c_77_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[8] == c_77_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[8] == c_77_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[9] == c_77_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[9] == c_77_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[10] == c_77_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[10] == c_77_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[11] == c_77_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[11] == c_77_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[12] == c_77_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[12] == c_77_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[13] == c_77_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[13] == c_77_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[14] == c_77_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[14] == c_77_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[15] == c_77_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[15] == c_77_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[16] == c_77_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[16] == c_77_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[17] == c_77_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[17] == c_77_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[18] == c_77_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[18] == c_77_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[19] == c_77_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[19] == c_77_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[20] == c_77_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[20] == c_77_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[21] == c_77_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[21] == c_77_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[22] == c_77_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[22] == c_77_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[23] == c_77_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[23] == c_77_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[24] == c_77_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[24] == c_77_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[25] == c_77_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[25] == c_77_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[26] == c_77_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[26] == c_77_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[27] == c_77_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[27] == c_77_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[28] == c_77_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[28] == c_77_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[29] == c_77_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[29] == c_77_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[30] == c_77_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[30] == c_77_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[31] == c_77_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[31] == c_77_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_77[32] == c_77_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_77[32] == c_77_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[0] == c_78_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[0] == c_78_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[1] == c_78_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[1] == c_78_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[2] == c_78_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[2] == c_78_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[3] == c_78_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[3] == c_78_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[4] == c_78_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[4] == c_78_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[5] == c_78_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[5] == c_78_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[6] == c_78_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[6] == c_78_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[7] == c_78_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[7] == c_78_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[8] == c_78_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[8] == c_78_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[9] == c_78_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[9] == c_78_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[10] == c_78_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[10] == c_78_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[11] == c_78_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[11] == c_78_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[12] == c_78_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[12] == c_78_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[13] == c_78_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[13] == c_78_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[14] == c_78_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[14] == c_78_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[15] == c_78_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[15] == c_78_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[16] == c_78_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[16] == c_78_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[17] == c_78_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[17] == c_78_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[18] == c_78_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[18] == c_78_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[19] == c_78_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[19] == c_78_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[20] == c_78_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[20] == c_78_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[21] == c_78_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[21] == c_78_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[22] == c_78_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[22] == c_78_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[23] == c_78_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[23] == c_78_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[24] == c_78_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[24] == c_78_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[25] == c_78_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[25] == c_78_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[26] == c_78_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[26] == c_78_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[27] == c_78_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[27] == c_78_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[28] == c_78_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[28] == c_78_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[29] == c_78_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[29] == c_78_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[30] == c_78_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[30] == c_78_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[31] == c_78_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[31] == c_78_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_78[32] == c_78_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_78[32] == c_78_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[0] == c_79_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[0] == c_79_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[1] == c_79_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[1] == c_79_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[2] == c_79_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[2] == c_79_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[3] == c_79_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[3] == c_79_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[4] == c_79_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[4] == c_79_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[5] == c_79_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[5] == c_79_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[6] == c_79_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[6] == c_79_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[7] == c_79_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[7] == c_79_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[8] == c_79_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[8] == c_79_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[9] == c_79_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[9] == c_79_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[10] == c_79_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[10] == c_79_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[11] == c_79_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[11] == c_79_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[12] == c_79_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[12] == c_79_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[13] == c_79_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[13] == c_79_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[14] == c_79_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[14] == c_79_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[15] == c_79_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[15] == c_79_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[16] == c_79_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[16] == c_79_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[17] == c_79_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[17] == c_79_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[18] == c_79_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[18] == c_79_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[19] == c_79_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[19] == c_79_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[20] == c_79_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[20] == c_79_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[21] == c_79_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[21] == c_79_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[22] == c_79_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[22] == c_79_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[23] == c_79_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[23] == c_79_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[24] == c_79_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[24] == c_79_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[25] == c_79_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[25] == c_79_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[26] == c_79_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[26] == c_79_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[27] == c_79_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[27] == c_79_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[28] == c_79_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[28] == c_79_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[29] == c_79_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[29] == c_79_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[30] == c_79_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[30] == c_79_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[31] == c_79_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[31] == c_79_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_79[32] == c_79_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_79[32] == c_79_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[0] == c_80_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[0] == c_80_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[1] == c_80_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[1] == c_80_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[2] == c_80_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[2] == c_80_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[3] == c_80_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[3] == c_80_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[4] == c_80_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[4] == c_80_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[5] == c_80_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[5] == c_80_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[6] == c_80_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[6] == c_80_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[7] == c_80_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[7] == c_80_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[8] == c_80_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[8] == c_80_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[9] == c_80_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[9] == c_80_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[10] == c_80_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[10] == c_80_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[11] == c_80_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[11] == c_80_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[12] == c_80_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[12] == c_80_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[13] == c_80_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[13] == c_80_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[14] == c_80_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[14] == c_80_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[15] == c_80_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[15] == c_80_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[16] == c_80_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[16] == c_80_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[17] == c_80_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[17] == c_80_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[18] == c_80_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[18] == c_80_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[19] == c_80_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[19] == c_80_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[20] == c_80_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[20] == c_80_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[21] == c_80_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[21] == c_80_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[22] == c_80_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[22] == c_80_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[23] == c_80_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[23] == c_80_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[24] == c_80_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[24] == c_80_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[25] == c_80_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[25] == c_80_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[26] == c_80_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[26] == c_80_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[27] == c_80_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[27] == c_80_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[28] == c_80_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[28] == c_80_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[29] == c_80_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[29] == c_80_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[30] == c_80_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[30] == c_80_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[31] == c_80_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[31] == c_80_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_80[32] == c_80_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_80[32] == c_80_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[0] == c_81_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[0] == c_81_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[1] == c_81_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[1] == c_81_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[2] == c_81_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[2] == c_81_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[3] == c_81_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[3] == c_81_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[4] == c_81_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[4] == c_81_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[5] == c_81_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[5] == c_81_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[6] == c_81_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[6] == c_81_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[7] == c_81_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[7] == c_81_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[8] == c_81_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[8] == c_81_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[9] == c_81_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[9] == c_81_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[10] == c_81_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[10] == c_81_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[11] == c_81_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[11] == c_81_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[12] == c_81_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[12] == c_81_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[13] == c_81_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[13] == c_81_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[14] == c_81_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[14] == c_81_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[15] == c_81_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[15] == c_81_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[16] == c_81_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[16] == c_81_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[17] == c_81_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[17] == c_81_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[18] == c_81_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[18] == c_81_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[19] == c_81_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[19] == c_81_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[20] == c_81_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[20] == c_81_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[21] == c_81_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[21] == c_81_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[22] == c_81_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[22] == c_81_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[23] == c_81_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[23] == c_81_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[24] == c_81_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[24] == c_81_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[25] == c_81_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[25] == c_81_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[26] == c_81_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[26] == c_81_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[27] == c_81_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[27] == c_81_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[28] == c_81_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[28] == c_81_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[29] == c_81_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[29] == c_81_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[30] == c_81_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[30] == c_81_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[31] == c_81_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[31] == c_81_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_81[32] == c_81_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_81[32] == c_81_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[0] == c_82_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[0] == c_82_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[1] == c_82_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[1] == c_82_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[2] == c_82_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[2] == c_82_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[3] == c_82_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[3] == c_82_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[4] == c_82_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[4] == c_82_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[5] == c_82_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[5] == c_82_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[6] == c_82_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[6] == c_82_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[7] == c_82_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[7] == c_82_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[8] == c_82_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[8] == c_82_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[9] == c_82_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[9] == c_82_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[10] == c_82_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[10] == c_82_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[11] == c_82_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[11] == c_82_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[12] == c_82_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[12] == c_82_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[13] == c_82_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[13] == c_82_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[14] == c_82_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[14] == c_82_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[15] == c_82_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[15] == c_82_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[16] == c_82_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[16] == c_82_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[17] == c_82_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[17] == c_82_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[18] == c_82_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[18] == c_82_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[19] == c_82_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[19] == c_82_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[20] == c_82_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[20] == c_82_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[21] == c_82_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[21] == c_82_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[22] == c_82_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[22] == c_82_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[23] == c_82_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[23] == c_82_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[24] == c_82_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[24] == c_82_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[25] == c_82_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[25] == c_82_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[26] == c_82_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[26] == c_82_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[27] == c_82_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[27] == c_82_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[28] == c_82_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[28] == c_82_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[29] == c_82_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[29] == c_82_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[30] == c_82_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[30] == c_82_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[31] == c_82_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[31] == c_82_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_82[32] == c_82_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_82[32] == c_82_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[0] == c_83_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[0] == c_83_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[1] == c_83_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[1] == c_83_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[2] == c_83_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[2] == c_83_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[3] == c_83_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[3] == c_83_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[4] == c_83_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[4] == c_83_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[5] == c_83_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[5] == c_83_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[6] == c_83_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[6] == c_83_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[7] == c_83_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[7] == c_83_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[8] == c_83_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[8] == c_83_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[9] == c_83_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[9] == c_83_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[10] == c_83_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[10] == c_83_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[11] == c_83_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[11] == c_83_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[12] == c_83_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[12] == c_83_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[13] == c_83_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[13] == c_83_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[14] == c_83_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[14] == c_83_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[15] == c_83_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[15] == c_83_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[16] == c_83_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[16] == c_83_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[17] == c_83_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[17] == c_83_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[18] == c_83_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[18] == c_83_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[19] == c_83_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[19] == c_83_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[20] == c_83_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[20] == c_83_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[21] == c_83_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[21] == c_83_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[22] == c_83_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[22] == c_83_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[23] == c_83_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[23] == c_83_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[24] == c_83_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[24] == c_83_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[25] == c_83_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[25] == c_83_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[26] == c_83_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[26] == c_83_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[27] == c_83_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[27] == c_83_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[28] == c_83_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[28] == c_83_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[29] == c_83_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[29] == c_83_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[30] == c_83_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[30] == c_83_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[31] == c_83_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[31] == c_83_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_83[32] == c_83_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_83[32] == c_83_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[0] == c_84_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[0] == c_84_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[1] == c_84_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[1] == c_84_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[2] == c_84_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[2] == c_84_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[3] == c_84_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[3] == c_84_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[4] == c_84_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[4] == c_84_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[5] == c_84_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[5] == c_84_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[6] == c_84_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[6] == c_84_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[7] == c_84_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[7] == c_84_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[8] == c_84_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[8] == c_84_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[9] == c_84_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[9] == c_84_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[10] == c_84_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[10] == c_84_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[11] == c_84_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[11] == c_84_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[12] == c_84_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[12] == c_84_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[13] == c_84_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[13] == c_84_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[14] == c_84_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[14] == c_84_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[15] == c_84_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[15] == c_84_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[16] == c_84_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[16] == c_84_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[17] == c_84_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[17] == c_84_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[18] == c_84_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[18] == c_84_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[19] == c_84_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[19] == c_84_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[20] == c_84_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[20] == c_84_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[21] == c_84_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[21] == c_84_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[22] == c_84_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[22] == c_84_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[23] == c_84_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[23] == c_84_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[24] == c_84_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[24] == c_84_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[25] == c_84_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[25] == c_84_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[26] == c_84_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[26] == c_84_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[27] == c_84_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[27] == c_84_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[28] == c_84_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[28] == c_84_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[29] == c_84_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[29] == c_84_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[30] == c_84_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[30] == c_84_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[31] == c_84_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[31] == c_84_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_84[32] == c_84_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_84[32] == c_84_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[0] == c_85_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[0] == c_85_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[1] == c_85_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[1] == c_85_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[2] == c_85_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[2] == c_85_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[3] == c_85_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[3] == c_85_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[4] == c_85_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[4] == c_85_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[5] == c_85_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[5] == c_85_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[6] == c_85_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[6] == c_85_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[7] == c_85_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[7] == c_85_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[8] == c_85_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[8] == c_85_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[9] == c_85_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[9] == c_85_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[10] == c_85_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[10] == c_85_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[11] == c_85_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[11] == c_85_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[12] == c_85_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[12] == c_85_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[13] == c_85_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[13] == c_85_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[14] == c_85_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[14] == c_85_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[15] == c_85_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[15] == c_85_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[16] == c_85_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[16] == c_85_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[17] == c_85_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[17] == c_85_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[18] == c_85_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[18] == c_85_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[19] == c_85_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[19] == c_85_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[20] == c_85_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[20] == c_85_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[21] == c_85_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[21] == c_85_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[22] == c_85_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[22] == c_85_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[23] == c_85_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[23] == c_85_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[24] == c_85_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[24] == c_85_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[25] == c_85_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[25] == c_85_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[26] == c_85_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[26] == c_85_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[27] == c_85_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[27] == c_85_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[28] == c_85_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[28] == c_85_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[29] == c_85_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[29] == c_85_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[30] == c_85_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[30] == c_85_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[31] == c_85_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[31] == c_85_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_85[32] == c_85_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_85[32] == c_85_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[0] == c_86_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[0] == c_86_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[1] == c_86_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[1] == c_86_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[2] == c_86_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[2] == c_86_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[3] == c_86_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[3] == c_86_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[4] == c_86_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[4] == c_86_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[5] == c_86_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[5] == c_86_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[6] == c_86_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[6] == c_86_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[7] == c_86_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[7] == c_86_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[8] == c_86_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[8] == c_86_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[9] == c_86_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[9] == c_86_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[10] == c_86_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[10] == c_86_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[11] == c_86_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[11] == c_86_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[12] == c_86_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[12] == c_86_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[13] == c_86_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[13] == c_86_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[14] == c_86_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[14] == c_86_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[15] == c_86_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[15] == c_86_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[16] == c_86_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[16] == c_86_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[17] == c_86_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[17] == c_86_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[18] == c_86_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[18] == c_86_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[19] == c_86_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[19] == c_86_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[20] == c_86_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[20] == c_86_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[21] == c_86_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[21] == c_86_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[22] == c_86_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[22] == c_86_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[23] == c_86_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[23] == c_86_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[24] == c_86_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[24] == c_86_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[25] == c_86_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[25] == c_86_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[26] == c_86_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[26] == c_86_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[27] == c_86_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[27] == c_86_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[28] == c_86_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[28] == c_86_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[29] == c_86_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[29] == c_86_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[30] == c_86_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[30] == c_86_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[31] == c_86_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[31] == c_86_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_86[32] == c_86_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_86[32] == c_86_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[0] == c_87_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[0] == c_87_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[1] == c_87_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[1] == c_87_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[2] == c_87_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[2] == c_87_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[3] == c_87_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[3] == c_87_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[4] == c_87_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[4] == c_87_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[5] == c_87_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[5] == c_87_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[6] == c_87_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[6] == c_87_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[7] == c_87_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[7] == c_87_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[8] == c_87_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[8] == c_87_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[9] == c_87_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[9] == c_87_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[10] == c_87_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[10] == c_87_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[11] == c_87_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[11] == c_87_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[12] == c_87_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[12] == c_87_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[13] == c_87_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[13] == c_87_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[14] == c_87_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[14] == c_87_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[15] == c_87_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[15] == c_87_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[16] == c_87_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[16] == c_87_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[17] == c_87_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[17] == c_87_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[18] == c_87_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[18] == c_87_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[19] == c_87_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[19] == c_87_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[20] == c_87_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[20] == c_87_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[21] == c_87_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[21] == c_87_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[22] == c_87_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[22] == c_87_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[23] == c_87_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[23] == c_87_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[24] == c_87_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[24] == c_87_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[25] == c_87_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[25] == c_87_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[26] == c_87_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[26] == c_87_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[27] == c_87_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[27] == c_87_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[28] == c_87_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[28] == c_87_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[29] == c_87_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[29] == c_87_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[30] == c_87_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[30] == c_87_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[31] == c_87_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[31] == c_87_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_87[32] == c_87_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_87[32] == c_87_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[0] == c_88_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[0] == c_88_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[1] == c_88_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[1] == c_88_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[2] == c_88_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[2] == c_88_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[3] == c_88_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[3] == c_88_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[4] == c_88_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[4] == c_88_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[5] == c_88_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[5] == c_88_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[6] == c_88_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[6] == c_88_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[7] == c_88_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[7] == c_88_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[8] == c_88_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[8] == c_88_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[9] == c_88_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[9] == c_88_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[10] == c_88_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[10] == c_88_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[11] == c_88_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[11] == c_88_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[12] == c_88_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[12] == c_88_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[13] == c_88_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[13] == c_88_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[14] == c_88_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[14] == c_88_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[15] == c_88_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[15] == c_88_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[16] == c_88_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[16] == c_88_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[17] == c_88_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[17] == c_88_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[18] == c_88_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[18] == c_88_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[19] == c_88_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[19] == c_88_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[20] == c_88_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[20] == c_88_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[21] == c_88_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[21] == c_88_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[22] == c_88_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[22] == c_88_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[23] == c_88_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[23] == c_88_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[24] == c_88_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[24] == c_88_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[25] == c_88_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[25] == c_88_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[26] == c_88_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[26] == c_88_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[27] == c_88_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[27] == c_88_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[28] == c_88_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[28] == c_88_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[29] == c_88_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[29] == c_88_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[30] == c_88_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[30] == c_88_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[31] == c_88_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[31] == c_88_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_88[32] == c_88_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_88[32] == c_88_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[0] == c_89_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[0] == c_89_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[1] == c_89_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[1] == c_89_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[2] == c_89_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[2] == c_89_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[3] == c_89_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[3] == c_89_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[4] == c_89_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[4] == c_89_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[5] == c_89_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[5] == c_89_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[6] == c_89_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[6] == c_89_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[7] == c_89_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[7] == c_89_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[8] == c_89_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[8] == c_89_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[9] == c_89_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[9] == c_89_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[10] == c_89_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[10] == c_89_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[11] == c_89_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[11] == c_89_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[12] == c_89_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[12] == c_89_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[13] == c_89_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[13] == c_89_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[14] == c_89_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[14] == c_89_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[15] == c_89_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[15] == c_89_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[16] == c_89_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[16] == c_89_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[17] == c_89_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[17] == c_89_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[18] == c_89_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[18] == c_89_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[19] == c_89_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[19] == c_89_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[20] == c_89_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[20] == c_89_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[21] == c_89_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[21] == c_89_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[22] == c_89_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[22] == c_89_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[23] == c_89_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[23] == c_89_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[24] == c_89_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[24] == c_89_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[25] == c_89_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[25] == c_89_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[26] == c_89_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[26] == c_89_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[27] == c_89_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[27] == c_89_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[28] == c_89_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[28] == c_89_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[29] == c_89_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[29] == c_89_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[30] == c_89_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[30] == c_89_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[31] == c_89_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[31] == c_89_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_89[32] == c_89_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_89[32] == c_89_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[0] == c_90_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[0] == c_90_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[1] == c_90_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[1] == c_90_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[2] == c_90_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[2] == c_90_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[3] == c_90_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[3] == c_90_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[4] == c_90_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[4] == c_90_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[5] == c_90_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[5] == c_90_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[6] == c_90_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[6] == c_90_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[7] == c_90_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[7] == c_90_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[8] == c_90_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[8] == c_90_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[9] == c_90_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[9] == c_90_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[10] == c_90_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[10] == c_90_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[11] == c_90_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[11] == c_90_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[12] == c_90_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[12] == c_90_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[13] == c_90_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[13] == c_90_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[14] == c_90_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[14] == c_90_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[15] == c_90_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[15] == c_90_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[16] == c_90_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[16] == c_90_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[17] == c_90_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[17] == c_90_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[18] == c_90_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[18] == c_90_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[19] == c_90_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[19] == c_90_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[20] == c_90_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[20] == c_90_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[21] == c_90_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[21] == c_90_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[22] == c_90_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[22] == c_90_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[23] == c_90_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[23] == c_90_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[24] == c_90_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[24] == c_90_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[25] == c_90_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[25] == c_90_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[26] == c_90_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[26] == c_90_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[27] == c_90_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[27] == c_90_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[28] == c_90_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[28] == c_90_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[29] == c_90_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[29] == c_90_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[30] == c_90_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[30] == c_90_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[31] == c_90_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[31] == c_90_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_90[32] == c_90_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_90[32] == c_90_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[0] == c_91_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[0] == c_91_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[1] == c_91_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[1] == c_91_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[2] == c_91_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[2] == c_91_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[3] == c_91_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[3] == c_91_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[4] == c_91_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[4] == c_91_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[5] == c_91_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[5] == c_91_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[6] == c_91_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[6] == c_91_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[7] == c_91_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[7] == c_91_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[8] == c_91_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[8] == c_91_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[9] == c_91_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[9] == c_91_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[10] == c_91_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[10] == c_91_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[11] == c_91_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[11] == c_91_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[12] == c_91_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[12] == c_91_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[13] == c_91_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[13] == c_91_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[14] == c_91_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[14] == c_91_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[15] == c_91_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[15] == c_91_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[16] == c_91_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[16] == c_91_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[17] == c_91_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[17] == c_91_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[18] == c_91_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[18] == c_91_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[19] == c_91_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[19] == c_91_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[20] == c_91_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[20] == c_91_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[21] == c_91_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[21] == c_91_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[22] == c_91_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[22] == c_91_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[23] == c_91_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[23] == c_91_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[24] == c_91_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[24] == c_91_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[25] == c_91_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[25] == c_91_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[26] == c_91_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[26] == c_91_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[27] == c_91_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[27] == c_91_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[28] == c_91_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[28] == c_91_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[29] == c_91_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[29] == c_91_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[30] == c_91_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[30] == c_91_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[31] == c_91_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[31] == c_91_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_91[32] == c_91_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_91[32] == c_91_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[0] == c_92_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[0] == c_92_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[1] == c_92_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[1] == c_92_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[2] == c_92_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[2] == c_92_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[3] == c_92_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[3] == c_92_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[4] == c_92_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[4] == c_92_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[5] == c_92_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[5] == c_92_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[6] == c_92_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[6] == c_92_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[7] == c_92_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[7] == c_92_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[8] == c_92_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[8] == c_92_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[9] == c_92_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[9] == c_92_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[10] == c_92_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[10] == c_92_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[11] == c_92_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[11] == c_92_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[12] == c_92_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[12] == c_92_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[13] == c_92_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[13] == c_92_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[14] == c_92_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[14] == c_92_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[15] == c_92_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[15] == c_92_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[16] == c_92_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[16] == c_92_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[17] == c_92_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[17] == c_92_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[18] == c_92_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[18] == c_92_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[19] == c_92_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[19] == c_92_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[20] == c_92_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[20] == c_92_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[21] == c_92_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[21] == c_92_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[22] == c_92_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[22] == c_92_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[23] == c_92_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[23] == c_92_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[24] == c_92_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[24] == c_92_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[25] == c_92_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[25] == c_92_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[26] == c_92_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[26] == c_92_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[27] == c_92_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[27] == c_92_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[28] == c_92_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[28] == c_92_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[29] == c_92_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[29] == c_92_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[30] == c_92_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[30] == c_92_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[31] == c_92_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[31] == c_92_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_92[32] == c_92_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_92[32] == c_92_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[0] == c_93_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[0] == c_93_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[1] == c_93_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[1] == c_93_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[2] == c_93_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[2] == c_93_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[3] == c_93_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[3] == c_93_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[4] == c_93_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[4] == c_93_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[5] == c_93_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[5] == c_93_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[6] == c_93_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[6] == c_93_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[7] == c_93_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[7] == c_93_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[8] == c_93_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[8] == c_93_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[9] == c_93_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[9] == c_93_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[10] == c_93_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[10] == c_93_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[11] == c_93_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[11] == c_93_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[12] == c_93_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[12] == c_93_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[13] == c_93_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[13] == c_93_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[14] == c_93_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[14] == c_93_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[15] == c_93_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[15] == c_93_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[16] == c_93_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[16] == c_93_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[17] == c_93_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[17] == c_93_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[18] == c_93_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[18] == c_93_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[19] == c_93_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[19] == c_93_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[20] == c_93_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[20] == c_93_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[21] == c_93_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[21] == c_93_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[22] == c_93_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[22] == c_93_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[23] == c_93_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[23] == c_93_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[24] == c_93_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[24] == c_93_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[25] == c_93_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[25] == c_93_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[26] == c_93_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[26] == c_93_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[27] == c_93_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[27] == c_93_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[28] == c_93_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[28] == c_93_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[29] == c_93_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[29] == c_93_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[30] == c_93_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[30] == c_93_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[31] == c_93_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[31] == c_93_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_93[32] == c_93_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_93[32] == c_93_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[0] == c_94_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[0] == c_94_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[1] == c_94_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[1] == c_94_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[2] == c_94_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[2] == c_94_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[3] == c_94_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[3] == c_94_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[4] == c_94_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[4] == c_94_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[5] == c_94_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[5] == c_94_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[6] == c_94_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[6] == c_94_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[7] == c_94_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[7] == c_94_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[8] == c_94_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[8] == c_94_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[9] == c_94_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[9] == c_94_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[10] == c_94_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[10] == c_94_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[11] == c_94_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[11] == c_94_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[12] == c_94_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[12] == c_94_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[13] == c_94_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[13] == c_94_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[14] == c_94_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[14] == c_94_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[15] == c_94_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[15] == c_94_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[16] == c_94_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[16] == c_94_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[17] == c_94_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[17] == c_94_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[18] == c_94_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[18] == c_94_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[19] == c_94_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[19] == c_94_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[20] == c_94_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[20] == c_94_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[21] == c_94_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[21] == c_94_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[22] == c_94_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[22] == c_94_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[23] == c_94_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[23] == c_94_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[24] == c_94_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[24] == c_94_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[25] == c_94_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[25] == c_94_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[26] == c_94_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[26] == c_94_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[27] == c_94_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[27] == c_94_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[28] == c_94_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[28] == c_94_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[29] == c_94_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[29] == c_94_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[30] == c_94_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[30] == c_94_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[31] == c_94_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[31] == c_94_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_94[32] == c_94_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_94[32] == c_94_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[0] == c_95_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[0] == c_95_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[1] == c_95_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[1] == c_95_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[2] == c_95_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[2] == c_95_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[3] == c_95_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[3] == c_95_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[4] == c_95_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[4] == c_95_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[5] == c_95_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[5] == c_95_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[6] == c_95_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[6] == c_95_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[7] == c_95_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[7] == c_95_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[8] == c_95_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[8] == c_95_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[9] == c_95_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[9] == c_95_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[10] == c_95_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[10] == c_95_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[11] == c_95_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[11] == c_95_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[12] == c_95_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[12] == c_95_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[13] == c_95_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[13] == c_95_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[14] == c_95_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[14] == c_95_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[15] == c_95_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[15] == c_95_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[16] == c_95_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[16] == c_95_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[17] == c_95_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[17] == c_95_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[18] == c_95_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[18] == c_95_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[19] == c_95_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[19] == c_95_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[20] == c_95_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[20] == c_95_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[21] == c_95_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[21] == c_95_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[22] == c_95_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[22] == c_95_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[23] == c_95_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[23] == c_95_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[24] == c_95_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[24] == c_95_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[25] == c_95_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[25] == c_95_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[26] == c_95_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[26] == c_95_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[27] == c_95_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[27] == c_95_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[28] == c_95_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[28] == c_95_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[29] == c_95_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[29] == c_95_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[30] == c_95_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[30] == c_95_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[31] == c_95_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[31] == c_95_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_95[32] == c_95_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_95[32] == c_95_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[0] == c_96_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[0] == c_96_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[1] == c_96_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[1] == c_96_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[2] == c_96_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[2] == c_96_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[3] == c_96_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[3] == c_96_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[4] == c_96_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[4] == c_96_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[5] == c_96_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[5] == c_96_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[6] == c_96_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[6] == c_96_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[7] == c_96_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[7] == c_96_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[8] == c_96_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[8] == c_96_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[9] == c_96_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[9] == c_96_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[10] == c_96_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[10] == c_96_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[11] == c_96_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[11] == c_96_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[12] == c_96_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[12] == c_96_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[13] == c_96_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[13] == c_96_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[14] == c_96_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[14] == c_96_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[15] == c_96_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[15] == c_96_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[16] == c_96_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[16] == c_96_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[17] == c_96_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[17] == c_96_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[18] == c_96_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[18] == c_96_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[19] == c_96_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[19] == c_96_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[20] == c_96_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[20] == c_96_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[21] == c_96_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[21] == c_96_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[22] == c_96_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[22] == c_96_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[23] == c_96_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[23] == c_96_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[24] == c_96_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[24] == c_96_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[25] == c_96_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[25] == c_96_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[26] == c_96_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[26] == c_96_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[27] == c_96_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[27] == c_96_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[28] == c_96_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[28] == c_96_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[29] == c_96_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[29] == c_96_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[30] == c_96_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[30] == c_96_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[31] == c_96_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[31] == c_96_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_96[32] == c_96_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_96[32] == c_96_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[0] == c_97_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[0] == c_97_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[1] == c_97_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[1] == c_97_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[2] == c_97_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[2] == c_97_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[3] == c_97_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[3] == c_97_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[4] == c_97_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[4] == c_97_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[5] == c_97_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[5] == c_97_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[6] == c_97_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[6] == c_97_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[7] == c_97_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[7] == c_97_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[8] == c_97_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[8] == c_97_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[9] == c_97_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[9] == c_97_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[10] == c_97_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[10] == c_97_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[11] == c_97_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[11] == c_97_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[12] == c_97_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[12] == c_97_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[13] == c_97_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[13] == c_97_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[14] == c_97_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[14] == c_97_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[15] == c_97_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[15] == c_97_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[16] == c_97_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[16] == c_97_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[17] == c_97_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[17] == c_97_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[18] == c_97_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[18] == c_97_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[19] == c_97_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[19] == c_97_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[20] == c_97_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[20] == c_97_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[21] == c_97_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[21] == c_97_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[22] == c_97_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[22] == c_97_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[23] == c_97_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[23] == c_97_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[24] == c_97_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[24] == c_97_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[25] == c_97_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[25] == c_97_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[26] == c_97_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[26] == c_97_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[27] == c_97_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[27] == c_97_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[28] == c_97_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[28] == c_97_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[29] == c_97_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[29] == c_97_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[30] == c_97_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[30] == c_97_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[31] == c_97_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[31] == c_97_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_97[32] == c_97_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_97[32] == c_97_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[0] == c_98_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[0] == c_98_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[1] == c_98_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[1] == c_98_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[2] == c_98_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[2] == c_98_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[3] == c_98_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[3] == c_98_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[4] == c_98_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[4] == c_98_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[5] == c_98_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[5] == c_98_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[6] == c_98_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[6] == c_98_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[7] == c_98_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[7] == c_98_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[8] == c_98_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[8] == c_98_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[9] == c_98_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[9] == c_98_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[10] == c_98_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[10] == c_98_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[11] == c_98_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[11] == c_98_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[12] == c_98_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[12] == c_98_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[13] == c_98_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[13] == c_98_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[14] == c_98_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[14] == c_98_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[15] == c_98_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[15] == c_98_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[16] == c_98_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[16] == c_98_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[17] == c_98_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[17] == c_98_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[18] == c_98_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[18] == c_98_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[19] == c_98_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[19] == c_98_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[20] == c_98_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[20] == c_98_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[21] == c_98_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[21] == c_98_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[22] == c_98_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[22] == c_98_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[23] == c_98_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[23] == c_98_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[24] == c_98_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[24] == c_98_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[25] == c_98_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[25] == c_98_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[26] == c_98_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[26] == c_98_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[27] == c_98_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[27] == c_98_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[28] == c_98_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[28] == c_98_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[29] == c_98_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[29] == c_98_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[30] == c_98_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[30] == c_98_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[31] == c_98_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[31] == c_98_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_98[32] == c_98_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_98[32] == c_98_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[0] == c_99_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[0] == c_99_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[1] == c_99_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[1] == c_99_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[2] == c_99_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[2] == c_99_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[3] == c_99_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[3] == c_99_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[4] == c_99_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[4] == c_99_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[5] == c_99_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[5] == c_99_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[6] == c_99_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[6] == c_99_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[7] == c_99_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[7] == c_99_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[8] == c_99_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[8] == c_99_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[9] == c_99_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[9] == c_99_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[10] == c_99_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[10] == c_99_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[11] == c_99_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[11] == c_99_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[12] == c_99_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[12] == c_99_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[13] == c_99_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[13] == c_99_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[14] == c_99_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[14] == c_99_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[15] == c_99_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[15] == c_99_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[16] == c_99_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[16] == c_99_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[17] == c_99_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[17] == c_99_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[18] == c_99_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[18] == c_99_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[19] == c_99_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[19] == c_99_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[20] == c_99_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[20] == c_99_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[21] == c_99_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[21] == c_99_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[22] == c_99_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[22] == c_99_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[23] == c_99_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[23] == c_99_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[24] == c_99_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[24] == c_99_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[25] == c_99_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[25] == c_99_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[26] == c_99_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[26] == c_99_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[27] == c_99_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[27] == c_99_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[28] == c_99_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[28] == c_99_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[29] == c_99_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[29] == c_99_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[30] == c_99_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[30] == c_99_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[31] == c_99_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[31] == c_99_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_99[32] == c_99_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_99[32] == c_99_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[0] == c_100_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[0] == c_100_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[1] == c_100_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[1] == c_100_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[2] == c_100_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[2] == c_100_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[3] == c_100_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[3] == c_100_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[4] == c_100_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[4] == c_100_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[5] == c_100_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[5] == c_100_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[6] == c_100_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[6] == c_100_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[7] == c_100_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[7] == c_100_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[8] == c_100_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[8] == c_100_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[9] == c_100_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[9] == c_100_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[10] == c_100_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[10] == c_100_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[11] == c_100_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[11] == c_100_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[12] == c_100_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[12] == c_100_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[13] == c_100_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[13] == c_100_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[14] == c_100_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[14] == c_100_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[15] == c_100_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[15] == c_100_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[16] == c_100_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[16] == c_100_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[17] == c_100_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[17] == c_100_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[18] == c_100_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[18] == c_100_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[19] == c_100_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[19] == c_100_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[20] == c_100_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[20] == c_100_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[21] == c_100_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[21] == c_100_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[22] == c_100_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[22] == c_100_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[23] == c_100_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[23] == c_100_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[24] == c_100_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[24] == c_100_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[25] == c_100_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[25] == c_100_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[26] == c_100_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[26] == c_100_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[27] == c_100_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[27] == c_100_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[28] == c_100_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[28] == c_100_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[29] == c_100_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[29] == c_100_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[30] == c_100_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[30] == c_100_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[31] == c_100_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[31] == c_100_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_100[32] == c_100_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_100[32] == c_100_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[0] == c_101_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[0] == c_101_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[1] == c_101_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[1] == c_101_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[2] == c_101_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[2] == c_101_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[3] == c_101_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[3] == c_101_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[4] == c_101_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[4] == c_101_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[5] == c_101_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[5] == c_101_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[6] == c_101_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[6] == c_101_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[7] == c_101_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[7] == c_101_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[8] == c_101_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[8] == c_101_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[9] == c_101_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[9] == c_101_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[10] == c_101_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[10] == c_101_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[11] == c_101_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[11] == c_101_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[12] == c_101_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[12] == c_101_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[13] == c_101_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[13] == c_101_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[14] == c_101_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[14] == c_101_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[15] == c_101_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[15] == c_101_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[16] == c_101_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[16] == c_101_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[17] == c_101_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[17] == c_101_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[18] == c_101_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[18] == c_101_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[19] == c_101_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[19] == c_101_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[20] == c_101_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[20] == c_101_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[21] == c_101_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[21] == c_101_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[22] == c_101_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[22] == c_101_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[23] == c_101_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[23] == c_101_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[24] == c_101_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[24] == c_101_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[25] == c_101_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[25] == c_101_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[26] == c_101_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[26] == c_101_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[27] == c_101_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[27] == c_101_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[28] == c_101_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[28] == c_101_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[29] == c_101_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[29] == c_101_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[30] == c_101_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[30] == c_101_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[31] == c_101_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[31] == c_101_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_101[32] == c_101_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_101[32] == c_101_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[0] == c_102_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[0] == c_102_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[1] == c_102_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[1] == c_102_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[2] == c_102_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[2] == c_102_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[3] == c_102_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[3] == c_102_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[4] == c_102_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[4] == c_102_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[5] == c_102_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[5] == c_102_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[6] == c_102_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[6] == c_102_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[7] == c_102_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[7] == c_102_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[8] == c_102_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[8] == c_102_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[9] == c_102_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[9] == c_102_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[10] == c_102_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[10] == c_102_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[11] == c_102_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[11] == c_102_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[12] == c_102_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[12] == c_102_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[13] == c_102_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[13] == c_102_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[14] == c_102_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[14] == c_102_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[15] == c_102_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[15] == c_102_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[16] == c_102_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[16] == c_102_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[17] == c_102_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[17] == c_102_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[18] == c_102_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[18] == c_102_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[19] == c_102_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[19] == c_102_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[20] == c_102_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[20] == c_102_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[21] == c_102_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[21] == c_102_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[22] == c_102_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[22] == c_102_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[23] == c_102_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[23] == c_102_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[24] == c_102_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[24] == c_102_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[25] == c_102_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[25] == c_102_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[26] == c_102_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[26] == c_102_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[27] == c_102_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[27] == c_102_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[28] == c_102_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[28] == c_102_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[29] == c_102_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[29] == c_102_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[30] == c_102_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[30] == c_102_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[31] == c_102_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[31] == c_102_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_102[32] == c_102_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_102[32] == c_102_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[0] == c_103_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[0] == c_103_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[1] == c_103_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[1] == c_103_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[2] == c_103_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[2] == c_103_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[3] == c_103_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[3] == c_103_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[4] == c_103_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[4] == c_103_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[5] == c_103_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[5] == c_103_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[6] == c_103_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[6] == c_103_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[7] == c_103_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[7] == c_103_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[8] == c_103_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[8] == c_103_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[9] == c_103_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[9] == c_103_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[10] == c_103_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[10] == c_103_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[11] == c_103_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[11] == c_103_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[12] == c_103_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[12] == c_103_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[13] == c_103_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[13] == c_103_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[14] == c_103_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[14] == c_103_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[15] == c_103_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[15] == c_103_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[16] == c_103_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[16] == c_103_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[17] == c_103_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[17] == c_103_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[18] == c_103_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[18] == c_103_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[19] == c_103_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[19] == c_103_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[20] == c_103_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[20] == c_103_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[21] == c_103_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[21] == c_103_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[22] == c_103_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[22] == c_103_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[23] == c_103_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[23] == c_103_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[24] == c_103_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[24] == c_103_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[25] == c_103_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[25] == c_103_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[26] == c_103_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[26] == c_103_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[27] == c_103_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[27] == c_103_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[28] == c_103_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[28] == c_103_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[29] == c_103_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[29] == c_103_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[30] == c_103_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[30] == c_103_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[31] == c_103_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[31] == c_103_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_103[32] == c_103_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_103[32] == c_103_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[0] == c_104_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[0] == c_104_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[1] == c_104_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[1] == c_104_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[2] == c_104_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[2] == c_104_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[3] == c_104_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[3] == c_104_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[4] == c_104_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[4] == c_104_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[5] == c_104_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[5] == c_104_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[6] == c_104_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[6] == c_104_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[7] == c_104_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[7] == c_104_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[8] == c_104_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[8] == c_104_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[9] == c_104_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[9] == c_104_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[10] == c_104_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[10] == c_104_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[11] == c_104_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[11] == c_104_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[12] == c_104_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[12] == c_104_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[13] == c_104_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[13] == c_104_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[14] == c_104_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[14] == c_104_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[15] == c_104_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[15] == c_104_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[16] == c_104_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[16] == c_104_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[17] == c_104_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[17] == c_104_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[18] == c_104_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[18] == c_104_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[19] == c_104_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[19] == c_104_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[20] == c_104_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[20] == c_104_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[21] == c_104_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[21] == c_104_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[22] == c_104_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[22] == c_104_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[23] == c_104_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[23] == c_104_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[24] == c_104_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[24] == c_104_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[25] == c_104_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[25] == c_104_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[26] == c_104_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[26] == c_104_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[27] == c_104_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[27] == c_104_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[28] == c_104_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[28] == c_104_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[29] == c_104_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[29] == c_104_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[30] == c_104_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[30] == c_104_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[31] == c_104_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[31] == c_104_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_104[32] == c_104_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_104[32] == c_104_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[0] == c_105_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[0] == c_105_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[1] == c_105_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[1] == c_105_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[2] == c_105_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[2] == c_105_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[3] == c_105_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[3] == c_105_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[4] == c_105_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[4] == c_105_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[5] == c_105_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[5] == c_105_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[6] == c_105_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[6] == c_105_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[7] == c_105_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[7] == c_105_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[8] == c_105_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[8] == c_105_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[9] == c_105_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[9] == c_105_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[10] == c_105_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[10] == c_105_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[11] == c_105_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[11] == c_105_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[12] == c_105_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[12] == c_105_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[13] == c_105_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[13] == c_105_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[14] == c_105_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[14] == c_105_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[15] == c_105_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[15] == c_105_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[16] == c_105_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[16] == c_105_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[17] == c_105_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[17] == c_105_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[18] == c_105_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[18] == c_105_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[19] == c_105_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[19] == c_105_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[20] == c_105_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[20] == c_105_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[21] == c_105_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[21] == c_105_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[22] == c_105_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[22] == c_105_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[23] == c_105_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[23] == c_105_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[24] == c_105_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[24] == c_105_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[25] == c_105_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[25] == c_105_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[26] == c_105_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[26] == c_105_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[27] == c_105_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[27] == c_105_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[28] == c_105_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[28] == c_105_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[29] == c_105_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[29] == c_105_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[30] == c_105_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[30] == c_105_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[31] == c_105_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[31] == c_105_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_105[32] == c_105_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_105[32] == c_105_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[0] == c_106_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[0] == c_106_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[1] == c_106_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[1] == c_106_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[2] == c_106_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[2] == c_106_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[3] == c_106_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[3] == c_106_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[4] == c_106_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[4] == c_106_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[5] == c_106_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[5] == c_106_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[6] == c_106_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[6] == c_106_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[7] == c_106_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[7] == c_106_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[8] == c_106_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[8] == c_106_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[9] == c_106_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[9] == c_106_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[10] == c_106_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[10] == c_106_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[11] == c_106_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[11] == c_106_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[12] == c_106_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[12] == c_106_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[13] == c_106_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[13] == c_106_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[14] == c_106_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[14] == c_106_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[15] == c_106_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[15] == c_106_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[16] == c_106_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[16] == c_106_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[17] == c_106_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[17] == c_106_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[18] == c_106_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[18] == c_106_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[19] == c_106_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[19] == c_106_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[20] == c_106_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[20] == c_106_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[21] == c_106_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[21] == c_106_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[22] == c_106_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[22] == c_106_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[23] == c_106_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[23] == c_106_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[24] == c_106_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[24] == c_106_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[25] == c_106_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[25] == c_106_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[26] == c_106_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[26] == c_106_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[27] == c_106_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[27] == c_106_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[28] == c_106_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[28] == c_106_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[29] == c_106_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[29] == c_106_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[30] == c_106_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[30] == c_106_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[31] == c_106_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[31] == c_106_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_106[32] == c_106_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_106[32] == c_106_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[0] == c_107_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[0] == c_107_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[1] == c_107_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[1] == c_107_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[2] == c_107_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[2] == c_107_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[3] == c_107_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[3] == c_107_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[4] == c_107_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[4] == c_107_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[5] == c_107_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[5] == c_107_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[6] == c_107_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[6] == c_107_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[7] == c_107_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[7] == c_107_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[8] == c_107_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[8] == c_107_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[9] == c_107_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[9] == c_107_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[10] == c_107_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[10] == c_107_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[11] == c_107_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[11] == c_107_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[12] == c_107_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[12] == c_107_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[13] == c_107_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[13] == c_107_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[14] == c_107_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[14] == c_107_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[15] == c_107_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[15] == c_107_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[16] == c_107_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[16] == c_107_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[17] == c_107_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[17] == c_107_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[18] == c_107_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[18] == c_107_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[19] == c_107_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[19] == c_107_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[20] == c_107_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[20] == c_107_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[21] == c_107_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[21] == c_107_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[22] == c_107_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[22] == c_107_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[23] == c_107_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[23] == c_107_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[24] == c_107_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[24] == c_107_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[25] == c_107_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[25] == c_107_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[26] == c_107_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[26] == c_107_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[27] == c_107_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[27] == c_107_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[28] == c_107_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[28] == c_107_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[29] == c_107_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[29] == c_107_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[30] == c_107_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[30] == c_107_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[31] == c_107_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[31] == c_107_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_107[32] == c_107_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_107[32] == c_107_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[0] == c_108_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[0] == c_108_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[1] == c_108_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[1] == c_108_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[2] == c_108_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[2] == c_108_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[3] == c_108_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[3] == c_108_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[4] == c_108_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[4] == c_108_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[5] == c_108_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[5] == c_108_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[6] == c_108_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[6] == c_108_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[7] == c_108_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[7] == c_108_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[8] == c_108_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[8] == c_108_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[9] == c_108_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[9] == c_108_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[10] == c_108_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[10] == c_108_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[11] == c_108_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[11] == c_108_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[12] == c_108_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[12] == c_108_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[13] == c_108_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[13] == c_108_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[14] == c_108_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[14] == c_108_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[15] == c_108_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[15] == c_108_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[16] == c_108_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[16] == c_108_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[17] == c_108_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[17] == c_108_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[18] == c_108_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[18] == c_108_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[19] == c_108_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[19] == c_108_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[20] == c_108_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[20] == c_108_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[21] == c_108_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[21] == c_108_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[22] == c_108_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[22] == c_108_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[23] == c_108_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[23] == c_108_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[24] == c_108_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[24] == c_108_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[25] == c_108_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[25] == c_108_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[26] == c_108_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[26] == c_108_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[27] == c_108_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[27] == c_108_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[28] == c_108_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[28] == c_108_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[29] == c_108_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[29] == c_108_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[30] == c_108_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[30] == c_108_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[31] == c_108_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[31] == c_108_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_108[32] == c_108_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_108[32] == c_108_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[0] == c_109_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[0] == c_109_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[1] == c_109_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[1] == c_109_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[2] == c_109_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[2] == c_109_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[3] == c_109_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[3] == c_109_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[4] == c_109_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[4] == c_109_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[5] == c_109_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[5] == c_109_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[6] == c_109_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[6] == c_109_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[7] == c_109_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[7] == c_109_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[8] == c_109_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[8] == c_109_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[9] == c_109_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[9] == c_109_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[10] == c_109_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[10] == c_109_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[11] == c_109_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[11] == c_109_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[12] == c_109_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[12] == c_109_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[13] == c_109_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[13] == c_109_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[14] == c_109_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[14] == c_109_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[15] == c_109_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[15] == c_109_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[16] == c_109_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[16] == c_109_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[17] == c_109_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[17] == c_109_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[18] == c_109_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[18] == c_109_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[19] == c_109_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[19] == c_109_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[20] == c_109_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[20] == c_109_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[21] == c_109_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[21] == c_109_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[22] == c_109_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[22] == c_109_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[23] == c_109_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[23] == c_109_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[24] == c_109_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[24] == c_109_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[25] == c_109_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[25] == c_109_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[26] == c_109_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[26] == c_109_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[27] == c_109_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[27] == c_109_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[28] == c_109_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[28] == c_109_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[29] == c_109_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[29] == c_109_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[30] == c_109_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[30] == c_109_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[31] == c_109_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[31] == c_109_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_109[32] == c_109_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_109[32] == c_109_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[0] == c_110_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[0] == c_110_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[1] == c_110_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[1] == c_110_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[2] == c_110_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[2] == c_110_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[3] == c_110_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[3] == c_110_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[4] == c_110_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[4] == c_110_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[5] == c_110_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[5] == c_110_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[6] == c_110_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[6] == c_110_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[7] == c_110_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[7] == c_110_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[8] == c_110_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[8] == c_110_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[9] == c_110_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[9] == c_110_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[10] == c_110_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[10] == c_110_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[11] == c_110_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[11] == c_110_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[12] == c_110_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[12] == c_110_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[13] == c_110_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[13] == c_110_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[14] == c_110_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[14] == c_110_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[15] == c_110_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[15] == c_110_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[16] == c_110_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[16] == c_110_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[17] == c_110_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[17] == c_110_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[18] == c_110_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[18] == c_110_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[19] == c_110_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[19] == c_110_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[20] == c_110_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[20] == c_110_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[21] == c_110_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[21] == c_110_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[22] == c_110_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[22] == c_110_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[23] == c_110_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[23] == c_110_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[24] == c_110_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[24] == c_110_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[25] == c_110_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[25] == c_110_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[26] == c_110_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[26] == c_110_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[27] == c_110_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[27] == c_110_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[28] == c_110_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[28] == c_110_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[29] == c_110_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[29] == c_110_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[30] == c_110_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[30] == c_110_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[31] == c_110_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[31] == c_110_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_110[32] == c_110_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_110[32] == c_110_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[0] == c_111_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[0] == c_111_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[1] == c_111_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[1] == c_111_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[2] == c_111_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[2] == c_111_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[3] == c_111_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[3] == c_111_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[4] == c_111_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[4] == c_111_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[5] == c_111_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[5] == c_111_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[6] == c_111_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[6] == c_111_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[7] == c_111_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[7] == c_111_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[8] == c_111_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[8] == c_111_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[9] == c_111_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[9] == c_111_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[10] == c_111_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[10] == c_111_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[11] == c_111_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[11] == c_111_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[12] == c_111_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[12] == c_111_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[13] == c_111_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[13] == c_111_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[14] == c_111_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[14] == c_111_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[15] == c_111_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[15] == c_111_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[16] == c_111_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[16] == c_111_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[17] == c_111_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[17] == c_111_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[18] == c_111_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[18] == c_111_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[19] == c_111_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[19] == c_111_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[20] == c_111_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[20] == c_111_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[21] == c_111_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[21] == c_111_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[22] == c_111_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[22] == c_111_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[23] == c_111_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[23] == c_111_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[24] == c_111_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[24] == c_111_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[25] == c_111_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[25] == c_111_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[26] == c_111_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[26] == c_111_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[27] == c_111_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[27] == c_111_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[28] == c_111_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[28] == c_111_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[29] == c_111_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[29] == c_111_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[30] == c_111_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[30] == c_111_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[31] == c_111_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[31] == c_111_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_111[32] == c_111_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_111[32] == c_111_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[0] == c_112_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[0] == c_112_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[1] == c_112_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[1] == c_112_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[2] == c_112_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[2] == c_112_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[3] == c_112_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[3] == c_112_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[4] == c_112_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[4] == c_112_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[5] == c_112_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[5] == c_112_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[6] == c_112_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[6] == c_112_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[7] == c_112_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[7] == c_112_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[8] == c_112_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[8] == c_112_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[9] == c_112_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[9] == c_112_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[10] == c_112_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[10] == c_112_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[11] == c_112_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[11] == c_112_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[12] == c_112_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[12] == c_112_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[13] == c_112_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[13] == c_112_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[14] == c_112_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[14] == c_112_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[15] == c_112_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[15] == c_112_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[16] == c_112_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[16] == c_112_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[17] == c_112_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[17] == c_112_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[18] == c_112_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[18] == c_112_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[19] == c_112_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[19] == c_112_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[20] == c_112_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[20] == c_112_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[21] == c_112_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[21] == c_112_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[22] == c_112_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[22] == c_112_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[23] == c_112_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[23] == c_112_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[24] == c_112_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[24] == c_112_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[25] == c_112_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[25] == c_112_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[26] == c_112_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[26] == c_112_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[27] == c_112_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[27] == c_112_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[28] == c_112_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[28] == c_112_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[29] == c_112_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[29] == c_112_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[30] == c_112_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[30] == c_112_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[31] == c_112_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[31] == c_112_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_112[32] == c_112_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_112[32] == c_112_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[0] == c_113_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[0] == c_113_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[1] == c_113_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[1] == c_113_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[2] == c_113_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[2] == c_113_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[3] == c_113_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[3] == c_113_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[4] == c_113_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[4] == c_113_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[5] == c_113_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[5] == c_113_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[6] == c_113_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[6] == c_113_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[7] == c_113_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[7] == c_113_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[8] == c_113_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[8] == c_113_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[9] == c_113_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[9] == c_113_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[10] == c_113_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[10] == c_113_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[11] == c_113_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[11] == c_113_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[12] == c_113_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[12] == c_113_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[13] == c_113_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[13] == c_113_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[14] == c_113_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[14] == c_113_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[15] == c_113_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[15] == c_113_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[16] == c_113_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[16] == c_113_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[17] == c_113_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[17] == c_113_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[18] == c_113_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[18] == c_113_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[19] == c_113_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[19] == c_113_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[20] == c_113_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[20] == c_113_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[21] == c_113_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[21] == c_113_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[22] == c_113_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[22] == c_113_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[23] == c_113_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[23] == c_113_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[24] == c_113_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[24] == c_113_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[25] == c_113_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[25] == c_113_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[26] == c_113_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[26] == c_113_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[27] == c_113_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[27] == c_113_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[28] == c_113_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[28] == c_113_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[29] == c_113_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[29] == c_113_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[30] == c_113_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[30] == c_113_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[31] == c_113_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[31] == c_113_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_113[32] == c_113_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_113[32] == c_113_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[0] == c_114_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[0] == c_114_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[1] == c_114_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[1] == c_114_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[2] == c_114_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[2] == c_114_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[3] == c_114_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[3] == c_114_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[4] == c_114_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[4] == c_114_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[5] == c_114_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[5] == c_114_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[6] == c_114_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[6] == c_114_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[7] == c_114_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[7] == c_114_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[8] == c_114_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[8] == c_114_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[9] == c_114_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[9] == c_114_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[10] == c_114_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[10] == c_114_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[11] == c_114_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[11] == c_114_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[12] == c_114_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[12] == c_114_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[13] == c_114_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[13] == c_114_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[14] == c_114_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[14] == c_114_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[15] == c_114_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[15] == c_114_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[16] == c_114_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[16] == c_114_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[17] == c_114_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[17] == c_114_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[18] == c_114_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[18] == c_114_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[19] == c_114_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[19] == c_114_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[20] == c_114_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[20] == c_114_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[21] == c_114_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[21] == c_114_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[22] == c_114_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[22] == c_114_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[23] == c_114_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[23] == c_114_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[24] == c_114_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[24] == c_114_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[25] == c_114_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[25] == c_114_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[26] == c_114_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[26] == c_114_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[27] == c_114_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[27] == c_114_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[28] == c_114_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[28] == c_114_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[29] == c_114_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[29] == c_114_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[30] == c_114_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[30] == c_114_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[31] == c_114_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[31] == c_114_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_114[32] == c_114_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_114[32] == c_114_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[0] == c_115_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[0] == c_115_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[1] == c_115_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[1] == c_115_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[2] == c_115_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[2] == c_115_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[3] == c_115_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[3] == c_115_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[4] == c_115_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[4] == c_115_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[5] == c_115_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[5] == c_115_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[6] == c_115_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[6] == c_115_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[7] == c_115_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[7] == c_115_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[8] == c_115_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[8] == c_115_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[9] == c_115_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[9] == c_115_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[10] == c_115_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[10] == c_115_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[11] == c_115_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[11] == c_115_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[12] == c_115_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[12] == c_115_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[13] == c_115_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[13] == c_115_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[14] == c_115_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[14] == c_115_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[15] == c_115_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[15] == c_115_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[16] == c_115_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[16] == c_115_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[17] == c_115_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[17] == c_115_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[18] == c_115_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[18] == c_115_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[19] == c_115_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[19] == c_115_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[20] == c_115_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[20] == c_115_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[21] == c_115_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[21] == c_115_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[22] == c_115_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[22] == c_115_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[23] == c_115_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[23] == c_115_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[24] == c_115_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[24] == c_115_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[25] == c_115_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[25] == c_115_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[26] == c_115_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[26] == c_115_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[27] == c_115_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[27] == c_115_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[28] == c_115_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[28] == c_115_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[29] == c_115_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[29] == c_115_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[30] == c_115_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[30] == c_115_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[31] == c_115_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[31] == c_115_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_115[32] == c_115_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_115[32] == c_115_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[0] == c_116_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[0] == c_116_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[1] == c_116_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[1] == c_116_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[2] == c_116_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[2] == c_116_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[3] == c_116_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[3] == c_116_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[4] == c_116_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[4] == c_116_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[5] == c_116_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[5] == c_116_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[6] == c_116_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[6] == c_116_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[7] == c_116_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[7] == c_116_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[8] == c_116_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[8] == c_116_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[9] == c_116_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[9] == c_116_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[10] == c_116_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[10] == c_116_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[11] == c_116_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[11] == c_116_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[12] == c_116_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[12] == c_116_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[13] == c_116_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[13] == c_116_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[14] == c_116_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[14] == c_116_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[15] == c_116_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[15] == c_116_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[16] == c_116_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[16] == c_116_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[17] == c_116_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[17] == c_116_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[18] == c_116_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[18] == c_116_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[19] == c_116_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[19] == c_116_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[20] == c_116_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[20] == c_116_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[21] == c_116_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[21] == c_116_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[22] == c_116_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[22] == c_116_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[23] == c_116_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[23] == c_116_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[24] == c_116_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[24] == c_116_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[25] == c_116_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[25] == c_116_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[26] == c_116_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[26] == c_116_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[27] == c_116_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[27] == c_116_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[28] == c_116_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[28] == c_116_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[29] == c_116_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[29] == c_116_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[30] == c_116_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[30] == c_116_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[31] == c_116_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[31] == c_116_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_116[32] == c_116_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_116[32] == c_116_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[0] == c_117_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[0] == c_117_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[1] == c_117_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[1] == c_117_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[2] == c_117_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[2] == c_117_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[3] == c_117_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[3] == c_117_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[4] == c_117_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[4] == c_117_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[5] == c_117_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[5] == c_117_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[6] == c_117_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[6] == c_117_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[7] == c_117_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[7] == c_117_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[8] == c_117_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[8] == c_117_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[9] == c_117_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[9] == c_117_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[10] == c_117_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[10] == c_117_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[11] == c_117_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[11] == c_117_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[12] == c_117_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[12] == c_117_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[13] == c_117_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[13] == c_117_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[14] == c_117_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[14] == c_117_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[15] == c_117_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[15] == c_117_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[16] == c_117_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[16] == c_117_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[17] == c_117_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[17] == c_117_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[18] == c_117_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[18] == c_117_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[19] == c_117_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[19] == c_117_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[20] == c_117_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[20] == c_117_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[21] == c_117_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[21] == c_117_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[22] == c_117_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[22] == c_117_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[23] == c_117_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[23] == c_117_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[24] == c_117_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[24] == c_117_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[25] == c_117_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[25] == c_117_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[26] == c_117_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[26] == c_117_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[27] == c_117_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[27] == c_117_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[28] == c_117_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[28] == c_117_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[29] == c_117_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[29] == c_117_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[30] == c_117_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[30] == c_117_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[31] == c_117_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[31] == c_117_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_117[32] == c_117_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_117[32] == c_117_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[0] == c_118_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[0] == c_118_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[1] == c_118_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[1] == c_118_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[2] == c_118_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[2] == c_118_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[3] == c_118_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[3] == c_118_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[4] == c_118_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[4] == c_118_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[5] == c_118_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[5] == c_118_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[6] == c_118_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[6] == c_118_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[7] == c_118_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[7] == c_118_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[8] == c_118_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[8] == c_118_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[9] == c_118_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[9] == c_118_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[10] == c_118_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[10] == c_118_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[11] == c_118_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[11] == c_118_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[12] == c_118_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[12] == c_118_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[13] == c_118_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[13] == c_118_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[14] == c_118_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[14] == c_118_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[15] == c_118_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[15] == c_118_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[16] == c_118_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[16] == c_118_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[17] == c_118_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[17] == c_118_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[18] == c_118_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[18] == c_118_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[19] == c_118_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[19] == c_118_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[20] == c_118_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[20] == c_118_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[21] == c_118_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[21] == c_118_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[22] == c_118_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[22] == c_118_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[23] == c_118_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[23] == c_118_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[24] == c_118_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[24] == c_118_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[25] == c_118_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[25] == c_118_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[26] == c_118_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[26] == c_118_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[27] == c_118_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[27] == c_118_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[28] == c_118_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[28] == c_118_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[29] == c_118_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[29] == c_118_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[30] == c_118_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[30] == c_118_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[31] == c_118_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[31] == c_118_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_118[32] == c_118_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_118[32] == c_118_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[0] == c_119_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[0] == c_119_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[1] == c_119_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[1] == c_119_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[2] == c_119_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[2] == c_119_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[3] == c_119_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[3] == c_119_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[4] == c_119_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[4] == c_119_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[5] == c_119_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[5] == c_119_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[6] == c_119_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[6] == c_119_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[7] == c_119_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[7] == c_119_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[8] == c_119_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[8] == c_119_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[9] == c_119_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[9] == c_119_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[10] == c_119_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[10] == c_119_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[11] == c_119_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[11] == c_119_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[12] == c_119_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[12] == c_119_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[13] == c_119_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[13] == c_119_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[14] == c_119_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[14] == c_119_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[15] == c_119_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[15] == c_119_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[16] == c_119_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[16] == c_119_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[17] == c_119_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[17] == c_119_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[18] == c_119_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[18] == c_119_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[19] == c_119_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[19] == c_119_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[20] == c_119_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[20] == c_119_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[21] == c_119_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[21] == c_119_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[22] == c_119_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[22] == c_119_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[23] == c_119_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[23] == c_119_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[24] == c_119_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[24] == c_119_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[25] == c_119_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[25] == c_119_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[26] == c_119_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[26] == c_119_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[27] == c_119_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[27] == c_119_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[28] == c_119_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[28] == c_119_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[29] == c_119_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[29] == c_119_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[30] == c_119_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[30] == c_119_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[31] == c_119_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[31] == c_119_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_119[32] == c_119_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_119[32] == c_119_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[0] == c_120_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[0] == c_120_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[1] == c_120_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[1] == c_120_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[2] == c_120_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[2] == c_120_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[3] == c_120_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[3] == c_120_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[4] == c_120_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[4] == c_120_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[5] == c_120_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[5] == c_120_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[6] == c_120_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[6] == c_120_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[7] == c_120_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[7] == c_120_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[8] == c_120_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[8] == c_120_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[9] == c_120_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[9] == c_120_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[10] == c_120_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[10] == c_120_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[11] == c_120_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[11] == c_120_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[12] == c_120_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[12] == c_120_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[13] == c_120_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[13] == c_120_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[14] == c_120_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[14] == c_120_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[15] == c_120_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[15] == c_120_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[16] == c_120_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[16] == c_120_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[17] == c_120_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[17] == c_120_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[18] == c_120_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[18] == c_120_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[19] == c_120_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[19] == c_120_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[20] == c_120_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[20] == c_120_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[21] == c_120_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[21] == c_120_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[22] == c_120_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[22] == c_120_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[23] == c_120_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[23] == c_120_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[24] == c_120_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[24] == c_120_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[25] == c_120_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[25] == c_120_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[26] == c_120_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[26] == c_120_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[27] == c_120_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[27] == c_120_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[28] == c_120_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[28] == c_120_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[29] == c_120_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[29] == c_120_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[30] == c_120_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[30] == c_120_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[31] == c_120_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[31] == c_120_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_120[32] == c_120_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_120[32] == c_120_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[0] == c_121_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[0] == c_121_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[1] == c_121_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[1] == c_121_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[2] == c_121_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[2] == c_121_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[3] == c_121_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[3] == c_121_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[4] == c_121_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[4] == c_121_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[5] == c_121_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[5] == c_121_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[6] == c_121_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[6] == c_121_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[7] == c_121_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[7] == c_121_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[8] == c_121_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[8] == c_121_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[9] == c_121_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[9] == c_121_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[10] == c_121_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[10] == c_121_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[11] == c_121_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[11] == c_121_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[12] == c_121_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[12] == c_121_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[13] == c_121_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[13] == c_121_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[14] == c_121_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[14] == c_121_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[15] == c_121_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[15] == c_121_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[16] == c_121_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[16] == c_121_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[17] == c_121_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[17] == c_121_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[18] == c_121_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[18] == c_121_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[19] == c_121_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[19] == c_121_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[20] == c_121_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[20] == c_121_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[21] == c_121_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[21] == c_121_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[22] == c_121_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[22] == c_121_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[23] == c_121_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[23] == c_121_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[24] == c_121_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[24] == c_121_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[25] == c_121_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[25] == c_121_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[26] == c_121_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[26] == c_121_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[27] == c_121_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[27] == c_121_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[28] == c_121_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[28] == c_121_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[29] == c_121_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[29] == c_121_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[30] == c_121_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[30] == c_121_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[31] == c_121_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[31] == c_121_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_121[32] == c_121_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_121[32] == c_121_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[0] == c_122_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[0] == c_122_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[1] == c_122_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[1] == c_122_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[2] == c_122_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[2] == c_122_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[3] == c_122_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[3] == c_122_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[4] == c_122_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[4] == c_122_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[5] == c_122_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[5] == c_122_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[6] == c_122_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[6] == c_122_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[7] == c_122_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[7] == c_122_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[8] == c_122_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[8] == c_122_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[9] == c_122_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[9] == c_122_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[10] == c_122_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[10] == c_122_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[11] == c_122_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[11] == c_122_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[12] == c_122_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[12] == c_122_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[13] == c_122_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[13] == c_122_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[14] == c_122_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[14] == c_122_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[15] == c_122_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[15] == c_122_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[16] == c_122_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[16] == c_122_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[17] == c_122_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[17] == c_122_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[18] == c_122_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[18] == c_122_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[19] == c_122_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[19] == c_122_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[20] == c_122_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[20] == c_122_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[21] == c_122_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[21] == c_122_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[22] == c_122_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[22] == c_122_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[23] == c_122_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[23] == c_122_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[24] == c_122_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[24] == c_122_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[25] == c_122_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[25] == c_122_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[26] == c_122_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[26] == c_122_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[27] == c_122_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[27] == c_122_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[28] == c_122_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[28] == c_122_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[29] == c_122_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[29] == c_122_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[30] == c_122_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[30] == c_122_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[31] == c_122_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[31] == c_122_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_122[32] == c_122_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_122[32] == c_122_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[0] == c_123_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[0] == c_123_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[1] == c_123_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[1] == c_123_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[2] == c_123_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[2] == c_123_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[3] == c_123_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[3] == c_123_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[4] == c_123_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[4] == c_123_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[5] == c_123_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[5] == c_123_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[6] == c_123_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[6] == c_123_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[7] == c_123_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[7] == c_123_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[8] == c_123_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[8] == c_123_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[9] == c_123_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[9] == c_123_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[10] == c_123_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[10] == c_123_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[11] == c_123_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[11] == c_123_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[12] == c_123_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[12] == c_123_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[13] == c_123_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[13] == c_123_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[14] == c_123_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[14] == c_123_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[15] == c_123_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[15] == c_123_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[16] == c_123_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[16] == c_123_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[17] == c_123_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[17] == c_123_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[18] == c_123_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[18] == c_123_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[19] == c_123_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[19] == c_123_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[20] == c_123_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[20] == c_123_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[21] == c_123_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[21] == c_123_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[22] == c_123_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[22] == c_123_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[23] == c_123_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[23] == c_123_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[24] == c_123_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[24] == c_123_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[25] == c_123_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[25] == c_123_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[26] == c_123_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[26] == c_123_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[27] == c_123_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[27] == c_123_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[28] == c_123_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[28] == c_123_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[29] == c_123_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[29] == c_123_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[30] == c_123_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[30] == c_123_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[31] == c_123_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[31] == c_123_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_123[32] == c_123_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_123[32] == c_123_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[0] == c_124_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[0] == c_124_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[1] == c_124_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[1] == c_124_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[2] == c_124_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[2] == c_124_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[3] == c_124_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[3] == c_124_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[4] == c_124_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[4] == c_124_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[5] == c_124_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[5] == c_124_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[6] == c_124_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[6] == c_124_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[7] == c_124_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[7] == c_124_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[8] == c_124_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[8] == c_124_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[9] == c_124_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[9] == c_124_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[10] == c_124_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[10] == c_124_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[11] == c_124_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[11] == c_124_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[12] == c_124_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[12] == c_124_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[13] == c_124_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[13] == c_124_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[14] == c_124_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[14] == c_124_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[15] == c_124_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[15] == c_124_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[16] == c_124_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[16] == c_124_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[17] == c_124_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[17] == c_124_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[18] == c_124_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[18] == c_124_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[19] == c_124_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[19] == c_124_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[20] == c_124_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[20] == c_124_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[21] == c_124_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[21] == c_124_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[22] == c_124_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[22] == c_124_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[23] == c_124_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[23] == c_124_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[24] == c_124_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[24] == c_124_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[25] == c_124_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[25] == c_124_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[26] == c_124_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[26] == c_124_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[27] == c_124_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[27] == c_124_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[28] == c_124_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[28] == c_124_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[29] == c_124_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[29] == c_124_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[30] == c_124_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[30] == c_124_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[31] == c_124_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[31] == c_124_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_124[32] == c_124_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_124[32] == c_124_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[0] == c_125_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[0] == c_125_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[1] == c_125_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[1] == c_125_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[2] == c_125_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[2] == c_125_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[3] == c_125_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[3] == c_125_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[4] == c_125_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[4] == c_125_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[5] == c_125_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[5] == c_125_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[6] == c_125_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[6] == c_125_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[7] == c_125_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[7] == c_125_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[8] == c_125_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[8] == c_125_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[9] == c_125_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[9] == c_125_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[10] == c_125_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[10] == c_125_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[11] == c_125_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[11] == c_125_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[12] == c_125_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[12] == c_125_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[13] == c_125_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[13] == c_125_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[14] == c_125_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[14] == c_125_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[15] == c_125_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[15] == c_125_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[16] == c_125_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[16] == c_125_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[17] == c_125_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[17] == c_125_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[18] == c_125_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[18] == c_125_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[19] == c_125_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[19] == c_125_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[20] == c_125_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[20] == c_125_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[21] == c_125_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[21] == c_125_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[22] == c_125_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[22] == c_125_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[23] == c_125_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[23] == c_125_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[24] == c_125_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[24] == c_125_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[25] == c_125_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[25] == c_125_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[26] == c_125_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[26] == c_125_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[27] == c_125_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[27] == c_125_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[28] == c_125_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[28] == c_125_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[29] == c_125_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[29] == c_125_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[30] == c_125_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[30] == c_125_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[31] == c_125_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[31] == c_125_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_125[32] == c_125_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_125[32] == c_125_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[0] == c_126_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[0] == c_126_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[1] == c_126_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[1] == c_126_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[2] == c_126_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[2] == c_126_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[3] == c_126_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[3] == c_126_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[4] == c_126_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[4] == c_126_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[5] == c_126_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[5] == c_126_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[6] == c_126_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[6] == c_126_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[7] == c_126_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[7] == c_126_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[8] == c_126_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[8] == c_126_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[9] == c_126_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[9] == c_126_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[10] == c_126_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[10] == c_126_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[11] == c_126_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[11] == c_126_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[12] == c_126_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[12] == c_126_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[13] == c_126_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[13] == c_126_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[14] == c_126_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[14] == c_126_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[15] == c_126_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[15] == c_126_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[16] == c_126_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[16] == c_126_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[17] == c_126_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[17] == c_126_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[18] == c_126_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[18] == c_126_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[19] == c_126_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[19] == c_126_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[20] == c_126_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[20] == c_126_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[21] == c_126_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[21] == c_126_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[22] == c_126_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[22] == c_126_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[23] == c_126_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[23] == c_126_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[24] == c_126_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[24] == c_126_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[25] == c_126_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[25] == c_126_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[26] == c_126_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[26] == c_126_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[27] == c_126_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[27] == c_126_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[28] == c_126_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[28] == c_126_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[29] == c_126_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[29] == c_126_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[30] == c_126_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[30] == c_126_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[31] == c_126_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[31] == c_126_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_126[32] == c_126_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_126[32] == c_126_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[0] == c_127_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[0] == c_127_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[1] == c_127_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[1] == c_127_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[2] == c_127_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[2] == c_127_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[3] == c_127_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[3] == c_127_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[4] == c_127_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[4] == c_127_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[5] == c_127_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[5] == c_127_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[6] == c_127_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[6] == c_127_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[7] == c_127_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[7] == c_127_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[8] == c_127_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[8] == c_127_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[9] == c_127_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[9] == c_127_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[10] == c_127_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[10] == c_127_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[11] == c_127_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[11] == c_127_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[12] == c_127_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[12] == c_127_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[13] == c_127_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[13] == c_127_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[14] == c_127_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[14] == c_127_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[15] == c_127_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[15] == c_127_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[16] == c_127_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[16] == c_127_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[17] == c_127_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[17] == c_127_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[18] == c_127_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[18] == c_127_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[19] == c_127_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[19] == c_127_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[20] == c_127_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[20] == c_127_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[21] == c_127_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[21] == c_127_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[22] == c_127_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[22] == c_127_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[23] == c_127_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[23] == c_127_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[24] == c_127_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[24] == c_127_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[25] == c_127_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[25] == c_127_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[26] == c_127_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[26] == c_127_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[27] == c_127_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[27] == c_127_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[28] == c_127_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[28] == c_127_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[29] == c_127_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[29] == c_127_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[30] == c_127_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[30] == c_127_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[31] == c_127_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[31] == c_127_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_127[32] == c_127_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_127[32] == c_127_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[0] == c_128_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[0] == c_128_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[1] == c_128_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[1] == c_128_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[2] == c_128_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[2] == c_128_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[3] == c_128_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[3] == c_128_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[4] == c_128_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[4] == c_128_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[5] == c_128_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[5] == c_128_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[6] == c_128_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[6] == c_128_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[7] == c_128_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[7] == c_128_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[8] == c_128_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[8] == c_128_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[9] == c_128_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[9] == c_128_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[10] == c_128_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[10] == c_128_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[11] == c_128_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[11] == c_128_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[12] == c_128_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[12] == c_128_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[13] == c_128_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[13] == c_128_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[14] == c_128_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[14] == c_128_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[15] == c_128_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[15] == c_128_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[16] == c_128_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[16] == c_128_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[17] == c_128_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[17] == c_128_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[18] == c_128_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[18] == c_128_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[19] == c_128_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[19] == c_128_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[20] == c_128_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[20] == c_128_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[21] == c_128_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[21] == c_128_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[22] == c_128_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[22] == c_128_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[23] == c_128_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[23] == c_128_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[24] == c_128_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[24] == c_128_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[25] == c_128_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[25] == c_128_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[26] == c_128_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[26] == c_128_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[27] == c_128_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[27] == c_128_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[28] == c_128_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[28] == c_128_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[29] == c_128_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[29] == c_128_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[30] == c_128_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[30] == c_128_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[31] == c_128_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[31] == c_128_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_128[32] == c_128_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_128[32] == c_128_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[0] == c_129_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[0] == c_129_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[1] == c_129_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[1] == c_129_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[2] == c_129_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[2] == c_129_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[3] == c_129_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[3] == c_129_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[4] == c_129_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[4] == c_129_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[5] == c_129_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[5] == c_129_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[6] == c_129_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[6] == c_129_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[7] == c_129_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[7] == c_129_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[8] == c_129_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[8] == c_129_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[9] == c_129_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[9] == c_129_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[10] == c_129_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[10] == c_129_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[11] == c_129_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[11] == c_129_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[12] == c_129_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[12] == c_129_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[13] == c_129_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[13] == c_129_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[14] == c_129_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[14] == c_129_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[15] == c_129_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[15] == c_129_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[16] == c_129_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[16] == c_129_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[17] == c_129_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[17] == c_129_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[18] == c_129_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[18] == c_129_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[19] == c_129_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[19] == c_129_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[20] == c_129_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[20] == c_129_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[21] == c_129_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[21] == c_129_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[22] == c_129_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[22] == c_129_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[23] == c_129_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[23] == c_129_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[24] == c_129_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[24] == c_129_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[25] == c_129_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[25] == c_129_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[26] == c_129_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[26] == c_129_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[27] == c_129_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[27] == c_129_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[28] == c_129_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[28] == c_129_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[29] == c_129_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[29] == c_129_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[30] == c_129_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[30] == c_129_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[31] == c_129_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[31] == c_129_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_129[32] == c_129_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_129[32] == c_129_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[0] == c_130_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[0] == c_130_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[1] == c_130_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[1] == c_130_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[2] == c_130_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[2] == c_130_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[3] == c_130_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[3] == c_130_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[4] == c_130_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[4] == c_130_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[5] == c_130_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[5] == c_130_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[6] == c_130_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[6] == c_130_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[7] == c_130_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[7] == c_130_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[8] == c_130_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[8] == c_130_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[9] == c_130_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[9] == c_130_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[10] == c_130_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[10] == c_130_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[11] == c_130_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[11] == c_130_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[12] == c_130_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[12] == c_130_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[13] == c_130_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[13] == c_130_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[14] == c_130_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[14] == c_130_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[15] == c_130_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[15] == c_130_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[16] == c_130_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[16] == c_130_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[17] == c_130_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[17] == c_130_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[18] == c_130_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[18] == c_130_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[19] == c_130_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[19] == c_130_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[20] == c_130_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[20] == c_130_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[21] == c_130_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[21] == c_130_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[22] == c_130_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[22] == c_130_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[23] == c_130_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[23] == c_130_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[24] == c_130_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[24] == c_130_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[25] == c_130_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[25] == c_130_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[26] == c_130_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[26] == c_130_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[27] == c_130_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[27] == c_130_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[28] == c_130_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[28] == c_130_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[29] == c_130_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[29] == c_130_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[30] == c_130_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[30] == c_130_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[31] == c_130_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[31] == c_130_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_130[32] == c_130_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_130[32] == c_130_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[0] == c_131_0)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[0] == c_131_0)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[1] == c_131_1)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[1] == c_131_1)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[2] == c_131_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[2] == c_131_2)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[3] == c_131_3)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[3] == c_131_3)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[4] == c_131_4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[4] == c_131_4)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[5] == c_131_5)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[5] == c_131_5)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[6] == c_131_6)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[6] == c_131_6)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[7] == c_131_7)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[7] == c_131_7)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[8] == c_131_8)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[8] == c_131_8)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[9] == c_131_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[9] == c_131_9)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[10] == c_131_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[10] == c_131_10)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[11] == c_131_11)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[11] == c_131_11)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[12] == c_131_12)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[12] == c_131_12)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[13] == c_131_13)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[13] == c_131_13)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[14] == c_131_14)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[14] == c_131_14)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[15] == c_131_15)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[15] == c_131_15)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[16] == c_131_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[16] == c_131_16)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[17] == c_131_17)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[17] == c_131_17)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[18] == c_131_18)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[18] == c_131_18)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[19] == c_131_19)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[19] == c_131_19)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[20] == c_131_20)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[20] == c_131_20)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[21] == c_131_21)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[21] == c_131_21)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[22] == c_131_22)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[22] == c_131_22)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[23] == c_131_23)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[23] == c_131_23)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[24] == c_131_24)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[24] == c_131_24)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[25] == c_131_25)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[25] == c_131_25)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[26] == c_131_26)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[26] == c_131_26)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[27] == c_131_27)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[27] == c_131_27)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[28] == c_131_28)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[28] == c_131_28)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[29] == c_131_29)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[29] == c_131_29)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[30] == c_131_30)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[30] == c_131_30)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[31] == c_131_31)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[31] == c_131_31)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_out_131[32] == c_131_32)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at WallaceTest.scala:112 chisel3.assert(io.out(j)(i) === io.in(i)(j))\n"); // @[WallaceTest.scala 112:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_out_131[32] == c_131_32)) begin
          $fatal; // @[WallaceTest.scala 112:21]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSA(
  input  [2:0] io_in,
  output [1:0] io_out
);
  wire  _out_1_T_6 = io_in[0] ^ io_in[1]; // @[WallaceTest.scala 27:59]
  wire  out_1 = io_in[0] & io_in[1] | io_in[2] & (io_in[0] ^ io_in[1]); // @[WallaceTest.scala 27:35]
  wire  out_0 = _out_1_T_6 ^ io_in[2]; // @[WallaceTest.scala 28:33]
  assign io_out = {out_1,out_0}; // @[Cat.scala 33:92]
endmodule
module Walloc33bits(
  input  [32:0] io_src_in,
  input  [29:0] io_cin,
  output        io_cout_group_0,
  output        io_cout_group_1,
  output        io_cout_group_2,
  output        io_cout_group_3,
  output        io_cout_group_4,
  output        io_cout_group_5,
  output        io_cout_group_6,
  output        io_cout_group_7,
  output        io_cout_group_8,
  output        io_cout_group_9,
  output        io_cout_group_10,
  output        io_cout_group_11,
  output        io_cout_group_12,
  output        io_cout_group_13,
  output        io_cout_group_14,
  output        io_cout_group_15,
  output        io_cout_group_16,
  output        io_cout_group_17,
  output        io_cout_group_18,
  output        io_cout_group_19,
  output        io_cout_group_20,
  output        io_cout_group_21,
  output        io_cout_group_22,
  output        io_cout_group_23,
  output        io_cout_group_24,
  output        io_cout_group_25,
  output        io_cout_group_26,
  output        io_cout_group_27,
  output        io_cout_group_28,
  output        io_cout_group_29,
  output        io_cout,
  output        io_s
);
  wire [2:0] csa_0_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_0_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_1_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_1_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_2_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_2_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_3_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_3_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_4_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_4_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_5_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_5_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_6_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_6_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_7_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_7_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_8_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_8_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_9_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_9_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_10_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_10_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_11_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_11_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_12_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_12_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_13_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_13_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_14_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_14_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_15_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_15_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_16_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_16_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_17_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_17_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_18_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_18_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_19_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_19_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_20_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_20_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_21_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_21_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_22_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_22_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_23_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_23_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_24_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_24_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_25_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_25_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_26_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_26_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_27_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_27_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_28_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_28_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_29_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_29_io_out; // @[WallaceTest.scala 128:33]
  wire [2:0] csa_30_io_in; // @[WallaceTest.scala 128:33]
  wire [1:0] csa_30_io_out; // @[WallaceTest.scala 128:33]
  wire  first_s_10 = csa_0_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_9 = csa_1_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_8 = csa_2_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_7 = csa_3_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_6 = csa_4_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_5 = csa_5_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_4 = csa_6_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_3 = csa_7_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_2 = csa_8_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_1 = csa_9_io_out[0]; // @[WallaceTest.scala 135:36]
  wire  first_s_0 = csa_10_io_out[0]; // @[WallaceTest.scala 135:36]
  wire [4:0] csa_11_io_in_lo = {first_s_4,first_s_3,first_s_2,first_s_1,first_s_0}; // @[WallaceTest.scala 140:30]
  wire [10:0] _csa_11_io_in_T = {first_s_10,first_s_9,first_s_8,first_s_7,first_s_6,first_s_5,csa_11_io_in_lo}; // @[WallaceTest.scala 140:30]
  wire  second_s_8 = csa_11_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_7 = csa_12_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_6 = csa_13_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_5 = csa_14_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_4 = csa_15_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_3 = csa_16_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_2 = csa_17_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_1 = csa_18_io_out[0]; // @[WallaceTest.scala 152:40]
  wire  second_s_0 = csa_19_io_out[0]; // @[WallaceTest.scala 152:40]
  wire [8:0] _csa_20_io_in_T = {second_s_8,second_s_7,second_s_6,second_s_5,second_s_4,second_s_3,second_s_2,second_s_1,
    second_s_0}; // @[WallaceTest.scala 159:30]
  wire  third_s_6 = csa_20_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_5 = csa_21_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_4 = csa_22_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_3 = csa_23_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_2 = csa_24_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_1 = csa_25_io_out[0]; // @[WallaceTest.scala 169:39]
  wire  third_s_0 = csa_26_io_out[0]; // @[WallaceTest.scala 169:39]
  wire [6:0] _csa_27_io_in_T = {third_s_6,third_s_5,third_s_4,third_s_3,third_s_2,third_s_1,third_s_0}; // @[WallaceTest.scala 176:28]
  wire  fourth_s_2 = csa_27_io_out[0]; // @[WallaceTest.scala 182:40]
  wire  fourth_s_1 = csa_28_io_out[0]; // @[WallaceTest.scala 182:40]
  wire  fourth_s_0 = csa_29_io_out[0]; // @[WallaceTest.scala 182:40]
  wire [1:0] csa_30_io_in_hi = {fourth_s_2,fourth_s_1}; // @[WallaceTest.scala 186:29]
  CSA csa_0 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_0_io_in),
    .io_out(csa_0_io_out)
  );
  CSA csa_1 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_1_io_in),
    .io_out(csa_1_io_out)
  );
  CSA csa_2 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_2_io_in),
    .io_out(csa_2_io_out)
  );
  CSA csa_3 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_3_io_in),
    .io_out(csa_3_io_out)
  );
  CSA csa_4 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_4_io_in),
    .io_out(csa_4_io_out)
  );
  CSA csa_5 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_5_io_in),
    .io_out(csa_5_io_out)
  );
  CSA csa_6 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_6_io_in),
    .io_out(csa_6_io_out)
  );
  CSA csa_7 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_7_io_in),
    .io_out(csa_7_io_out)
  );
  CSA csa_8 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_8_io_in),
    .io_out(csa_8_io_out)
  );
  CSA csa_9 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_9_io_in),
    .io_out(csa_9_io_out)
  );
  CSA csa_10 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_10_io_in),
    .io_out(csa_10_io_out)
  );
  CSA csa_11 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_11_io_in),
    .io_out(csa_11_io_out)
  );
  CSA csa_12 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_12_io_in),
    .io_out(csa_12_io_out)
  );
  CSA csa_13 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_13_io_in),
    .io_out(csa_13_io_out)
  );
  CSA csa_14 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_14_io_in),
    .io_out(csa_14_io_out)
  );
  CSA csa_15 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_15_io_in),
    .io_out(csa_15_io_out)
  );
  CSA csa_16 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_16_io_in),
    .io_out(csa_16_io_out)
  );
  CSA csa_17 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_17_io_in),
    .io_out(csa_17_io_out)
  );
  CSA csa_18 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_18_io_in),
    .io_out(csa_18_io_out)
  );
  CSA csa_19 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_19_io_in),
    .io_out(csa_19_io_out)
  );
  CSA csa_20 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_20_io_in),
    .io_out(csa_20_io_out)
  );
  CSA csa_21 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_21_io_in),
    .io_out(csa_21_io_out)
  );
  CSA csa_22 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_22_io_in),
    .io_out(csa_22_io_out)
  );
  CSA csa_23 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_23_io_in),
    .io_out(csa_23_io_out)
  );
  CSA csa_24 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_24_io_in),
    .io_out(csa_24_io_out)
  );
  CSA csa_25 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_25_io_in),
    .io_out(csa_25_io_out)
  );
  CSA csa_26 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_26_io_in),
    .io_out(csa_26_io_out)
  );
  CSA csa_27 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_27_io_in),
    .io_out(csa_27_io_out)
  );
  CSA csa_28 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_28_io_in),
    .io_out(csa_28_io_out)
  );
  CSA csa_29 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_29_io_in),
    .io_out(csa_29_io_out)
  );
  CSA csa_30 ( // @[WallaceTest.scala 128:33]
    .io_in(csa_30_io_in),
    .io_out(csa_30_io_out)
  );
  assign io_cout_group_0 = csa_10_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_1 = csa_9_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_2 = csa_8_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_3 = csa_7_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_4 = csa_6_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_5 = csa_5_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_6 = csa_4_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_7 = csa_3_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_8 = csa_2_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_9 = csa_1_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_10 = csa_0_io_out[1]; // @[WallaceTest.scala 134:28]
  assign io_cout_group_11 = csa_19_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_12 = csa_18_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_13 = csa_17_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_14 = csa_16_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_15 = csa_15_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_16 = csa_14_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_17 = csa_13_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_18 = csa_12_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_19 = csa_11_io_out[1]; // @[WallaceTest.scala 151:32]
  assign io_cout_group_20 = csa_26_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_21 = csa_25_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_22 = csa_24_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_23 = csa_23_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_24 = csa_22_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_25 = csa_21_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_26 = csa_20_io_out[1]; // @[WallaceTest.scala 168:32]
  assign io_cout_group_27 = csa_29_io_out[1]; // @[WallaceTest.scala 181:32]
  assign io_cout_group_28 = csa_28_io_out[1]; // @[WallaceTest.scala 181:32]
  assign io_cout_group_29 = csa_27_io_out[1]; // @[WallaceTest.scala 181:32]
  assign io_cout = csa_30_io_out[1]; // @[WallaceTest.scala 187:26]
  assign io_s = csa_30_io_out[0]; // @[WallaceTest.scala 188:25]
  assign csa_0_io_in = io_src_in[32:30]; // @[WallaceTest.scala 133:30]
  assign csa_1_io_in = io_src_in[29:27]; // @[WallaceTest.scala 133:30]
  assign csa_2_io_in = io_src_in[26:24]; // @[WallaceTest.scala 133:30]
  assign csa_3_io_in = io_src_in[23:21]; // @[WallaceTest.scala 133:30]
  assign csa_4_io_in = io_src_in[20:18]; // @[WallaceTest.scala 133:30]
  assign csa_5_io_in = io_src_in[17:15]; // @[WallaceTest.scala 133:30]
  assign csa_6_io_in = io_src_in[14:12]; // @[WallaceTest.scala 133:30]
  assign csa_7_io_in = io_src_in[11:9]; // @[WallaceTest.scala 133:30]
  assign csa_8_io_in = io_src_in[8:6]; // @[WallaceTest.scala 133:30]
  assign csa_9_io_in = io_src_in[5:3]; // @[WallaceTest.scala 133:30]
  assign csa_10_io_in = io_src_in[2:0]; // @[WallaceTest.scala 133:30]
  assign csa_11_io_in = _csa_11_io_in_T[10:8]; // @[WallaceTest.scala 140:36]
  assign csa_12_io_in = _csa_11_io_in_T[7:5]; // @[WallaceTest.scala 141:36]
  assign csa_13_io_in = _csa_11_io_in_T[4:2]; // @[WallaceTest.scala 142:36]
  assign csa_14_io_in = {_csa_11_io_in_T[1:0],io_cin[15]}; // @[Cat.scala 33:92]
  assign csa_15_io_in = io_cin[14:12]; // @[WallaceTest.scala 144:25]
  assign csa_16_io_in = io_cin[11:9]; // @[WallaceTest.scala 145:25]
  assign csa_17_io_in = io_cin[8:6]; // @[WallaceTest.scala 146:25]
  assign csa_18_io_in = io_cin[5:3]; // @[WallaceTest.scala 147:25]
  assign csa_19_io_in = io_cin[2:0]; // @[WallaceTest.scala 148:25]
  assign csa_20_io_in = _csa_20_io_in_T[8:6]; // @[WallaceTest.scala 159:36]
  assign csa_21_io_in = _csa_20_io_in_T[5:3]; // @[WallaceTest.scala 160:36]
  assign csa_22_io_in = _csa_20_io_in_T[2:0]; // @[WallaceTest.scala 161:36]
  assign csa_23_io_in = io_cin[27:25]; // @[WallaceTest.scala 162:24]
  assign csa_24_io_in = io_cin[24:22]; // @[WallaceTest.scala 163:24]
  assign csa_25_io_in = io_cin[21:19]; // @[WallaceTest.scala 164:24]
  assign csa_26_io_in = io_cin[18:16]; // @[WallaceTest.scala 165:24]
  assign csa_27_io_in = _csa_27_io_in_T[6:4]; // @[WallaceTest.scala 176:34]
  assign csa_28_io_in = _csa_27_io_in_T[3:1]; // @[WallaceTest.scala 177:34]
  assign csa_29_io_in = {_csa_27_io_in_T[0],io_cin[29:28]}; // @[Cat.scala 33:92]
  assign csa_30_io_in = {csa_30_io_in_hi,fourth_s_0}; // @[WallaceTest.scala 186:29]
endmodule
module walloc_64_mul(
  input          clock,
  input          reset,
  input  [131:0] io_multiplicand,
  input  [65:0]  io_multiplier,
  output [63:0]  io_result_hi,
  output [63:0]  io_result_lo
);
  wire [2:0] gen_p_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_1_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_1_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_1_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_1_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_2_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_2_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_2_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_2_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_3_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_3_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_3_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_3_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_4_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_4_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_4_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_4_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_5_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_5_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_5_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_5_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_6_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_6_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_6_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_6_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_7_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_7_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_7_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_7_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_8_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_8_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_8_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_8_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_9_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_9_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_9_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_9_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_10_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_10_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_10_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_10_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_11_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_11_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_11_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_11_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_12_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_12_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_12_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_12_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_13_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_13_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_13_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_13_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_14_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_14_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_14_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_14_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_15_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_15_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_15_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_15_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_16_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_16_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_16_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_16_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_17_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_17_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_17_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_17_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_18_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_18_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_18_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_18_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_19_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_19_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_19_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_19_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_20_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_20_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_20_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_20_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_21_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_21_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_21_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_21_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_22_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_22_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_22_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_22_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_23_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_23_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_23_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_23_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_24_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_24_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_24_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_24_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_25_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_25_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_25_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_25_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_26_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_26_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_26_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_26_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_27_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_27_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_27_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_27_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_28_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_28_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_28_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_28_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_29_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_29_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_29_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_29_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_30_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_30_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_30_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_30_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_31_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_31_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_31_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_31_io_c; // @[WallaceTest.scala 204:30]
  wire [2:0] gen_p_32_io_src; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_32_io_x; // @[WallaceTest.scala 204:30]
  wire [131:0] gen_p_32_io_p; // @[WallaceTest.scala 204:30]
  wire  gen_p_32_io_c; // @[WallaceTest.scala 204:30]
  wire  switch_clock; // @[WallaceTest.scala 205:16]
  wire  switch_reset; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_0; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_1; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_2; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_3; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_4; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_5; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_6; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_7; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_8; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_9; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_10; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_11; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_12; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_13; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_14; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_15; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_16; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_17; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_18; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_19; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_20; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_21; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_22; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_23; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_24; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_25; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_26; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_27; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_28; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_29; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_30; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_31; // @[WallaceTest.scala 205:16]
  wire [131:0] switch_io_in_32; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_0; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_1; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_2; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_3; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_4; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_5; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_6; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_7; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_8; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_9; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_10; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_11; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_12; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_13; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_14; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_15; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_16; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_17; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_18; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_19; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_20; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_21; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_22; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_23; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_24; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_25; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_26; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_27; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_28; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_29; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_30; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_31; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_32; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_33; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_34; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_35; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_36; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_37; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_38; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_39; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_40; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_41; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_42; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_43; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_44; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_45; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_46; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_47; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_48; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_49; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_50; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_51; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_52; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_53; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_54; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_55; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_56; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_57; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_58; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_59; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_60; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_61; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_62; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_63; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_64; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_65; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_66; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_67; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_68; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_69; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_70; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_71; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_72; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_73; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_74; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_75; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_76; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_77; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_78; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_79; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_80; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_81; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_82; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_83; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_84; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_85; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_86; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_87; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_88; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_89; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_90; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_91; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_92; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_93; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_94; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_95; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_96; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_97; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_98; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_99; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_100; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_101; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_102; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_103; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_104; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_105; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_106; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_107; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_108; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_109; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_110; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_111; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_112; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_113; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_114; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_115; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_116; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_117; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_118; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_119; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_120; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_121; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_122; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_123; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_124; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_125; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_126; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_127; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_128; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_129; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_130; // @[WallaceTest.scala 205:16]
  wire [32:0] switch_io_out_131; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_0; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_1; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_2; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_3; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_4; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_5; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_6; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_7; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_8; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_9; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_10; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_11; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_12; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_13; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_14; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_15; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_16; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_17; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_18; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_19; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_20; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_21; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_22; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_23; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_24; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_25; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_26; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_27; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_28; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_29; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_30; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_31; // @[WallaceTest.scala 205:16]
  wire  switch_io_cin_32; // @[WallaceTest.scala 205:16]
  wire [31:0] switch_io_cout; // @[WallaceTest.scala 205:16]
  wire [32:0] Walloc33bits_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_1_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_1_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_1_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_2_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_2_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_2_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_3_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_3_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_3_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_4_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_4_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_4_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_5_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_5_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_5_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_6_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_6_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_6_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_7_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_7_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_7_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_8_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_8_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_8_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_9_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_9_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_9_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_10_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_10_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_10_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_11_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_11_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_11_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_12_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_12_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_12_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_13_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_13_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_13_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_14_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_14_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_14_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_15_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_15_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_15_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_16_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_16_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_16_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_17_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_17_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_17_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_18_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_18_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_18_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_19_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_19_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_19_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_20_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_20_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_20_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_21_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_21_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_21_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_22_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_22_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_22_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_23_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_23_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_23_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_24_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_24_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_24_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_25_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_25_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_25_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_26_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_26_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_26_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_27_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_27_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_27_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_28_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_28_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_28_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_29_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_29_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_29_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_30_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_30_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_30_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_31_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_31_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_31_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_32_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_32_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_32_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_33_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_33_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_33_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_34_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_34_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_34_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_35_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_35_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_35_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_36_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_36_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_36_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_37_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_37_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_37_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_38_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_38_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_38_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_39_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_39_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_39_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_40_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_40_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_40_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_41_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_41_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_41_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_42_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_42_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_42_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_43_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_43_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_43_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_44_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_44_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_44_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_45_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_45_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_45_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_46_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_46_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_46_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_47_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_47_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_47_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_48_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_48_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_48_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_49_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_49_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_49_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_50_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_50_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_50_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_51_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_51_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_51_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_52_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_52_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_52_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_53_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_53_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_53_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_54_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_54_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_54_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_55_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_55_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_55_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_56_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_56_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_56_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_57_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_57_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_57_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_58_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_58_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_58_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_59_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_59_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_59_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_60_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_60_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_60_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_61_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_61_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_61_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_62_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_62_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_62_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_63_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_63_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_63_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_64_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_64_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_64_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_65_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_65_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_65_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_66_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_66_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_66_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_67_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_67_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_67_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_68_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_68_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_68_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_69_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_69_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_69_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_70_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_70_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_70_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_71_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_71_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_71_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_72_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_72_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_72_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_73_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_73_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_73_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_74_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_74_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_74_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_75_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_75_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_75_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_76_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_76_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_76_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_77_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_77_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_77_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_78_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_78_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_78_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_79_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_79_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_79_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_80_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_80_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_80_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_81_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_81_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_81_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_82_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_82_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_82_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_83_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_83_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_83_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_84_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_84_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_84_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_85_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_85_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_85_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_86_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_86_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_86_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_87_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_87_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_87_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_88_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_88_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_88_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_89_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_89_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_89_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_90_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_90_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_90_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_91_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_91_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_91_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_92_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_92_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_92_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_93_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_93_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_93_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_94_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_94_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_94_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_95_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_95_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_95_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_96_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_96_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_96_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_97_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_97_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_97_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_98_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_98_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_98_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_99_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_99_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_99_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_100_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_100_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_100_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_101_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_101_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_101_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_102_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_102_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_102_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_103_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_103_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_103_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_104_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_104_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_104_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_105_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_105_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_105_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_106_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_106_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_106_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_107_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_107_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_107_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_108_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_108_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_108_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_109_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_109_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_109_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_110_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_110_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_110_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_111_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_111_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_111_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_112_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_112_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_112_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_113_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_113_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_113_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_114_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_114_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_114_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_115_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_115_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_115_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_116_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_116_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_116_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_117_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_117_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_117_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_118_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_118_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_118_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_119_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_119_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_119_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_120_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_120_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_120_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_121_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_121_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_121_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_122_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_122_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_122_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_123_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_123_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_123_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_124_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_124_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_124_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_125_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_125_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_125_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_126_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_126_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_126_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_127_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_127_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_127_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_128_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_128_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_128_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_129_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_129_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_129_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_130_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_130_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_130_io_s; // @[WallaceTest.scala 206:30]
  wire [32:0] Walloc33bits_131_io_src_in; // @[WallaceTest.scala 206:30]
  wire [29:0] Walloc33bits_131_io_cin; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_0; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_1; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_2; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_3; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_4; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_5; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_6; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_7; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_8; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_9; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_10; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_11; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_12; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_13; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_14; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_15; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_16; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_17; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_18; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_19; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_20; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_21; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_22; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_23; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_24; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_25; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_26; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_27; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_28; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout_group_29; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_cout; // @[WallaceTest.scala 206:30]
  wire  Walloc33bits_131_io_s; // @[WallaceTest.scala 206:30]
  wire [66:0] mulb = {io_multiplier,1'h0}; // @[Cat.scala 33:92]
  wire [6:0] lo_lo = {Walloc33bits_io_cout_group_6,Walloc33bits_io_cout_group_5,Walloc33bits_io_cout_group_4,
    Walloc33bits_io_cout_group_3,Walloc33bits_io_cout_group_2,Walloc33bits_io_cout_group_1,Walloc33bits_io_cout_group_0}
    ; // @[WallaceTest.scala 224:37]
  wire [14:0] lo = {Walloc33bits_io_cout_group_14,Walloc33bits_io_cout_group_13,Walloc33bits_io_cout_group_12,
    Walloc33bits_io_cout_group_11,Walloc33bits_io_cout_group_10,Walloc33bits_io_cout_group_9,
    Walloc33bits_io_cout_group_8,Walloc33bits_io_cout_group_7,lo_lo}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo = {Walloc33bits_io_cout_group_21,Walloc33bits_io_cout_group_20,Walloc33bits_io_cout_group_19,
    Walloc33bits_io_cout_group_18,Walloc33bits_io_cout_group_17,Walloc33bits_io_cout_group_16,
    Walloc33bits_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi = {Walloc33bits_io_cout_group_29,Walloc33bits_io_cout_group_28,Walloc33bits_io_cout_group_27,
    Walloc33bits_io_cout_group_26,Walloc33bits_io_cout_group_25,Walloc33bits_io_cout_group_24,
    Walloc33bits_io_cout_group_23,Walloc33bits_io_cout_group_22,hi_lo}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_1 = {Walloc33bits_1_io_cout_group_6,Walloc33bits_1_io_cout_group_5,Walloc33bits_1_io_cout_group_4,
    Walloc33bits_1_io_cout_group_3,Walloc33bits_1_io_cout_group_2,Walloc33bits_1_io_cout_group_1,
    Walloc33bits_1_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_1 = {Walloc33bits_1_io_cout_group_14,Walloc33bits_1_io_cout_group_13,Walloc33bits_1_io_cout_group_12,
    Walloc33bits_1_io_cout_group_11,Walloc33bits_1_io_cout_group_10,Walloc33bits_1_io_cout_group_9,
    Walloc33bits_1_io_cout_group_8,Walloc33bits_1_io_cout_group_7,lo_lo_1}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_1 = {Walloc33bits_1_io_cout_group_21,Walloc33bits_1_io_cout_group_20,Walloc33bits_1_io_cout_group_19,
    Walloc33bits_1_io_cout_group_18,Walloc33bits_1_io_cout_group_17,Walloc33bits_1_io_cout_group_16,
    Walloc33bits_1_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_1 = {Walloc33bits_1_io_cout_group_29,Walloc33bits_1_io_cout_group_28,Walloc33bits_1_io_cout_group_27,
    Walloc33bits_1_io_cout_group_26,Walloc33bits_1_io_cout_group_25,Walloc33bits_1_io_cout_group_24,
    Walloc33bits_1_io_cout_group_23,Walloc33bits_1_io_cout_group_22,hi_lo_1}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_2 = {Walloc33bits_2_io_cout_group_6,Walloc33bits_2_io_cout_group_5,Walloc33bits_2_io_cout_group_4,
    Walloc33bits_2_io_cout_group_3,Walloc33bits_2_io_cout_group_2,Walloc33bits_2_io_cout_group_1,
    Walloc33bits_2_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_2 = {Walloc33bits_2_io_cout_group_14,Walloc33bits_2_io_cout_group_13,Walloc33bits_2_io_cout_group_12,
    Walloc33bits_2_io_cout_group_11,Walloc33bits_2_io_cout_group_10,Walloc33bits_2_io_cout_group_9,
    Walloc33bits_2_io_cout_group_8,Walloc33bits_2_io_cout_group_7,lo_lo_2}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_2 = {Walloc33bits_2_io_cout_group_21,Walloc33bits_2_io_cout_group_20,Walloc33bits_2_io_cout_group_19,
    Walloc33bits_2_io_cout_group_18,Walloc33bits_2_io_cout_group_17,Walloc33bits_2_io_cout_group_16,
    Walloc33bits_2_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_2 = {Walloc33bits_2_io_cout_group_29,Walloc33bits_2_io_cout_group_28,Walloc33bits_2_io_cout_group_27,
    Walloc33bits_2_io_cout_group_26,Walloc33bits_2_io_cout_group_25,Walloc33bits_2_io_cout_group_24,
    Walloc33bits_2_io_cout_group_23,Walloc33bits_2_io_cout_group_22,hi_lo_2}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_3 = {Walloc33bits_3_io_cout_group_6,Walloc33bits_3_io_cout_group_5,Walloc33bits_3_io_cout_group_4,
    Walloc33bits_3_io_cout_group_3,Walloc33bits_3_io_cout_group_2,Walloc33bits_3_io_cout_group_1,
    Walloc33bits_3_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_3 = {Walloc33bits_3_io_cout_group_14,Walloc33bits_3_io_cout_group_13,Walloc33bits_3_io_cout_group_12,
    Walloc33bits_3_io_cout_group_11,Walloc33bits_3_io_cout_group_10,Walloc33bits_3_io_cout_group_9,
    Walloc33bits_3_io_cout_group_8,Walloc33bits_3_io_cout_group_7,lo_lo_3}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_3 = {Walloc33bits_3_io_cout_group_21,Walloc33bits_3_io_cout_group_20,Walloc33bits_3_io_cout_group_19,
    Walloc33bits_3_io_cout_group_18,Walloc33bits_3_io_cout_group_17,Walloc33bits_3_io_cout_group_16,
    Walloc33bits_3_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_3 = {Walloc33bits_3_io_cout_group_29,Walloc33bits_3_io_cout_group_28,Walloc33bits_3_io_cout_group_27,
    Walloc33bits_3_io_cout_group_26,Walloc33bits_3_io_cout_group_25,Walloc33bits_3_io_cout_group_24,
    Walloc33bits_3_io_cout_group_23,Walloc33bits_3_io_cout_group_22,hi_lo_3}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_4 = {Walloc33bits_4_io_cout_group_6,Walloc33bits_4_io_cout_group_5,Walloc33bits_4_io_cout_group_4,
    Walloc33bits_4_io_cout_group_3,Walloc33bits_4_io_cout_group_2,Walloc33bits_4_io_cout_group_1,
    Walloc33bits_4_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_4 = {Walloc33bits_4_io_cout_group_14,Walloc33bits_4_io_cout_group_13,Walloc33bits_4_io_cout_group_12,
    Walloc33bits_4_io_cout_group_11,Walloc33bits_4_io_cout_group_10,Walloc33bits_4_io_cout_group_9,
    Walloc33bits_4_io_cout_group_8,Walloc33bits_4_io_cout_group_7,lo_lo_4}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_4 = {Walloc33bits_4_io_cout_group_21,Walloc33bits_4_io_cout_group_20,Walloc33bits_4_io_cout_group_19,
    Walloc33bits_4_io_cout_group_18,Walloc33bits_4_io_cout_group_17,Walloc33bits_4_io_cout_group_16,
    Walloc33bits_4_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_4 = {Walloc33bits_4_io_cout_group_29,Walloc33bits_4_io_cout_group_28,Walloc33bits_4_io_cout_group_27,
    Walloc33bits_4_io_cout_group_26,Walloc33bits_4_io_cout_group_25,Walloc33bits_4_io_cout_group_24,
    Walloc33bits_4_io_cout_group_23,Walloc33bits_4_io_cout_group_22,hi_lo_4}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_5 = {Walloc33bits_5_io_cout_group_6,Walloc33bits_5_io_cout_group_5,Walloc33bits_5_io_cout_group_4,
    Walloc33bits_5_io_cout_group_3,Walloc33bits_5_io_cout_group_2,Walloc33bits_5_io_cout_group_1,
    Walloc33bits_5_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_5 = {Walloc33bits_5_io_cout_group_14,Walloc33bits_5_io_cout_group_13,Walloc33bits_5_io_cout_group_12,
    Walloc33bits_5_io_cout_group_11,Walloc33bits_5_io_cout_group_10,Walloc33bits_5_io_cout_group_9,
    Walloc33bits_5_io_cout_group_8,Walloc33bits_5_io_cout_group_7,lo_lo_5}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_5 = {Walloc33bits_5_io_cout_group_21,Walloc33bits_5_io_cout_group_20,Walloc33bits_5_io_cout_group_19,
    Walloc33bits_5_io_cout_group_18,Walloc33bits_5_io_cout_group_17,Walloc33bits_5_io_cout_group_16,
    Walloc33bits_5_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_5 = {Walloc33bits_5_io_cout_group_29,Walloc33bits_5_io_cout_group_28,Walloc33bits_5_io_cout_group_27,
    Walloc33bits_5_io_cout_group_26,Walloc33bits_5_io_cout_group_25,Walloc33bits_5_io_cout_group_24,
    Walloc33bits_5_io_cout_group_23,Walloc33bits_5_io_cout_group_22,hi_lo_5}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_6 = {Walloc33bits_6_io_cout_group_6,Walloc33bits_6_io_cout_group_5,Walloc33bits_6_io_cout_group_4,
    Walloc33bits_6_io_cout_group_3,Walloc33bits_6_io_cout_group_2,Walloc33bits_6_io_cout_group_1,
    Walloc33bits_6_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_6 = {Walloc33bits_6_io_cout_group_14,Walloc33bits_6_io_cout_group_13,Walloc33bits_6_io_cout_group_12,
    Walloc33bits_6_io_cout_group_11,Walloc33bits_6_io_cout_group_10,Walloc33bits_6_io_cout_group_9,
    Walloc33bits_6_io_cout_group_8,Walloc33bits_6_io_cout_group_7,lo_lo_6}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_6 = {Walloc33bits_6_io_cout_group_21,Walloc33bits_6_io_cout_group_20,Walloc33bits_6_io_cout_group_19,
    Walloc33bits_6_io_cout_group_18,Walloc33bits_6_io_cout_group_17,Walloc33bits_6_io_cout_group_16,
    Walloc33bits_6_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_6 = {Walloc33bits_6_io_cout_group_29,Walloc33bits_6_io_cout_group_28,Walloc33bits_6_io_cout_group_27,
    Walloc33bits_6_io_cout_group_26,Walloc33bits_6_io_cout_group_25,Walloc33bits_6_io_cout_group_24,
    Walloc33bits_6_io_cout_group_23,Walloc33bits_6_io_cout_group_22,hi_lo_6}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_7 = {Walloc33bits_7_io_cout_group_6,Walloc33bits_7_io_cout_group_5,Walloc33bits_7_io_cout_group_4,
    Walloc33bits_7_io_cout_group_3,Walloc33bits_7_io_cout_group_2,Walloc33bits_7_io_cout_group_1,
    Walloc33bits_7_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_7 = {Walloc33bits_7_io_cout_group_14,Walloc33bits_7_io_cout_group_13,Walloc33bits_7_io_cout_group_12,
    Walloc33bits_7_io_cout_group_11,Walloc33bits_7_io_cout_group_10,Walloc33bits_7_io_cout_group_9,
    Walloc33bits_7_io_cout_group_8,Walloc33bits_7_io_cout_group_7,lo_lo_7}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_7 = {Walloc33bits_7_io_cout_group_21,Walloc33bits_7_io_cout_group_20,Walloc33bits_7_io_cout_group_19,
    Walloc33bits_7_io_cout_group_18,Walloc33bits_7_io_cout_group_17,Walloc33bits_7_io_cout_group_16,
    Walloc33bits_7_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_7 = {Walloc33bits_7_io_cout_group_29,Walloc33bits_7_io_cout_group_28,Walloc33bits_7_io_cout_group_27,
    Walloc33bits_7_io_cout_group_26,Walloc33bits_7_io_cout_group_25,Walloc33bits_7_io_cout_group_24,
    Walloc33bits_7_io_cout_group_23,Walloc33bits_7_io_cout_group_22,hi_lo_7}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_8 = {Walloc33bits_8_io_cout_group_6,Walloc33bits_8_io_cout_group_5,Walloc33bits_8_io_cout_group_4,
    Walloc33bits_8_io_cout_group_3,Walloc33bits_8_io_cout_group_2,Walloc33bits_8_io_cout_group_1,
    Walloc33bits_8_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_8 = {Walloc33bits_8_io_cout_group_14,Walloc33bits_8_io_cout_group_13,Walloc33bits_8_io_cout_group_12,
    Walloc33bits_8_io_cout_group_11,Walloc33bits_8_io_cout_group_10,Walloc33bits_8_io_cout_group_9,
    Walloc33bits_8_io_cout_group_8,Walloc33bits_8_io_cout_group_7,lo_lo_8}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_8 = {Walloc33bits_8_io_cout_group_21,Walloc33bits_8_io_cout_group_20,Walloc33bits_8_io_cout_group_19,
    Walloc33bits_8_io_cout_group_18,Walloc33bits_8_io_cout_group_17,Walloc33bits_8_io_cout_group_16,
    Walloc33bits_8_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_8 = {Walloc33bits_8_io_cout_group_29,Walloc33bits_8_io_cout_group_28,Walloc33bits_8_io_cout_group_27,
    Walloc33bits_8_io_cout_group_26,Walloc33bits_8_io_cout_group_25,Walloc33bits_8_io_cout_group_24,
    Walloc33bits_8_io_cout_group_23,Walloc33bits_8_io_cout_group_22,hi_lo_8}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_9 = {Walloc33bits_9_io_cout_group_6,Walloc33bits_9_io_cout_group_5,Walloc33bits_9_io_cout_group_4,
    Walloc33bits_9_io_cout_group_3,Walloc33bits_9_io_cout_group_2,Walloc33bits_9_io_cout_group_1,
    Walloc33bits_9_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_9 = {Walloc33bits_9_io_cout_group_14,Walloc33bits_9_io_cout_group_13,Walloc33bits_9_io_cout_group_12,
    Walloc33bits_9_io_cout_group_11,Walloc33bits_9_io_cout_group_10,Walloc33bits_9_io_cout_group_9,
    Walloc33bits_9_io_cout_group_8,Walloc33bits_9_io_cout_group_7,lo_lo_9}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_9 = {Walloc33bits_9_io_cout_group_21,Walloc33bits_9_io_cout_group_20,Walloc33bits_9_io_cout_group_19,
    Walloc33bits_9_io_cout_group_18,Walloc33bits_9_io_cout_group_17,Walloc33bits_9_io_cout_group_16,
    Walloc33bits_9_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_9 = {Walloc33bits_9_io_cout_group_29,Walloc33bits_9_io_cout_group_28,Walloc33bits_9_io_cout_group_27,
    Walloc33bits_9_io_cout_group_26,Walloc33bits_9_io_cout_group_25,Walloc33bits_9_io_cout_group_24,
    Walloc33bits_9_io_cout_group_23,Walloc33bits_9_io_cout_group_22,hi_lo_9}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_10 = {Walloc33bits_10_io_cout_group_6,Walloc33bits_10_io_cout_group_5,Walloc33bits_10_io_cout_group_4
    ,Walloc33bits_10_io_cout_group_3,Walloc33bits_10_io_cout_group_2,Walloc33bits_10_io_cout_group_1,
    Walloc33bits_10_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_10 = {Walloc33bits_10_io_cout_group_14,Walloc33bits_10_io_cout_group_13,
    Walloc33bits_10_io_cout_group_12,Walloc33bits_10_io_cout_group_11,Walloc33bits_10_io_cout_group_10,
    Walloc33bits_10_io_cout_group_9,Walloc33bits_10_io_cout_group_8,Walloc33bits_10_io_cout_group_7,lo_lo_10}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_10 = {Walloc33bits_10_io_cout_group_21,Walloc33bits_10_io_cout_group_20,
    Walloc33bits_10_io_cout_group_19,Walloc33bits_10_io_cout_group_18,Walloc33bits_10_io_cout_group_17,
    Walloc33bits_10_io_cout_group_16,Walloc33bits_10_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_10 = {Walloc33bits_10_io_cout_group_29,Walloc33bits_10_io_cout_group_28,
    Walloc33bits_10_io_cout_group_27,Walloc33bits_10_io_cout_group_26,Walloc33bits_10_io_cout_group_25,
    Walloc33bits_10_io_cout_group_24,Walloc33bits_10_io_cout_group_23,Walloc33bits_10_io_cout_group_22,hi_lo_10}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_11 = {Walloc33bits_11_io_cout_group_6,Walloc33bits_11_io_cout_group_5,Walloc33bits_11_io_cout_group_4
    ,Walloc33bits_11_io_cout_group_3,Walloc33bits_11_io_cout_group_2,Walloc33bits_11_io_cout_group_1,
    Walloc33bits_11_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_11 = {Walloc33bits_11_io_cout_group_14,Walloc33bits_11_io_cout_group_13,
    Walloc33bits_11_io_cout_group_12,Walloc33bits_11_io_cout_group_11,Walloc33bits_11_io_cout_group_10,
    Walloc33bits_11_io_cout_group_9,Walloc33bits_11_io_cout_group_8,Walloc33bits_11_io_cout_group_7,lo_lo_11}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_11 = {Walloc33bits_11_io_cout_group_21,Walloc33bits_11_io_cout_group_20,
    Walloc33bits_11_io_cout_group_19,Walloc33bits_11_io_cout_group_18,Walloc33bits_11_io_cout_group_17,
    Walloc33bits_11_io_cout_group_16,Walloc33bits_11_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_11 = {Walloc33bits_11_io_cout_group_29,Walloc33bits_11_io_cout_group_28,
    Walloc33bits_11_io_cout_group_27,Walloc33bits_11_io_cout_group_26,Walloc33bits_11_io_cout_group_25,
    Walloc33bits_11_io_cout_group_24,Walloc33bits_11_io_cout_group_23,Walloc33bits_11_io_cout_group_22,hi_lo_11}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_12 = {Walloc33bits_12_io_cout_group_6,Walloc33bits_12_io_cout_group_5,Walloc33bits_12_io_cout_group_4
    ,Walloc33bits_12_io_cout_group_3,Walloc33bits_12_io_cout_group_2,Walloc33bits_12_io_cout_group_1,
    Walloc33bits_12_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_12 = {Walloc33bits_12_io_cout_group_14,Walloc33bits_12_io_cout_group_13,
    Walloc33bits_12_io_cout_group_12,Walloc33bits_12_io_cout_group_11,Walloc33bits_12_io_cout_group_10,
    Walloc33bits_12_io_cout_group_9,Walloc33bits_12_io_cout_group_8,Walloc33bits_12_io_cout_group_7,lo_lo_12}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_12 = {Walloc33bits_12_io_cout_group_21,Walloc33bits_12_io_cout_group_20,
    Walloc33bits_12_io_cout_group_19,Walloc33bits_12_io_cout_group_18,Walloc33bits_12_io_cout_group_17,
    Walloc33bits_12_io_cout_group_16,Walloc33bits_12_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_12 = {Walloc33bits_12_io_cout_group_29,Walloc33bits_12_io_cout_group_28,
    Walloc33bits_12_io_cout_group_27,Walloc33bits_12_io_cout_group_26,Walloc33bits_12_io_cout_group_25,
    Walloc33bits_12_io_cout_group_24,Walloc33bits_12_io_cout_group_23,Walloc33bits_12_io_cout_group_22,hi_lo_12}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_13 = {Walloc33bits_13_io_cout_group_6,Walloc33bits_13_io_cout_group_5,Walloc33bits_13_io_cout_group_4
    ,Walloc33bits_13_io_cout_group_3,Walloc33bits_13_io_cout_group_2,Walloc33bits_13_io_cout_group_1,
    Walloc33bits_13_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_13 = {Walloc33bits_13_io_cout_group_14,Walloc33bits_13_io_cout_group_13,
    Walloc33bits_13_io_cout_group_12,Walloc33bits_13_io_cout_group_11,Walloc33bits_13_io_cout_group_10,
    Walloc33bits_13_io_cout_group_9,Walloc33bits_13_io_cout_group_8,Walloc33bits_13_io_cout_group_7,lo_lo_13}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_13 = {Walloc33bits_13_io_cout_group_21,Walloc33bits_13_io_cout_group_20,
    Walloc33bits_13_io_cout_group_19,Walloc33bits_13_io_cout_group_18,Walloc33bits_13_io_cout_group_17,
    Walloc33bits_13_io_cout_group_16,Walloc33bits_13_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_13 = {Walloc33bits_13_io_cout_group_29,Walloc33bits_13_io_cout_group_28,
    Walloc33bits_13_io_cout_group_27,Walloc33bits_13_io_cout_group_26,Walloc33bits_13_io_cout_group_25,
    Walloc33bits_13_io_cout_group_24,Walloc33bits_13_io_cout_group_23,Walloc33bits_13_io_cout_group_22,hi_lo_13}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_14 = {Walloc33bits_14_io_cout_group_6,Walloc33bits_14_io_cout_group_5,Walloc33bits_14_io_cout_group_4
    ,Walloc33bits_14_io_cout_group_3,Walloc33bits_14_io_cout_group_2,Walloc33bits_14_io_cout_group_1,
    Walloc33bits_14_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_14 = {Walloc33bits_14_io_cout_group_14,Walloc33bits_14_io_cout_group_13,
    Walloc33bits_14_io_cout_group_12,Walloc33bits_14_io_cout_group_11,Walloc33bits_14_io_cout_group_10,
    Walloc33bits_14_io_cout_group_9,Walloc33bits_14_io_cout_group_8,Walloc33bits_14_io_cout_group_7,lo_lo_14}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_14 = {Walloc33bits_14_io_cout_group_21,Walloc33bits_14_io_cout_group_20,
    Walloc33bits_14_io_cout_group_19,Walloc33bits_14_io_cout_group_18,Walloc33bits_14_io_cout_group_17,
    Walloc33bits_14_io_cout_group_16,Walloc33bits_14_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_14 = {Walloc33bits_14_io_cout_group_29,Walloc33bits_14_io_cout_group_28,
    Walloc33bits_14_io_cout_group_27,Walloc33bits_14_io_cout_group_26,Walloc33bits_14_io_cout_group_25,
    Walloc33bits_14_io_cout_group_24,Walloc33bits_14_io_cout_group_23,Walloc33bits_14_io_cout_group_22,hi_lo_14}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_15 = {Walloc33bits_15_io_cout_group_6,Walloc33bits_15_io_cout_group_5,Walloc33bits_15_io_cout_group_4
    ,Walloc33bits_15_io_cout_group_3,Walloc33bits_15_io_cout_group_2,Walloc33bits_15_io_cout_group_1,
    Walloc33bits_15_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_15 = {Walloc33bits_15_io_cout_group_14,Walloc33bits_15_io_cout_group_13,
    Walloc33bits_15_io_cout_group_12,Walloc33bits_15_io_cout_group_11,Walloc33bits_15_io_cout_group_10,
    Walloc33bits_15_io_cout_group_9,Walloc33bits_15_io_cout_group_8,Walloc33bits_15_io_cout_group_7,lo_lo_15}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_15 = {Walloc33bits_15_io_cout_group_21,Walloc33bits_15_io_cout_group_20,
    Walloc33bits_15_io_cout_group_19,Walloc33bits_15_io_cout_group_18,Walloc33bits_15_io_cout_group_17,
    Walloc33bits_15_io_cout_group_16,Walloc33bits_15_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_15 = {Walloc33bits_15_io_cout_group_29,Walloc33bits_15_io_cout_group_28,
    Walloc33bits_15_io_cout_group_27,Walloc33bits_15_io_cout_group_26,Walloc33bits_15_io_cout_group_25,
    Walloc33bits_15_io_cout_group_24,Walloc33bits_15_io_cout_group_23,Walloc33bits_15_io_cout_group_22,hi_lo_15}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_16 = {Walloc33bits_16_io_cout_group_6,Walloc33bits_16_io_cout_group_5,Walloc33bits_16_io_cout_group_4
    ,Walloc33bits_16_io_cout_group_3,Walloc33bits_16_io_cout_group_2,Walloc33bits_16_io_cout_group_1,
    Walloc33bits_16_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_16 = {Walloc33bits_16_io_cout_group_14,Walloc33bits_16_io_cout_group_13,
    Walloc33bits_16_io_cout_group_12,Walloc33bits_16_io_cout_group_11,Walloc33bits_16_io_cout_group_10,
    Walloc33bits_16_io_cout_group_9,Walloc33bits_16_io_cout_group_8,Walloc33bits_16_io_cout_group_7,lo_lo_16}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_16 = {Walloc33bits_16_io_cout_group_21,Walloc33bits_16_io_cout_group_20,
    Walloc33bits_16_io_cout_group_19,Walloc33bits_16_io_cout_group_18,Walloc33bits_16_io_cout_group_17,
    Walloc33bits_16_io_cout_group_16,Walloc33bits_16_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_16 = {Walloc33bits_16_io_cout_group_29,Walloc33bits_16_io_cout_group_28,
    Walloc33bits_16_io_cout_group_27,Walloc33bits_16_io_cout_group_26,Walloc33bits_16_io_cout_group_25,
    Walloc33bits_16_io_cout_group_24,Walloc33bits_16_io_cout_group_23,Walloc33bits_16_io_cout_group_22,hi_lo_16}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_17 = {Walloc33bits_17_io_cout_group_6,Walloc33bits_17_io_cout_group_5,Walloc33bits_17_io_cout_group_4
    ,Walloc33bits_17_io_cout_group_3,Walloc33bits_17_io_cout_group_2,Walloc33bits_17_io_cout_group_1,
    Walloc33bits_17_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_17 = {Walloc33bits_17_io_cout_group_14,Walloc33bits_17_io_cout_group_13,
    Walloc33bits_17_io_cout_group_12,Walloc33bits_17_io_cout_group_11,Walloc33bits_17_io_cout_group_10,
    Walloc33bits_17_io_cout_group_9,Walloc33bits_17_io_cout_group_8,Walloc33bits_17_io_cout_group_7,lo_lo_17}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_17 = {Walloc33bits_17_io_cout_group_21,Walloc33bits_17_io_cout_group_20,
    Walloc33bits_17_io_cout_group_19,Walloc33bits_17_io_cout_group_18,Walloc33bits_17_io_cout_group_17,
    Walloc33bits_17_io_cout_group_16,Walloc33bits_17_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_17 = {Walloc33bits_17_io_cout_group_29,Walloc33bits_17_io_cout_group_28,
    Walloc33bits_17_io_cout_group_27,Walloc33bits_17_io_cout_group_26,Walloc33bits_17_io_cout_group_25,
    Walloc33bits_17_io_cout_group_24,Walloc33bits_17_io_cout_group_23,Walloc33bits_17_io_cout_group_22,hi_lo_17}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_18 = {Walloc33bits_18_io_cout_group_6,Walloc33bits_18_io_cout_group_5,Walloc33bits_18_io_cout_group_4
    ,Walloc33bits_18_io_cout_group_3,Walloc33bits_18_io_cout_group_2,Walloc33bits_18_io_cout_group_1,
    Walloc33bits_18_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_18 = {Walloc33bits_18_io_cout_group_14,Walloc33bits_18_io_cout_group_13,
    Walloc33bits_18_io_cout_group_12,Walloc33bits_18_io_cout_group_11,Walloc33bits_18_io_cout_group_10,
    Walloc33bits_18_io_cout_group_9,Walloc33bits_18_io_cout_group_8,Walloc33bits_18_io_cout_group_7,lo_lo_18}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_18 = {Walloc33bits_18_io_cout_group_21,Walloc33bits_18_io_cout_group_20,
    Walloc33bits_18_io_cout_group_19,Walloc33bits_18_io_cout_group_18,Walloc33bits_18_io_cout_group_17,
    Walloc33bits_18_io_cout_group_16,Walloc33bits_18_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_18 = {Walloc33bits_18_io_cout_group_29,Walloc33bits_18_io_cout_group_28,
    Walloc33bits_18_io_cout_group_27,Walloc33bits_18_io_cout_group_26,Walloc33bits_18_io_cout_group_25,
    Walloc33bits_18_io_cout_group_24,Walloc33bits_18_io_cout_group_23,Walloc33bits_18_io_cout_group_22,hi_lo_18}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_19 = {Walloc33bits_19_io_cout_group_6,Walloc33bits_19_io_cout_group_5,Walloc33bits_19_io_cout_group_4
    ,Walloc33bits_19_io_cout_group_3,Walloc33bits_19_io_cout_group_2,Walloc33bits_19_io_cout_group_1,
    Walloc33bits_19_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_19 = {Walloc33bits_19_io_cout_group_14,Walloc33bits_19_io_cout_group_13,
    Walloc33bits_19_io_cout_group_12,Walloc33bits_19_io_cout_group_11,Walloc33bits_19_io_cout_group_10,
    Walloc33bits_19_io_cout_group_9,Walloc33bits_19_io_cout_group_8,Walloc33bits_19_io_cout_group_7,lo_lo_19}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_19 = {Walloc33bits_19_io_cout_group_21,Walloc33bits_19_io_cout_group_20,
    Walloc33bits_19_io_cout_group_19,Walloc33bits_19_io_cout_group_18,Walloc33bits_19_io_cout_group_17,
    Walloc33bits_19_io_cout_group_16,Walloc33bits_19_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_19 = {Walloc33bits_19_io_cout_group_29,Walloc33bits_19_io_cout_group_28,
    Walloc33bits_19_io_cout_group_27,Walloc33bits_19_io_cout_group_26,Walloc33bits_19_io_cout_group_25,
    Walloc33bits_19_io_cout_group_24,Walloc33bits_19_io_cout_group_23,Walloc33bits_19_io_cout_group_22,hi_lo_19}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_20 = {Walloc33bits_20_io_cout_group_6,Walloc33bits_20_io_cout_group_5,Walloc33bits_20_io_cout_group_4
    ,Walloc33bits_20_io_cout_group_3,Walloc33bits_20_io_cout_group_2,Walloc33bits_20_io_cout_group_1,
    Walloc33bits_20_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_20 = {Walloc33bits_20_io_cout_group_14,Walloc33bits_20_io_cout_group_13,
    Walloc33bits_20_io_cout_group_12,Walloc33bits_20_io_cout_group_11,Walloc33bits_20_io_cout_group_10,
    Walloc33bits_20_io_cout_group_9,Walloc33bits_20_io_cout_group_8,Walloc33bits_20_io_cout_group_7,lo_lo_20}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_20 = {Walloc33bits_20_io_cout_group_21,Walloc33bits_20_io_cout_group_20,
    Walloc33bits_20_io_cout_group_19,Walloc33bits_20_io_cout_group_18,Walloc33bits_20_io_cout_group_17,
    Walloc33bits_20_io_cout_group_16,Walloc33bits_20_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_20 = {Walloc33bits_20_io_cout_group_29,Walloc33bits_20_io_cout_group_28,
    Walloc33bits_20_io_cout_group_27,Walloc33bits_20_io_cout_group_26,Walloc33bits_20_io_cout_group_25,
    Walloc33bits_20_io_cout_group_24,Walloc33bits_20_io_cout_group_23,Walloc33bits_20_io_cout_group_22,hi_lo_20}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_21 = {Walloc33bits_21_io_cout_group_6,Walloc33bits_21_io_cout_group_5,Walloc33bits_21_io_cout_group_4
    ,Walloc33bits_21_io_cout_group_3,Walloc33bits_21_io_cout_group_2,Walloc33bits_21_io_cout_group_1,
    Walloc33bits_21_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_21 = {Walloc33bits_21_io_cout_group_14,Walloc33bits_21_io_cout_group_13,
    Walloc33bits_21_io_cout_group_12,Walloc33bits_21_io_cout_group_11,Walloc33bits_21_io_cout_group_10,
    Walloc33bits_21_io_cout_group_9,Walloc33bits_21_io_cout_group_8,Walloc33bits_21_io_cout_group_7,lo_lo_21}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_21 = {Walloc33bits_21_io_cout_group_21,Walloc33bits_21_io_cout_group_20,
    Walloc33bits_21_io_cout_group_19,Walloc33bits_21_io_cout_group_18,Walloc33bits_21_io_cout_group_17,
    Walloc33bits_21_io_cout_group_16,Walloc33bits_21_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_21 = {Walloc33bits_21_io_cout_group_29,Walloc33bits_21_io_cout_group_28,
    Walloc33bits_21_io_cout_group_27,Walloc33bits_21_io_cout_group_26,Walloc33bits_21_io_cout_group_25,
    Walloc33bits_21_io_cout_group_24,Walloc33bits_21_io_cout_group_23,Walloc33bits_21_io_cout_group_22,hi_lo_21}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_22 = {Walloc33bits_22_io_cout_group_6,Walloc33bits_22_io_cout_group_5,Walloc33bits_22_io_cout_group_4
    ,Walloc33bits_22_io_cout_group_3,Walloc33bits_22_io_cout_group_2,Walloc33bits_22_io_cout_group_1,
    Walloc33bits_22_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_22 = {Walloc33bits_22_io_cout_group_14,Walloc33bits_22_io_cout_group_13,
    Walloc33bits_22_io_cout_group_12,Walloc33bits_22_io_cout_group_11,Walloc33bits_22_io_cout_group_10,
    Walloc33bits_22_io_cout_group_9,Walloc33bits_22_io_cout_group_8,Walloc33bits_22_io_cout_group_7,lo_lo_22}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_22 = {Walloc33bits_22_io_cout_group_21,Walloc33bits_22_io_cout_group_20,
    Walloc33bits_22_io_cout_group_19,Walloc33bits_22_io_cout_group_18,Walloc33bits_22_io_cout_group_17,
    Walloc33bits_22_io_cout_group_16,Walloc33bits_22_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_22 = {Walloc33bits_22_io_cout_group_29,Walloc33bits_22_io_cout_group_28,
    Walloc33bits_22_io_cout_group_27,Walloc33bits_22_io_cout_group_26,Walloc33bits_22_io_cout_group_25,
    Walloc33bits_22_io_cout_group_24,Walloc33bits_22_io_cout_group_23,Walloc33bits_22_io_cout_group_22,hi_lo_22}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_23 = {Walloc33bits_23_io_cout_group_6,Walloc33bits_23_io_cout_group_5,Walloc33bits_23_io_cout_group_4
    ,Walloc33bits_23_io_cout_group_3,Walloc33bits_23_io_cout_group_2,Walloc33bits_23_io_cout_group_1,
    Walloc33bits_23_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_23 = {Walloc33bits_23_io_cout_group_14,Walloc33bits_23_io_cout_group_13,
    Walloc33bits_23_io_cout_group_12,Walloc33bits_23_io_cout_group_11,Walloc33bits_23_io_cout_group_10,
    Walloc33bits_23_io_cout_group_9,Walloc33bits_23_io_cout_group_8,Walloc33bits_23_io_cout_group_7,lo_lo_23}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_23 = {Walloc33bits_23_io_cout_group_21,Walloc33bits_23_io_cout_group_20,
    Walloc33bits_23_io_cout_group_19,Walloc33bits_23_io_cout_group_18,Walloc33bits_23_io_cout_group_17,
    Walloc33bits_23_io_cout_group_16,Walloc33bits_23_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_23 = {Walloc33bits_23_io_cout_group_29,Walloc33bits_23_io_cout_group_28,
    Walloc33bits_23_io_cout_group_27,Walloc33bits_23_io_cout_group_26,Walloc33bits_23_io_cout_group_25,
    Walloc33bits_23_io_cout_group_24,Walloc33bits_23_io_cout_group_23,Walloc33bits_23_io_cout_group_22,hi_lo_23}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_24 = {Walloc33bits_24_io_cout_group_6,Walloc33bits_24_io_cout_group_5,Walloc33bits_24_io_cout_group_4
    ,Walloc33bits_24_io_cout_group_3,Walloc33bits_24_io_cout_group_2,Walloc33bits_24_io_cout_group_1,
    Walloc33bits_24_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_24 = {Walloc33bits_24_io_cout_group_14,Walloc33bits_24_io_cout_group_13,
    Walloc33bits_24_io_cout_group_12,Walloc33bits_24_io_cout_group_11,Walloc33bits_24_io_cout_group_10,
    Walloc33bits_24_io_cout_group_9,Walloc33bits_24_io_cout_group_8,Walloc33bits_24_io_cout_group_7,lo_lo_24}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_24 = {Walloc33bits_24_io_cout_group_21,Walloc33bits_24_io_cout_group_20,
    Walloc33bits_24_io_cout_group_19,Walloc33bits_24_io_cout_group_18,Walloc33bits_24_io_cout_group_17,
    Walloc33bits_24_io_cout_group_16,Walloc33bits_24_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_24 = {Walloc33bits_24_io_cout_group_29,Walloc33bits_24_io_cout_group_28,
    Walloc33bits_24_io_cout_group_27,Walloc33bits_24_io_cout_group_26,Walloc33bits_24_io_cout_group_25,
    Walloc33bits_24_io_cout_group_24,Walloc33bits_24_io_cout_group_23,Walloc33bits_24_io_cout_group_22,hi_lo_24}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_25 = {Walloc33bits_25_io_cout_group_6,Walloc33bits_25_io_cout_group_5,Walloc33bits_25_io_cout_group_4
    ,Walloc33bits_25_io_cout_group_3,Walloc33bits_25_io_cout_group_2,Walloc33bits_25_io_cout_group_1,
    Walloc33bits_25_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_25 = {Walloc33bits_25_io_cout_group_14,Walloc33bits_25_io_cout_group_13,
    Walloc33bits_25_io_cout_group_12,Walloc33bits_25_io_cout_group_11,Walloc33bits_25_io_cout_group_10,
    Walloc33bits_25_io_cout_group_9,Walloc33bits_25_io_cout_group_8,Walloc33bits_25_io_cout_group_7,lo_lo_25}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_25 = {Walloc33bits_25_io_cout_group_21,Walloc33bits_25_io_cout_group_20,
    Walloc33bits_25_io_cout_group_19,Walloc33bits_25_io_cout_group_18,Walloc33bits_25_io_cout_group_17,
    Walloc33bits_25_io_cout_group_16,Walloc33bits_25_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_25 = {Walloc33bits_25_io_cout_group_29,Walloc33bits_25_io_cout_group_28,
    Walloc33bits_25_io_cout_group_27,Walloc33bits_25_io_cout_group_26,Walloc33bits_25_io_cout_group_25,
    Walloc33bits_25_io_cout_group_24,Walloc33bits_25_io_cout_group_23,Walloc33bits_25_io_cout_group_22,hi_lo_25}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_26 = {Walloc33bits_26_io_cout_group_6,Walloc33bits_26_io_cout_group_5,Walloc33bits_26_io_cout_group_4
    ,Walloc33bits_26_io_cout_group_3,Walloc33bits_26_io_cout_group_2,Walloc33bits_26_io_cout_group_1,
    Walloc33bits_26_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_26 = {Walloc33bits_26_io_cout_group_14,Walloc33bits_26_io_cout_group_13,
    Walloc33bits_26_io_cout_group_12,Walloc33bits_26_io_cout_group_11,Walloc33bits_26_io_cout_group_10,
    Walloc33bits_26_io_cout_group_9,Walloc33bits_26_io_cout_group_8,Walloc33bits_26_io_cout_group_7,lo_lo_26}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_26 = {Walloc33bits_26_io_cout_group_21,Walloc33bits_26_io_cout_group_20,
    Walloc33bits_26_io_cout_group_19,Walloc33bits_26_io_cout_group_18,Walloc33bits_26_io_cout_group_17,
    Walloc33bits_26_io_cout_group_16,Walloc33bits_26_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_26 = {Walloc33bits_26_io_cout_group_29,Walloc33bits_26_io_cout_group_28,
    Walloc33bits_26_io_cout_group_27,Walloc33bits_26_io_cout_group_26,Walloc33bits_26_io_cout_group_25,
    Walloc33bits_26_io_cout_group_24,Walloc33bits_26_io_cout_group_23,Walloc33bits_26_io_cout_group_22,hi_lo_26}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_27 = {Walloc33bits_27_io_cout_group_6,Walloc33bits_27_io_cout_group_5,Walloc33bits_27_io_cout_group_4
    ,Walloc33bits_27_io_cout_group_3,Walloc33bits_27_io_cout_group_2,Walloc33bits_27_io_cout_group_1,
    Walloc33bits_27_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_27 = {Walloc33bits_27_io_cout_group_14,Walloc33bits_27_io_cout_group_13,
    Walloc33bits_27_io_cout_group_12,Walloc33bits_27_io_cout_group_11,Walloc33bits_27_io_cout_group_10,
    Walloc33bits_27_io_cout_group_9,Walloc33bits_27_io_cout_group_8,Walloc33bits_27_io_cout_group_7,lo_lo_27}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_27 = {Walloc33bits_27_io_cout_group_21,Walloc33bits_27_io_cout_group_20,
    Walloc33bits_27_io_cout_group_19,Walloc33bits_27_io_cout_group_18,Walloc33bits_27_io_cout_group_17,
    Walloc33bits_27_io_cout_group_16,Walloc33bits_27_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_27 = {Walloc33bits_27_io_cout_group_29,Walloc33bits_27_io_cout_group_28,
    Walloc33bits_27_io_cout_group_27,Walloc33bits_27_io_cout_group_26,Walloc33bits_27_io_cout_group_25,
    Walloc33bits_27_io_cout_group_24,Walloc33bits_27_io_cout_group_23,Walloc33bits_27_io_cout_group_22,hi_lo_27}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_28 = {Walloc33bits_28_io_cout_group_6,Walloc33bits_28_io_cout_group_5,Walloc33bits_28_io_cout_group_4
    ,Walloc33bits_28_io_cout_group_3,Walloc33bits_28_io_cout_group_2,Walloc33bits_28_io_cout_group_1,
    Walloc33bits_28_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_28 = {Walloc33bits_28_io_cout_group_14,Walloc33bits_28_io_cout_group_13,
    Walloc33bits_28_io_cout_group_12,Walloc33bits_28_io_cout_group_11,Walloc33bits_28_io_cout_group_10,
    Walloc33bits_28_io_cout_group_9,Walloc33bits_28_io_cout_group_8,Walloc33bits_28_io_cout_group_7,lo_lo_28}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_28 = {Walloc33bits_28_io_cout_group_21,Walloc33bits_28_io_cout_group_20,
    Walloc33bits_28_io_cout_group_19,Walloc33bits_28_io_cout_group_18,Walloc33bits_28_io_cout_group_17,
    Walloc33bits_28_io_cout_group_16,Walloc33bits_28_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_28 = {Walloc33bits_28_io_cout_group_29,Walloc33bits_28_io_cout_group_28,
    Walloc33bits_28_io_cout_group_27,Walloc33bits_28_io_cout_group_26,Walloc33bits_28_io_cout_group_25,
    Walloc33bits_28_io_cout_group_24,Walloc33bits_28_io_cout_group_23,Walloc33bits_28_io_cout_group_22,hi_lo_28}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_29 = {Walloc33bits_29_io_cout_group_6,Walloc33bits_29_io_cout_group_5,Walloc33bits_29_io_cout_group_4
    ,Walloc33bits_29_io_cout_group_3,Walloc33bits_29_io_cout_group_2,Walloc33bits_29_io_cout_group_1,
    Walloc33bits_29_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_29 = {Walloc33bits_29_io_cout_group_14,Walloc33bits_29_io_cout_group_13,
    Walloc33bits_29_io_cout_group_12,Walloc33bits_29_io_cout_group_11,Walloc33bits_29_io_cout_group_10,
    Walloc33bits_29_io_cout_group_9,Walloc33bits_29_io_cout_group_8,Walloc33bits_29_io_cout_group_7,lo_lo_29}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_29 = {Walloc33bits_29_io_cout_group_21,Walloc33bits_29_io_cout_group_20,
    Walloc33bits_29_io_cout_group_19,Walloc33bits_29_io_cout_group_18,Walloc33bits_29_io_cout_group_17,
    Walloc33bits_29_io_cout_group_16,Walloc33bits_29_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_29 = {Walloc33bits_29_io_cout_group_29,Walloc33bits_29_io_cout_group_28,
    Walloc33bits_29_io_cout_group_27,Walloc33bits_29_io_cout_group_26,Walloc33bits_29_io_cout_group_25,
    Walloc33bits_29_io_cout_group_24,Walloc33bits_29_io_cout_group_23,Walloc33bits_29_io_cout_group_22,hi_lo_29}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_30 = {Walloc33bits_30_io_cout_group_6,Walloc33bits_30_io_cout_group_5,Walloc33bits_30_io_cout_group_4
    ,Walloc33bits_30_io_cout_group_3,Walloc33bits_30_io_cout_group_2,Walloc33bits_30_io_cout_group_1,
    Walloc33bits_30_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_30 = {Walloc33bits_30_io_cout_group_14,Walloc33bits_30_io_cout_group_13,
    Walloc33bits_30_io_cout_group_12,Walloc33bits_30_io_cout_group_11,Walloc33bits_30_io_cout_group_10,
    Walloc33bits_30_io_cout_group_9,Walloc33bits_30_io_cout_group_8,Walloc33bits_30_io_cout_group_7,lo_lo_30}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_30 = {Walloc33bits_30_io_cout_group_21,Walloc33bits_30_io_cout_group_20,
    Walloc33bits_30_io_cout_group_19,Walloc33bits_30_io_cout_group_18,Walloc33bits_30_io_cout_group_17,
    Walloc33bits_30_io_cout_group_16,Walloc33bits_30_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_30 = {Walloc33bits_30_io_cout_group_29,Walloc33bits_30_io_cout_group_28,
    Walloc33bits_30_io_cout_group_27,Walloc33bits_30_io_cout_group_26,Walloc33bits_30_io_cout_group_25,
    Walloc33bits_30_io_cout_group_24,Walloc33bits_30_io_cout_group_23,Walloc33bits_30_io_cout_group_22,hi_lo_30}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_31 = {Walloc33bits_31_io_cout_group_6,Walloc33bits_31_io_cout_group_5,Walloc33bits_31_io_cout_group_4
    ,Walloc33bits_31_io_cout_group_3,Walloc33bits_31_io_cout_group_2,Walloc33bits_31_io_cout_group_1,
    Walloc33bits_31_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_31 = {Walloc33bits_31_io_cout_group_14,Walloc33bits_31_io_cout_group_13,
    Walloc33bits_31_io_cout_group_12,Walloc33bits_31_io_cout_group_11,Walloc33bits_31_io_cout_group_10,
    Walloc33bits_31_io_cout_group_9,Walloc33bits_31_io_cout_group_8,Walloc33bits_31_io_cout_group_7,lo_lo_31}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_31 = {Walloc33bits_31_io_cout_group_21,Walloc33bits_31_io_cout_group_20,
    Walloc33bits_31_io_cout_group_19,Walloc33bits_31_io_cout_group_18,Walloc33bits_31_io_cout_group_17,
    Walloc33bits_31_io_cout_group_16,Walloc33bits_31_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_31 = {Walloc33bits_31_io_cout_group_29,Walloc33bits_31_io_cout_group_28,
    Walloc33bits_31_io_cout_group_27,Walloc33bits_31_io_cout_group_26,Walloc33bits_31_io_cout_group_25,
    Walloc33bits_31_io_cout_group_24,Walloc33bits_31_io_cout_group_23,Walloc33bits_31_io_cout_group_22,hi_lo_31}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_32 = {Walloc33bits_32_io_cout_group_6,Walloc33bits_32_io_cout_group_5,Walloc33bits_32_io_cout_group_4
    ,Walloc33bits_32_io_cout_group_3,Walloc33bits_32_io_cout_group_2,Walloc33bits_32_io_cout_group_1,
    Walloc33bits_32_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_32 = {Walloc33bits_32_io_cout_group_14,Walloc33bits_32_io_cout_group_13,
    Walloc33bits_32_io_cout_group_12,Walloc33bits_32_io_cout_group_11,Walloc33bits_32_io_cout_group_10,
    Walloc33bits_32_io_cout_group_9,Walloc33bits_32_io_cout_group_8,Walloc33bits_32_io_cout_group_7,lo_lo_32}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_32 = {Walloc33bits_32_io_cout_group_21,Walloc33bits_32_io_cout_group_20,
    Walloc33bits_32_io_cout_group_19,Walloc33bits_32_io_cout_group_18,Walloc33bits_32_io_cout_group_17,
    Walloc33bits_32_io_cout_group_16,Walloc33bits_32_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_32 = {Walloc33bits_32_io_cout_group_29,Walloc33bits_32_io_cout_group_28,
    Walloc33bits_32_io_cout_group_27,Walloc33bits_32_io_cout_group_26,Walloc33bits_32_io_cout_group_25,
    Walloc33bits_32_io_cout_group_24,Walloc33bits_32_io_cout_group_23,Walloc33bits_32_io_cout_group_22,hi_lo_32}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_33 = {Walloc33bits_33_io_cout_group_6,Walloc33bits_33_io_cout_group_5,Walloc33bits_33_io_cout_group_4
    ,Walloc33bits_33_io_cout_group_3,Walloc33bits_33_io_cout_group_2,Walloc33bits_33_io_cout_group_1,
    Walloc33bits_33_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_33 = {Walloc33bits_33_io_cout_group_14,Walloc33bits_33_io_cout_group_13,
    Walloc33bits_33_io_cout_group_12,Walloc33bits_33_io_cout_group_11,Walloc33bits_33_io_cout_group_10,
    Walloc33bits_33_io_cout_group_9,Walloc33bits_33_io_cout_group_8,Walloc33bits_33_io_cout_group_7,lo_lo_33}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_33 = {Walloc33bits_33_io_cout_group_21,Walloc33bits_33_io_cout_group_20,
    Walloc33bits_33_io_cout_group_19,Walloc33bits_33_io_cout_group_18,Walloc33bits_33_io_cout_group_17,
    Walloc33bits_33_io_cout_group_16,Walloc33bits_33_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_33 = {Walloc33bits_33_io_cout_group_29,Walloc33bits_33_io_cout_group_28,
    Walloc33bits_33_io_cout_group_27,Walloc33bits_33_io_cout_group_26,Walloc33bits_33_io_cout_group_25,
    Walloc33bits_33_io_cout_group_24,Walloc33bits_33_io_cout_group_23,Walloc33bits_33_io_cout_group_22,hi_lo_33}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_34 = {Walloc33bits_34_io_cout_group_6,Walloc33bits_34_io_cout_group_5,Walloc33bits_34_io_cout_group_4
    ,Walloc33bits_34_io_cout_group_3,Walloc33bits_34_io_cout_group_2,Walloc33bits_34_io_cout_group_1,
    Walloc33bits_34_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_34 = {Walloc33bits_34_io_cout_group_14,Walloc33bits_34_io_cout_group_13,
    Walloc33bits_34_io_cout_group_12,Walloc33bits_34_io_cout_group_11,Walloc33bits_34_io_cout_group_10,
    Walloc33bits_34_io_cout_group_9,Walloc33bits_34_io_cout_group_8,Walloc33bits_34_io_cout_group_7,lo_lo_34}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_34 = {Walloc33bits_34_io_cout_group_21,Walloc33bits_34_io_cout_group_20,
    Walloc33bits_34_io_cout_group_19,Walloc33bits_34_io_cout_group_18,Walloc33bits_34_io_cout_group_17,
    Walloc33bits_34_io_cout_group_16,Walloc33bits_34_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_34 = {Walloc33bits_34_io_cout_group_29,Walloc33bits_34_io_cout_group_28,
    Walloc33bits_34_io_cout_group_27,Walloc33bits_34_io_cout_group_26,Walloc33bits_34_io_cout_group_25,
    Walloc33bits_34_io_cout_group_24,Walloc33bits_34_io_cout_group_23,Walloc33bits_34_io_cout_group_22,hi_lo_34}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_35 = {Walloc33bits_35_io_cout_group_6,Walloc33bits_35_io_cout_group_5,Walloc33bits_35_io_cout_group_4
    ,Walloc33bits_35_io_cout_group_3,Walloc33bits_35_io_cout_group_2,Walloc33bits_35_io_cout_group_1,
    Walloc33bits_35_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_35 = {Walloc33bits_35_io_cout_group_14,Walloc33bits_35_io_cout_group_13,
    Walloc33bits_35_io_cout_group_12,Walloc33bits_35_io_cout_group_11,Walloc33bits_35_io_cout_group_10,
    Walloc33bits_35_io_cout_group_9,Walloc33bits_35_io_cout_group_8,Walloc33bits_35_io_cout_group_7,lo_lo_35}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_35 = {Walloc33bits_35_io_cout_group_21,Walloc33bits_35_io_cout_group_20,
    Walloc33bits_35_io_cout_group_19,Walloc33bits_35_io_cout_group_18,Walloc33bits_35_io_cout_group_17,
    Walloc33bits_35_io_cout_group_16,Walloc33bits_35_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_35 = {Walloc33bits_35_io_cout_group_29,Walloc33bits_35_io_cout_group_28,
    Walloc33bits_35_io_cout_group_27,Walloc33bits_35_io_cout_group_26,Walloc33bits_35_io_cout_group_25,
    Walloc33bits_35_io_cout_group_24,Walloc33bits_35_io_cout_group_23,Walloc33bits_35_io_cout_group_22,hi_lo_35}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_36 = {Walloc33bits_36_io_cout_group_6,Walloc33bits_36_io_cout_group_5,Walloc33bits_36_io_cout_group_4
    ,Walloc33bits_36_io_cout_group_3,Walloc33bits_36_io_cout_group_2,Walloc33bits_36_io_cout_group_1,
    Walloc33bits_36_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_36 = {Walloc33bits_36_io_cout_group_14,Walloc33bits_36_io_cout_group_13,
    Walloc33bits_36_io_cout_group_12,Walloc33bits_36_io_cout_group_11,Walloc33bits_36_io_cout_group_10,
    Walloc33bits_36_io_cout_group_9,Walloc33bits_36_io_cout_group_8,Walloc33bits_36_io_cout_group_7,lo_lo_36}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_36 = {Walloc33bits_36_io_cout_group_21,Walloc33bits_36_io_cout_group_20,
    Walloc33bits_36_io_cout_group_19,Walloc33bits_36_io_cout_group_18,Walloc33bits_36_io_cout_group_17,
    Walloc33bits_36_io_cout_group_16,Walloc33bits_36_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_36 = {Walloc33bits_36_io_cout_group_29,Walloc33bits_36_io_cout_group_28,
    Walloc33bits_36_io_cout_group_27,Walloc33bits_36_io_cout_group_26,Walloc33bits_36_io_cout_group_25,
    Walloc33bits_36_io_cout_group_24,Walloc33bits_36_io_cout_group_23,Walloc33bits_36_io_cout_group_22,hi_lo_36}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_37 = {Walloc33bits_37_io_cout_group_6,Walloc33bits_37_io_cout_group_5,Walloc33bits_37_io_cout_group_4
    ,Walloc33bits_37_io_cout_group_3,Walloc33bits_37_io_cout_group_2,Walloc33bits_37_io_cout_group_1,
    Walloc33bits_37_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_37 = {Walloc33bits_37_io_cout_group_14,Walloc33bits_37_io_cout_group_13,
    Walloc33bits_37_io_cout_group_12,Walloc33bits_37_io_cout_group_11,Walloc33bits_37_io_cout_group_10,
    Walloc33bits_37_io_cout_group_9,Walloc33bits_37_io_cout_group_8,Walloc33bits_37_io_cout_group_7,lo_lo_37}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_37 = {Walloc33bits_37_io_cout_group_21,Walloc33bits_37_io_cout_group_20,
    Walloc33bits_37_io_cout_group_19,Walloc33bits_37_io_cout_group_18,Walloc33bits_37_io_cout_group_17,
    Walloc33bits_37_io_cout_group_16,Walloc33bits_37_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_37 = {Walloc33bits_37_io_cout_group_29,Walloc33bits_37_io_cout_group_28,
    Walloc33bits_37_io_cout_group_27,Walloc33bits_37_io_cout_group_26,Walloc33bits_37_io_cout_group_25,
    Walloc33bits_37_io_cout_group_24,Walloc33bits_37_io_cout_group_23,Walloc33bits_37_io_cout_group_22,hi_lo_37}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_38 = {Walloc33bits_38_io_cout_group_6,Walloc33bits_38_io_cout_group_5,Walloc33bits_38_io_cout_group_4
    ,Walloc33bits_38_io_cout_group_3,Walloc33bits_38_io_cout_group_2,Walloc33bits_38_io_cout_group_1,
    Walloc33bits_38_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_38 = {Walloc33bits_38_io_cout_group_14,Walloc33bits_38_io_cout_group_13,
    Walloc33bits_38_io_cout_group_12,Walloc33bits_38_io_cout_group_11,Walloc33bits_38_io_cout_group_10,
    Walloc33bits_38_io_cout_group_9,Walloc33bits_38_io_cout_group_8,Walloc33bits_38_io_cout_group_7,lo_lo_38}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_38 = {Walloc33bits_38_io_cout_group_21,Walloc33bits_38_io_cout_group_20,
    Walloc33bits_38_io_cout_group_19,Walloc33bits_38_io_cout_group_18,Walloc33bits_38_io_cout_group_17,
    Walloc33bits_38_io_cout_group_16,Walloc33bits_38_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_38 = {Walloc33bits_38_io_cout_group_29,Walloc33bits_38_io_cout_group_28,
    Walloc33bits_38_io_cout_group_27,Walloc33bits_38_io_cout_group_26,Walloc33bits_38_io_cout_group_25,
    Walloc33bits_38_io_cout_group_24,Walloc33bits_38_io_cout_group_23,Walloc33bits_38_io_cout_group_22,hi_lo_38}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_39 = {Walloc33bits_39_io_cout_group_6,Walloc33bits_39_io_cout_group_5,Walloc33bits_39_io_cout_group_4
    ,Walloc33bits_39_io_cout_group_3,Walloc33bits_39_io_cout_group_2,Walloc33bits_39_io_cout_group_1,
    Walloc33bits_39_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_39 = {Walloc33bits_39_io_cout_group_14,Walloc33bits_39_io_cout_group_13,
    Walloc33bits_39_io_cout_group_12,Walloc33bits_39_io_cout_group_11,Walloc33bits_39_io_cout_group_10,
    Walloc33bits_39_io_cout_group_9,Walloc33bits_39_io_cout_group_8,Walloc33bits_39_io_cout_group_7,lo_lo_39}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_39 = {Walloc33bits_39_io_cout_group_21,Walloc33bits_39_io_cout_group_20,
    Walloc33bits_39_io_cout_group_19,Walloc33bits_39_io_cout_group_18,Walloc33bits_39_io_cout_group_17,
    Walloc33bits_39_io_cout_group_16,Walloc33bits_39_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_39 = {Walloc33bits_39_io_cout_group_29,Walloc33bits_39_io_cout_group_28,
    Walloc33bits_39_io_cout_group_27,Walloc33bits_39_io_cout_group_26,Walloc33bits_39_io_cout_group_25,
    Walloc33bits_39_io_cout_group_24,Walloc33bits_39_io_cout_group_23,Walloc33bits_39_io_cout_group_22,hi_lo_39}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_40 = {Walloc33bits_40_io_cout_group_6,Walloc33bits_40_io_cout_group_5,Walloc33bits_40_io_cout_group_4
    ,Walloc33bits_40_io_cout_group_3,Walloc33bits_40_io_cout_group_2,Walloc33bits_40_io_cout_group_1,
    Walloc33bits_40_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_40 = {Walloc33bits_40_io_cout_group_14,Walloc33bits_40_io_cout_group_13,
    Walloc33bits_40_io_cout_group_12,Walloc33bits_40_io_cout_group_11,Walloc33bits_40_io_cout_group_10,
    Walloc33bits_40_io_cout_group_9,Walloc33bits_40_io_cout_group_8,Walloc33bits_40_io_cout_group_7,lo_lo_40}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_40 = {Walloc33bits_40_io_cout_group_21,Walloc33bits_40_io_cout_group_20,
    Walloc33bits_40_io_cout_group_19,Walloc33bits_40_io_cout_group_18,Walloc33bits_40_io_cout_group_17,
    Walloc33bits_40_io_cout_group_16,Walloc33bits_40_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_40 = {Walloc33bits_40_io_cout_group_29,Walloc33bits_40_io_cout_group_28,
    Walloc33bits_40_io_cout_group_27,Walloc33bits_40_io_cout_group_26,Walloc33bits_40_io_cout_group_25,
    Walloc33bits_40_io_cout_group_24,Walloc33bits_40_io_cout_group_23,Walloc33bits_40_io_cout_group_22,hi_lo_40}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_41 = {Walloc33bits_41_io_cout_group_6,Walloc33bits_41_io_cout_group_5,Walloc33bits_41_io_cout_group_4
    ,Walloc33bits_41_io_cout_group_3,Walloc33bits_41_io_cout_group_2,Walloc33bits_41_io_cout_group_1,
    Walloc33bits_41_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_41 = {Walloc33bits_41_io_cout_group_14,Walloc33bits_41_io_cout_group_13,
    Walloc33bits_41_io_cout_group_12,Walloc33bits_41_io_cout_group_11,Walloc33bits_41_io_cout_group_10,
    Walloc33bits_41_io_cout_group_9,Walloc33bits_41_io_cout_group_8,Walloc33bits_41_io_cout_group_7,lo_lo_41}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_41 = {Walloc33bits_41_io_cout_group_21,Walloc33bits_41_io_cout_group_20,
    Walloc33bits_41_io_cout_group_19,Walloc33bits_41_io_cout_group_18,Walloc33bits_41_io_cout_group_17,
    Walloc33bits_41_io_cout_group_16,Walloc33bits_41_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_41 = {Walloc33bits_41_io_cout_group_29,Walloc33bits_41_io_cout_group_28,
    Walloc33bits_41_io_cout_group_27,Walloc33bits_41_io_cout_group_26,Walloc33bits_41_io_cout_group_25,
    Walloc33bits_41_io_cout_group_24,Walloc33bits_41_io_cout_group_23,Walloc33bits_41_io_cout_group_22,hi_lo_41}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_42 = {Walloc33bits_42_io_cout_group_6,Walloc33bits_42_io_cout_group_5,Walloc33bits_42_io_cout_group_4
    ,Walloc33bits_42_io_cout_group_3,Walloc33bits_42_io_cout_group_2,Walloc33bits_42_io_cout_group_1,
    Walloc33bits_42_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_42 = {Walloc33bits_42_io_cout_group_14,Walloc33bits_42_io_cout_group_13,
    Walloc33bits_42_io_cout_group_12,Walloc33bits_42_io_cout_group_11,Walloc33bits_42_io_cout_group_10,
    Walloc33bits_42_io_cout_group_9,Walloc33bits_42_io_cout_group_8,Walloc33bits_42_io_cout_group_7,lo_lo_42}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_42 = {Walloc33bits_42_io_cout_group_21,Walloc33bits_42_io_cout_group_20,
    Walloc33bits_42_io_cout_group_19,Walloc33bits_42_io_cout_group_18,Walloc33bits_42_io_cout_group_17,
    Walloc33bits_42_io_cout_group_16,Walloc33bits_42_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_42 = {Walloc33bits_42_io_cout_group_29,Walloc33bits_42_io_cout_group_28,
    Walloc33bits_42_io_cout_group_27,Walloc33bits_42_io_cout_group_26,Walloc33bits_42_io_cout_group_25,
    Walloc33bits_42_io_cout_group_24,Walloc33bits_42_io_cout_group_23,Walloc33bits_42_io_cout_group_22,hi_lo_42}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_43 = {Walloc33bits_43_io_cout_group_6,Walloc33bits_43_io_cout_group_5,Walloc33bits_43_io_cout_group_4
    ,Walloc33bits_43_io_cout_group_3,Walloc33bits_43_io_cout_group_2,Walloc33bits_43_io_cout_group_1,
    Walloc33bits_43_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_43 = {Walloc33bits_43_io_cout_group_14,Walloc33bits_43_io_cout_group_13,
    Walloc33bits_43_io_cout_group_12,Walloc33bits_43_io_cout_group_11,Walloc33bits_43_io_cout_group_10,
    Walloc33bits_43_io_cout_group_9,Walloc33bits_43_io_cout_group_8,Walloc33bits_43_io_cout_group_7,lo_lo_43}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_43 = {Walloc33bits_43_io_cout_group_21,Walloc33bits_43_io_cout_group_20,
    Walloc33bits_43_io_cout_group_19,Walloc33bits_43_io_cout_group_18,Walloc33bits_43_io_cout_group_17,
    Walloc33bits_43_io_cout_group_16,Walloc33bits_43_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_43 = {Walloc33bits_43_io_cout_group_29,Walloc33bits_43_io_cout_group_28,
    Walloc33bits_43_io_cout_group_27,Walloc33bits_43_io_cout_group_26,Walloc33bits_43_io_cout_group_25,
    Walloc33bits_43_io_cout_group_24,Walloc33bits_43_io_cout_group_23,Walloc33bits_43_io_cout_group_22,hi_lo_43}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_44 = {Walloc33bits_44_io_cout_group_6,Walloc33bits_44_io_cout_group_5,Walloc33bits_44_io_cout_group_4
    ,Walloc33bits_44_io_cout_group_3,Walloc33bits_44_io_cout_group_2,Walloc33bits_44_io_cout_group_1,
    Walloc33bits_44_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_44 = {Walloc33bits_44_io_cout_group_14,Walloc33bits_44_io_cout_group_13,
    Walloc33bits_44_io_cout_group_12,Walloc33bits_44_io_cout_group_11,Walloc33bits_44_io_cout_group_10,
    Walloc33bits_44_io_cout_group_9,Walloc33bits_44_io_cout_group_8,Walloc33bits_44_io_cout_group_7,lo_lo_44}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_44 = {Walloc33bits_44_io_cout_group_21,Walloc33bits_44_io_cout_group_20,
    Walloc33bits_44_io_cout_group_19,Walloc33bits_44_io_cout_group_18,Walloc33bits_44_io_cout_group_17,
    Walloc33bits_44_io_cout_group_16,Walloc33bits_44_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_44 = {Walloc33bits_44_io_cout_group_29,Walloc33bits_44_io_cout_group_28,
    Walloc33bits_44_io_cout_group_27,Walloc33bits_44_io_cout_group_26,Walloc33bits_44_io_cout_group_25,
    Walloc33bits_44_io_cout_group_24,Walloc33bits_44_io_cout_group_23,Walloc33bits_44_io_cout_group_22,hi_lo_44}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_45 = {Walloc33bits_45_io_cout_group_6,Walloc33bits_45_io_cout_group_5,Walloc33bits_45_io_cout_group_4
    ,Walloc33bits_45_io_cout_group_3,Walloc33bits_45_io_cout_group_2,Walloc33bits_45_io_cout_group_1,
    Walloc33bits_45_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_45 = {Walloc33bits_45_io_cout_group_14,Walloc33bits_45_io_cout_group_13,
    Walloc33bits_45_io_cout_group_12,Walloc33bits_45_io_cout_group_11,Walloc33bits_45_io_cout_group_10,
    Walloc33bits_45_io_cout_group_9,Walloc33bits_45_io_cout_group_8,Walloc33bits_45_io_cout_group_7,lo_lo_45}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_45 = {Walloc33bits_45_io_cout_group_21,Walloc33bits_45_io_cout_group_20,
    Walloc33bits_45_io_cout_group_19,Walloc33bits_45_io_cout_group_18,Walloc33bits_45_io_cout_group_17,
    Walloc33bits_45_io_cout_group_16,Walloc33bits_45_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_45 = {Walloc33bits_45_io_cout_group_29,Walloc33bits_45_io_cout_group_28,
    Walloc33bits_45_io_cout_group_27,Walloc33bits_45_io_cout_group_26,Walloc33bits_45_io_cout_group_25,
    Walloc33bits_45_io_cout_group_24,Walloc33bits_45_io_cout_group_23,Walloc33bits_45_io_cout_group_22,hi_lo_45}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_46 = {Walloc33bits_46_io_cout_group_6,Walloc33bits_46_io_cout_group_5,Walloc33bits_46_io_cout_group_4
    ,Walloc33bits_46_io_cout_group_3,Walloc33bits_46_io_cout_group_2,Walloc33bits_46_io_cout_group_1,
    Walloc33bits_46_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_46 = {Walloc33bits_46_io_cout_group_14,Walloc33bits_46_io_cout_group_13,
    Walloc33bits_46_io_cout_group_12,Walloc33bits_46_io_cout_group_11,Walloc33bits_46_io_cout_group_10,
    Walloc33bits_46_io_cout_group_9,Walloc33bits_46_io_cout_group_8,Walloc33bits_46_io_cout_group_7,lo_lo_46}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_46 = {Walloc33bits_46_io_cout_group_21,Walloc33bits_46_io_cout_group_20,
    Walloc33bits_46_io_cout_group_19,Walloc33bits_46_io_cout_group_18,Walloc33bits_46_io_cout_group_17,
    Walloc33bits_46_io_cout_group_16,Walloc33bits_46_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_46 = {Walloc33bits_46_io_cout_group_29,Walloc33bits_46_io_cout_group_28,
    Walloc33bits_46_io_cout_group_27,Walloc33bits_46_io_cout_group_26,Walloc33bits_46_io_cout_group_25,
    Walloc33bits_46_io_cout_group_24,Walloc33bits_46_io_cout_group_23,Walloc33bits_46_io_cout_group_22,hi_lo_46}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_47 = {Walloc33bits_47_io_cout_group_6,Walloc33bits_47_io_cout_group_5,Walloc33bits_47_io_cout_group_4
    ,Walloc33bits_47_io_cout_group_3,Walloc33bits_47_io_cout_group_2,Walloc33bits_47_io_cout_group_1,
    Walloc33bits_47_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_47 = {Walloc33bits_47_io_cout_group_14,Walloc33bits_47_io_cout_group_13,
    Walloc33bits_47_io_cout_group_12,Walloc33bits_47_io_cout_group_11,Walloc33bits_47_io_cout_group_10,
    Walloc33bits_47_io_cout_group_9,Walloc33bits_47_io_cout_group_8,Walloc33bits_47_io_cout_group_7,lo_lo_47}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_47 = {Walloc33bits_47_io_cout_group_21,Walloc33bits_47_io_cout_group_20,
    Walloc33bits_47_io_cout_group_19,Walloc33bits_47_io_cout_group_18,Walloc33bits_47_io_cout_group_17,
    Walloc33bits_47_io_cout_group_16,Walloc33bits_47_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_47 = {Walloc33bits_47_io_cout_group_29,Walloc33bits_47_io_cout_group_28,
    Walloc33bits_47_io_cout_group_27,Walloc33bits_47_io_cout_group_26,Walloc33bits_47_io_cout_group_25,
    Walloc33bits_47_io_cout_group_24,Walloc33bits_47_io_cout_group_23,Walloc33bits_47_io_cout_group_22,hi_lo_47}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_48 = {Walloc33bits_48_io_cout_group_6,Walloc33bits_48_io_cout_group_5,Walloc33bits_48_io_cout_group_4
    ,Walloc33bits_48_io_cout_group_3,Walloc33bits_48_io_cout_group_2,Walloc33bits_48_io_cout_group_1,
    Walloc33bits_48_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_48 = {Walloc33bits_48_io_cout_group_14,Walloc33bits_48_io_cout_group_13,
    Walloc33bits_48_io_cout_group_12,Walloc33bits_48_io_cout_group_11,Walloc33bits_48_io_cout_group_10,
    Walloc33bits_48_io_cout_group_9,Walloc33bits_48_io_cout_group_8,Walloc33bits_48_io_cout_group_7,lo_lo_48}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_48 = {Walloc33bits_48_io_cout_group_21,Walloc33bits_48_io_cout_group_20,
    Walloc33bits_48_io_cout_group_19,Walloc33bits_48_io_cout_group_18,Walloc33bits_48_io_cout_group_17,
    Walloc33bits_48_io_cout_group_16,Walloc33bits_48_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_48 = {Walloc33bits_48_io_cout_group_29,Walloc33bits_48_io_cout_group_28,
    Walloc33bits_48_io_cout_group_27,Walloc33bits_48_io_cout_group_26,Walloc33bits_48_io_cout_group_25,
    Walloc33bits_48_io_cout_group_24,Walloc33bits_48_io_cout_group_23,Walloc33bits_48_io_cout_group_22,hi_lo_48}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_49 = {Walloc33bits_49_io_cout_group_6,Walloc33bits_49_io_cout_group_5,Walloc33bits_49_io_cout_group_4
    ,Walloc33bits_49_io_cout_group_3,Walloc33bits_49_io_cout_group_2,Walloc33bits_49_io_cout_group_1,
    Walloc33bits_49_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_49 = {Walloc33bits_49_io_cout_group_14,Walloc33bits_49_io_cout_group_13,
    Walloc33bits_49_io_cout_group_12,Walloc33bits_49_io_cout_group_11,Walloc33bits_49_io_cout_group_10,
    Walloc33bits_49_io_cout_group_9,Walloc33bits_49_io_cout_group_8,Walloc33bits_49_io_cout_group_7,lo_lo_49}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_49 = {Walloc33bits_49_io_cout_group_21,Walloc33bits_49_io_cout_group_20,
    Walloc33bits_49_io_cout_group_19,Walloc33bits_49_io_cout_group_18,Walloc33bits_49_io_cout_group_17,
    Walloc33bits_49_io_cout_group_16,Walloc33bits_49_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_49 = {Walloc33bits_49_io_cout_group_29,Walloc33bits_49_io_cout_group_28,
    Walloc33bits_49_io_cout_group_27,Walloc33bits_49_io_cout_group_26,Walloc33bits_49_io_cout_group_25,
    Walloc33bits_49_io_cout_group_24,Walloc33bits_49_io_cout_group_23,Walloc33bits_49_io_cout_group_22,hi_lo_49}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_50 = {Walloc33bits_50_io_cout_group_6,Walloc33bits_50_io_cout_group_5,Walloc33bits_50_io_cout_group_4
    ,Walloc33bits_50_io_cout_group_3,Walloc33bits_50_io_cout_group_2,Walloc33bits_50_io_cout_group_1,
    Walloc33bits_50_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_50 = {Walloc33bits_50_io_cout_group_14,Walloc33bits_50_io_cout_group_13,
    Walloc33bits_50_io_cout_group_12,Walloc33bits_50_io_cout_group_11,Walloc33bits_50_io_cout_group_10,
    Walloc33bits_50_io_cout_group_9,Walloc33bits_50_io_cout_group_8,Walloc33bits_50_io_cout_group_7,lo_lo_50}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_50 = {Walloc33bits_50_io_cout_group_21,Walloc33bits_50_io_cout_group_20,
    Walloc33bits_50_io_cout_group_19,Walloc33bits_50_io_cout_group_18,Walloc33bits_50_io_cout_group_17,
    Walloc33bits_50_io_cout_group_16,Walloc33bits_50_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_50 = {Walloc33bits_50_io_cout_group_29,Walloc33bits_50_io_cout_group_28,
    Walloc33bits_50_io_cout_group_27,Walloc33bits_50_io_cout_group_26,Walloc33bits_50_io_cout_group_25,
    Walloc33bits_50_io_cout_group_24,Walloc33bits_50_io_cout_group_23,Walloc33bits_50_io_cout_group_22,hi_lo_50}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_51 = {Walloc33bits_51_io_cout_group_6,Walloc33bits_51_io_cout_group_5,Walloc33bits_51_io_cout_group_4
    ,Walloc33bits_51_io_cout_group_3,Walloc33bits_51_io_cout_group_2,Walloc33bits_51_io_cout_group_1,
    Walloc33bits_51_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_51 = {Walloc33bits_51_io_cout_group_14,Walloc33bits_51_io_cout_group_13,
    Walloc33bits_51_io_cout_group_12,Walloc33bits_51_io_cout_group_11,Walloc33bits_51_io_cout_group_10,
    Walloc33bits_51_io_cout_group_9,Walloc33bits_51_io_cout_group_8,Walloc33bits_51_io_cout_group_7,lo_lo_51}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_51 = {Walloc33bits_51_io_cout_group_21,Walloc33bits_51_io_cout_group_20,
    Walloc33bits_51_io_cout_group_19,Walloc33bits_51_io_cout_group_18,Walloc33bits_51_io_cout_group_17,
    Walloc33bits_51_io_cout_group_16,Walloc33bits_51_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_51 = {Walloc33bits_51_io_cout_group_29,Walloc33bits_51_io_cout_group_28,
    Walloc33bits_51_io_cout_group_27,Walloc33bits_51_io_cout_group_26,Walloc33bits_51_io_cout_group_25,
    Walloc33bits_51_io_cout_group_24,Walloc33bits_51_io_cout_group_23,Walloc33bits_51_io_cout_group_22,hi_lo_51}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_52 = {Walloc33bits_52_io_cout_group_6,Walloc33bits_52_io_cout_group_5,Walloc33bits_52_io_cout_group_4
    ,Walloc33bits_52_io_cout_group_3,Walloc33bits_52_io_cout_group_2,Walloc33bits_52_io_cout_group_1,
    Walloc33bits_52_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_52 = {Walloc33bits_52_io_cout_group_14,Walloc33bits_52_io_cout_group_13,
    Walloc33bits_52_io_cout_group_12,Walloc33bits_52_io_cout_group_11,Walloc33bits_52_io_cout_group_10,
    Walloc33bits_52_io_cout_group_9,Walloc33bits_52_io_cout_group_8,Walloc33bits_52_io_cout_group_7,lo_lo_52}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_52 = {Walloc33bits_52_io_cout_group_21,Walloc33bits_52_io_cout_group_20,
    Walloc33bits_52_io_cout_group_19,Walloc33bits_52_io_cout_group_18,Walloc33bits_52_io_cout_group_17,
    Walloc33bits_52_io_cout_group_16,Walloc33bits_52_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_52 = {Walloc33bits_52_io_cout_group_29,Walloc33bits_52_io_cout_group_28,
    Walloc33bits_52_io_cout_group_27,Walloc33bits_52_io_cout_group_26,Walloc33bits_52_io_cout_group_25,
    Walloc33bits_52_io_cout_group_24,Walloc33bits_52_io_cout_group_23,Walloc33bits_52_io_cout_group_22,hi_lo_52}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_53 = {Walloc33bits_53_io_cout_group_6,Walloc33bits_53_io_cout_group_5,Walloc33bits_53_io_cout_group_4
    ,Walloc33bits_53_io_cout_group_3,Walloc33bits_53_io_cout_group_2,Walloc33bits_53_io_cout_group_1,
    Walloc33bits_53_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_53 = {Walloc33bits_53_io_cout_group_14,Walloc33bits_53_io_cout_group_13,
    Walloc33bits_53_io_cout_group_12,Walloc33bits_53_io_cout_group_11,Walloc33bits_53_io_cout_group_10,
    Walloc33bits_53_io_cout_group_9,Walloc33bits_53_io_cout_group_8,Walloc33bits_53_io_cout_group_7,lo_lo_53}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_53 = {Walloc33bits_53_io_cout_group_21,Walloc33bits_53_io_cout_group_20,
    Walloc33bits_53_io_cout_group_19,Walloc33bits_53_io_cout_group_18,Walloc33bits_53_io_cout_group_17,
    Walloc33bits_53_io_cout_group_16,Walloc33bits_53_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_53 = {Walloc33bits_53_io_cout_group_29,Walloc33bits_53_io_cout_group_28,
    Walloc33bits_53_io_cout_group_27,Walloc33bits_53_io_cout_group_26,Walloc33bits_53_io_cout_group_25,
    Walloc33bits_53_io_cout_group_24,Walloc33bits_53_io_cout_group_23,Walloc33bits_53_io_cout_group_22,hi_lo_53}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_54 = {Walloc33bits_54_io_cout_group_6,Walloc33bits_54_io_cout_group_5,Walloc33bits_54_io_cout_group_4
    ,Walloc33bits_54_io_cout_group_3,Walloc33bits_54_io_cout_group_2,Walloc33bits_54_io_cout_group_1,
    Walloc33bits_54_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_54 = {Walloc33bits_54_io_cout_group_14,Walloc33bits_54_io_cout_group_13,
    Walloc33bits_54_io_cout_group_12,Walloc33bits_54_io_cout_group_11,Walloc33bits_54_io_cout_group_10,
    Walloc33bits_54_io_cout_group_9,Walloc33bits_54_io_cout_group_8,Walloc33bits_54_io_cout_group_7,lo_lo_54}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_54 = {Walloc33bits_54_io_cout_group_21,Walloc33bits_54_io_cout_group_20,
    Walloc33bits_54_io_cout_group_19,Walloc33bits_54_io_cout_group_18,Walloc33bits_54_io_cout_group_17,
    Walloc33bits_54_io_cout_group_16,Walloc33bits_54_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_54 = {Walloc33bits_54_io_cout_group_29,Walloc33bits_54_io_cout_group_28,
    Walloc33bits_54_io_cout_group_27,Walloc33bits_54_io_cout_group_26,Walloc33bits_54_io_cout_group_25,
    Walloc33bits_54_io_cout_group_24,Walloc33bits_54_io_cout_group_23,Walloc33bits_54_io_cout_group_22,hi_lo_54}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_55 = {Walloc33bits_55_io_cout_group_6,Walloc33bits_55_io_cout_group_5,Walloc33bits_55_io_cout_group_4
    ,Walloc33bits_55_io_cout_group_3,Walloc33bits_55_io_cout_group_2,Walloc33bits_55_io_cout_group_1,
    Walloc33bits_55_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_55 = {Walloc33bits_55_io_cout_group_14,Walloc33bits_55_io_cout_group_13,
    Walloc33bits_55_io_cout_group_12,Walloc33bits_55_io_cout_group_11,Walloc33bits_55_io_cout_group_10,
    Walloc33bits_55_io_cout_group_9,Walloc33bits_55_io_cout_group_8,Walloc33bits_55_io_cout_group_7,lo_lo_55}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_55 = {Walloc33bits_55_io_cout_group_21,Walloc33bits_55_io_cout_group_20,
    Walloc33bits_55_io_cout_group_19,Walloc33bits_55_io_cout_group_18,Walloc33bits_55_io_cout_group_17,
    Walloc33bits_55_io_cout_group_16,Walloc33bits_55_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_55 = {Walloc33bits_55_io_cout_group_29,Walloc33bits_55_io_cout_group_28,
    Walloc33bits_55_io_cout_group_27,Walloc33bits_55_io_cout_group_26,Walloc33bits_55_io_cout_group_25,
    Walloc33bits_55_io_cout_group_24,Walloc33bits_55_io_cout_group_23,Walloc33bits_55_io_cout_group_22,hi_lo_55}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_56 = {Walloc33bits_56_io_cout_group_6,Walloc33bits_56_io_cout_group_5,Walloc33bits_56_io_cout_group_4
    ,Walloc33bits_56_io_cout_group_3,Walloc33bits_56_io_cout_group_2,Walloc33bits_56_io_cout_group_1,
    Walloc33bits_56_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_56 = {Walloc33bits_56_io_cout_group_14,Walloc33bits_56_io_cout_group_13,
    Walloc33bits_56_io_cout_group_12,Walloc33bits_56_io_cout_group_11,Walloc33bits_56_io_cout_group_10,
    Walloc33bits_56_io_cout_group_9,Walloc33bits_56_io_cout_group_8,Walloc33bits_56_io_cout_group_7,lo_lo_56}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_56 = {Walloc33bits_56_io_cout_group_21,Walloc33bits_56_io_cout_group_20,
    Walloc33bits_56_io_cout_group_19,Walloc33bits_56_io_cout_group_18,Walloc33bits_56_io_cout_group_17,
    Walloc33bits_56_io_cout_group_16,Walloc33bits_56_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_56 = {Walloc33bits_56_io_cout_group_29,Walloc33bits_56_io_cout_group_28,
    Walloc33bits_56_io_cout_group_27,Walloc33bits_56_io_cout_group_26,Walloc33bits_56_io_cout_group_25,
    Walloc33bits_56_io_cout_group_24,Walloc33bits_56_io_cout_group_23,Walloc33bits_56_io_cout_group_22,hi_lo_56}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_57 = {Walloc33bits_57_io_cout_group_6,Walloc33bits_57_io_cout_group_5,Walloc33bits_57_io_cout_group_4
    ,Walloc33bits_57_io_cout_group_3,Walloc33bits_57_io_cout_group_2,Walloc33bits_57_io_cout_group_1,
    Walloc33bits_57_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_57 = {Walloc33bits_57_io_cout_group_14,Walloc33bits_57_io_cout_group_13,
    Walloc33bits_57_io_cout_group_12,Walloc33bits_57_io_cout_group_11,Walloc33bits_57_io_cout_group_10,
    Walloc33bits_57_io_cout_group_9,Walloc33bits_57_io_cout_group_8,Walloc33bits_57_io_cout_group_7,lo_lo_57}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_57 = {Walloc33bits_57_io_cout_group_21,Walloc33bits_57_io_cout_group_20,
    Walloc33bits_57_io_cout_group_19,Walloc33bits_57_io_cout_group_18,Walloc33bits_57_io_cout_group_17,
    Walloc33bits_57_io_cout_group_16,Walloc33bits_57_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_57 = {Walloc33bits_57_io_cout_group_29,Walloc33bits_57_io_cout_group_28,
    Walloc33bits_57_io_cout_group_27,Walloc33bits_57_io_cout_group_26,Walloc33bits_57_io_cout_group_25,
    Walloc33bits_57_io_cout_group_24,Walloc33bits_57_io_cout_group_23,Walloc33bits_57_io_cout_group_22,hi_lo_57}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_58 = {Walloc33bits_58_io_cout_group_6,Walloc33bits_58_io_cout_group_5,Walloc33bits_58_io_cout_group_4
    ,Walloc33bits_58_io_cout_group_3,Walloc33bits_58_io_cout_group_2,Walloc33bits_58_io_cout_group_1,
    Walloc33bits_58_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_58 = {Walloc33bits_58_io_cout_group_14,Walloc33bits_58_io_cout_group_13,
    Walloc33bits_58_io_cout_group_12,Walloc33bits_58_io_cout_group_11,Walloc33bits_58_io_cout_group_10,
    Walloc33bits_58_io_cout_group_9,Walloc33bits_58_io_cout_group_8,Walloc33bits_58_io_cout_group_7,lo_lo_58}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_58 = {Walloc33bits_58_io_cout_group_21,Walloc33bits_58_io_cout_group_20,
    Walloc33bits_58_io_cout_group_19,Walloc33bits_58_io_cout_group_18,Walloc33bits_58_io_cout_group_17,
    Walloc33bits_58_io_cout_group_16,Walloc33bits_58_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_58 = {Walloc33bits_58_io_cout_group_29,Walloc33bits_58_io_cout_group_28,
    Walloc33bits_58_io_cout_group_27,Walloc33bits_58_io_cout_group_26,Walloc33bits_58_io_cout_group_25,
    Walloc33bits_58_io_cout_group_24,Walloc33bits_58_io_cout_group_23,Walloc33bits_58_io_cout_group_22,hi_lo_58}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_59 = {Walloc33bits_59_io_cout_group_6,Walloc33bits_59_io_cout_group_5,Walloc33bits_59_io_cout_group_4
    ,Walloc33bits_59_io_cout_group_3,Walloc33bits_59_io_cout_group_2,Walloc33bits_59_io_cout_group_1,
    Walloc33bits_59_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_59 = {Walloc33bits_59_io_cout_group_14,Walloc33bits_59_io_cout_group_13,
    Walloc33bits_59_io_cout_group_12,Walloc33bits_59_io_cout_group_11,Walloc33bits_59_io_cout_group_10,
    Walloc33bits_59_io_cout_group_9,Walloc33bits_59_io_cout_group_8,Walloc33bits_59_io_cout_group_7,lo_lo_59}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_59 = {Walloc33bits_59_io_cout_group_21,Walloc33bits_59_io_cout_group_20,
    Walloc33bits_59_io_cout_group_19,Walloc33bits_59_io_cout_group_18,Walloc33bits_59_io_cout_group_17,
    Walloc33bits_59_io_cout_group_16,Walloc33bits_59_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_59 = {Walloc33bits_59_io_cout_group_29,Walloc33bits_59_io_cout_group_28,
    Walloc33bits_59_io_cout_group_27,Walloc33bits_59_io_cout_group_26,Walloc33bits_59_io_cout_group_25,
    Walloc33bits_59_io_cout_group_24,Walloc33bits_59_io_cout_group_23,Walloc33bits_59_io_cout_group_22,hi_lo_59}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_60 = {Walloc33bits_60_io_cout_group_6,Walloc33bits_60_io_cout_group_5,Walloc33bits_60_io_cout_group_4
    ,Walloc33bits_60_io_cout_group_3,Walloc33bits_60_io_cout_group_2,Walloc33bits_60_io_cout_group_1,
    Walloc33bits_60_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_60 = {Walloc33bits_60_io_cout_group_14,Walloc33bits_60_io_cout_group_13,
    Walloc33bits_60_io_cout_group_12,Walloc33bits_60_io_cout_group_11,Walloc33bits_60_io_cout_group_10,
    Walloc33bits_60_io_cout_group_9,Walloc33bits_60_io_cout_group_8,Walloc33bits_60_io_cout_group_7,lo_lo_60}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_60 = {Walloc33bits_60_io_cout_group_21,Walloc33bits_60_io_cout_group_20,
    Walloc33bits_60_io_cout_group_19,Walloc33bits_60_io_cout_group_18,Walloc33bits_60_io_cout_group_17,
    Walloc33bits_60_io_cout_group_16,Walloc33bits_60_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_60 = {Walloc33bits_60_io_cout_group_29,Walloc33bits_60_io_cout_group_28,
    Walloc33bits_60_io_cout_group_27,Walloc33bits_60_io_cout_group_26,Walloc33bits_60_io_cout_group_25,
    Walloc33bits_60_io_cout_group_24,Walloc33bits_60_io_cout_group_23,Walloc33bits_60_io_cout_group_22,hi_lo_60}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_61 = {Walloc33bits_61_io_cout_group_6,Walloc33bits_61_io_cout_group_5,Walloc33bits_61_io_cout_group_4
    ,Walloc33bits_61_io_cout_group_3,Walloc33bits_61_io_cout_group_2,Walloc33bits_61_io_cout_group_1,
    Walloc33bits_61_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_61 = {Walloc33bits_61_io_cout_group_14,Walloc33bits_61_io_cout_group_13,
    Walloc33bits_61_io_cout_group_12,Walloc33bits_61_io_cout_group_11,Walloc33bits_61_io_cout_group_10,
    Walloc33bits_61_io_cout_group_9,Walloc33bits_61_io_cout_group_8,Walloc33bits_61_io_cout_group_7,lo_lo_61}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_61 = {Walloc33bits_61_io_cout_group_21,Walloc33bits_61_io_cout_group_20,
    Walloc33bits_61_io_cout_group_19,Walloc33bits_61_io_cout_group_18,Walloc33bits_61_io_cout_group_17,
    Walloc33bits_61_io_cout_group_16,Walloc33bits_61_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_61 = {Walloc33bits_61_io_cout_group_29,Walloc33bits_61_io_cout_group_28,
    Walloc33bits_61_io_cout_group_27,Walloc33bits_61_io_cout_group_26,Walloc33bits_61_io_cout_group_25,
    Walloc33bits_61_io_cout_group_24,Walloc33bits_61_io_cout_group_23,Walloc33bits_61_io_cout_group_22,hi_lo_61}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_62 = {Walloc33bits_62_io_cout_group_6,Walloc33bits_62_io_cout_group_5,Walloc33bits_62_io_cout_group_4
    ,Walloc33bits_62_io_cout_group_3,Walloc33bits_62_io_cout_group_2,Walloc33bits_62_io_cout_group_1,
    Walloc33bits_62_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_62 = {Walloc33bits_62_io_cout_group_14,Walloc33bits_62_io_cout_group_13,
    Walloc33bits_62_io_cout_group_12,Walloc33bits_62_io_cout_group_11,Walloc33bits_62_io_cout_group_10,
    Walloc33bits_62_io_cout_group_9,Walloc33bits_62_io_cout_group_8,Walloc33bits_62_io_cout_group_7,lo_lo_62}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_62 = {Walloc33bits_62_io_cout_group_21,Walloc33bits_62_io_cout_group_20,
    Walloc33bits_62_io_cout_group_19,Walloc33bits_62_io_cout_group_18,Walloc33bits_62_io_cout_group_17,
    Walloc33bits_62_io_cout_group_16,Walloc33bits_62_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_62 = {Walloc33bits_62_io_cout_group_29,Walloc33bits_62_io_cout_group_28,
    Walloc33bits_62_io_cout_group_27,Walloc33bits_62_io_cout_group_26,Walloc33bits_62_io_cout_group_25,
    Walloc33bits_62_io_cout_group_24,Walloc33bits_62_io_cout_group_23,Walloc33bits_62_io_cout_group_22,hi_lo_62}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_63 = {Walloc33bits_63_io_cout_group_6,Walloc33bits_63_io_cout_group_5,Walloc33bits_63_io_cout_group_4
    ,Walloc33bits_63_io_cout_group_3,Walloc33bits_63_io_cout_group_2,Walloc33bits_63_io_cout_group_1,
    Walloc33bits_63_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_63 = {Walloc33bits_63_io_cout_group_14,Walloc33bits_63_io_cout_group_13,
    Walloc33bits_63_io_cout_group_12,Walloc33bits_63_io_cout_group_11,Walloc33bits_63_io_cout_group_10,
    Walloc33bits_63_io_cout_group_9,Walloc33bits_63_io_cout_group_8,Walloc33bits_63_io_cout_group_7,lo_lo_63}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_63 = {Walloc33bits_63_io_cout_group_21,Walloc33bits_63_io_cout_group_20,
    Walloc33bits_63_io_cout_group_19,Walloc33bits_63_io_cout_group_18,Walloc33bits_63_io_cout_group_17,
    Walloc33bits_63_io_cout_group_16,Walloc33bits_63_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_63 = {Walloc33bits_63_io_cout_group_29,Walloc33bits_63_io_cout_group_28,
    Walloc33bits_63_io_cout_group_27,Walloc33bits_63_io_cout_group_26,Walloc33bits_63_io_cout_group_25,
    Walloc33bits_63_io_cout_group_24,Walloc33bits_63_io_cout_group_23,Walloc33bits_63_io_cout_group_22,hi_lo_63}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_64 = {Walloc33bits_64_io_cout_group_6,Walloc33bits_64_io_cout_group_5,Walloc33bits_64_io_cout_group_4
    ,Walloc33bits_64_io_cout_group_3,Walloc33bits_64_io_cout_group_2,Walloc33bits_64_io_cout_group_1,
    Walloc33bits_64_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_64 = {Walloc33bits_64_io_cout_group_14,Walloc33bits_64_io_cout_group_13,
    Walloc33bits_64_io_cout_group_12,Walloc33bits_64_io_cout_group_11,Walloc33bits_64_io_cout_group_10,
    Walloc33bits_64_io_cout_group_9,Walloc33bits_64_io_cout_group_8,Walloc33bits_64_io_cout_group_7,lo_lo_64}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_64 = {Walloc33bits_64_io_cout_group_21,Walloc33bits_64_io_cout_group_20,
    Walloc33bits_64_io_cout_group_19,Walloc33bits_64_io_cout_group_18,Walloc33bits_64_io_cout_group_17,
    Walloc33bits_64_io_cout_group_16,Walloc33bits_64_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_64 = {Walloc33bits_64_io_cout_group_29,Walloc33bits_64_io_cout_group_28,
    Walloc33bits_64_io_cout_group_27,Walloc33bits_64_io_cout_group_26,Walloc33bits_64_io_cout_group_25,
    Walloc33bits_64_io_cout_group_24,Walloc33bits_64_io_cout_group_23,Walloc33bits_64_io_cout_group_22,hi_lo_64}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_65 = {Walloc33bits_65_io_cout_group_6,Walloc33bits_65_io_cout_group_5,Walloc33bits_65_io_cout_group_4
    ,Walloc33bits_65_io_cout_group_3,Walloc33bits_65_io_cout_group_2,Walloc33bits_65_io_cout_group_1,
    Walloc33bits_65_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_65 = {Walloc33bits_65_io_cout_group_14,Walloc33bits_65_io_cout_group_13,
    Walloc33bits_65_io_cout_group_12,Walloc33bits_65_io_cout_group_11,Walloc33bits_65_io_cout_group_10,
    Walloc33bits_65_io_cout_group_9,Walloc33bits_65_io_cout_group_8,Walloc33bits_65_io_cout_group_7,lo_lo_65}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_65 = {Walloc33bits_65_io_cout_group_21,Walloc33bits_65_io_cout_group_20,
    Walloc33bits_65_io_cout_group_19,Walloc33bits_65_io_cout_group_18,Walloc33bits_65_io_cout_group_17,
    Walloc33bits_65_io_cout_group_16,Walloc33bits_65_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_65 = {Walloc33bits_65_io_cout_group_29,Walloc33bits_65_io_cout_group_28,
    Walloc33bits_65_io_cout_group_27,Walloc33bits_65_io_cout_group_26,Walloc33bits_65_io_cout_group_25,
    Walloc33bits_65_io_cout_group_24,Walloc33bits_65_io_cout_group_23,Walloc33bits_65_io_cout_group_22,hi_lo_65}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_66 = {Walloc33bits_66_io_cout_group_6,Walloc33bits_66_io_cout_group_5,Walloc33bits_66_io_cout_group_4
    ,Walloc33bits_66_io_cout_group_3,Walloc33bits_66_io_cout_group_2,Walloc33bits_66_io_cout_group_1,
    Walloc33bits_66_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_66 = {Walloc33bits_66_io_cout_group_14,Walloc33bits_66_io_cout_group_13,
    Walloc33bits_66_io_cout_group_12,Walloc33bits_66_io_cout_group_11,Walloc33bits_66_io_cout_group_10,
    Walloc33bits_66_io_cout_group_9,Walloc33bits_66_io_cout_group_8,Walloc33bits_66_io_cout_group_7,lo_lo_66}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_66 = {Walloc33bits_66_io_cout_group_21,Walloc33bits_66_io_cout_group_20,
    Walloc33bits_66_io_cout_group_19,Walloc33bits_66_io_cout_group_18,Walloc33bits_66_io_cout_group_17,
    Walloc33bits_66_io_cout_group_16,Walloc33bits_66_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_66 = {Walloc33bits_66_io_cout_group_29,Walloc33bits_66_io_cout_group_28,
    Walloc33bits_66_io_cout_group_27,Walloc33bits_66_io_cout_group_26,Walloc33bits_66_io_cout_group_25,
    Walloc33bits_66_io_cout_group_24,Walloc33bits_66_io_cout_group_23,Walloc33bits_66_io_cout_group_22,hi_lo_66}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_67 = {Walloc33bits_67_io_cout_group_6,Walloc33bits_67_io_cout_group_5,Walloc33bits_67_io_cout_group_4
    ,Walloc33bits_67_io_cout_group_3,Walloc33bits_67_io_cout_group_2,Walloc33bits_67_io_cout_group_1,
    Walloc33bits_67_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_67 = {Walloc33bits_67_io_cout_group_14,Walloc33bits_67_io_cout_group_13,
    Walloc33bits_67_io_cout_group_12,Walloc33bits_67_io_cout_group_11,Walloc33bits_67_io_cout_group_10,
    Walloc33bits_67_io_cout_group_9,Walloc33bits_67_io_cout_group_8,Walloc33bits_67_io_cout_group_7,lo_lo_67}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_67 = {Walloc33bits_67_io_cout_group_21,Walloc33bits_67_io_cout_group_20,
    Walloc33bits_67_io_cout_group_19,Walloc33bits_67_io_cout_group_18,Walloc33bits_67_io_cout_group_17,
    Walloc33bits_67_io_cout_group_16,Walloc33bits_67_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_67 = {Walloc33bits_67_io_cout_group_29,Walloc33bits_67_io_cout_group_28,
    Walloc33bits_67_io_cout_group_27,Walloc33bits_67_io_cout_group_26,Walloc33bits_67_io_cout_group_25,
    Walloc33bits_67_io_cout_group_24,Walloc33bits_67_io_cout_group_23,Walloc33bits_67_io_cout_group_22,hi_lo_67}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_68 = {Walloc33bits_68_io_cout_group_6,Walloc33bits_68_io_cout_group_5,Walloc33bits_68_io_cout_group_4
    ,Walloc33bits_68_io_cout_group_3,Walloc33bits_68_io_cout_group_2,Walloc33bits_68_io_cout_group_1,
    Walloc33bits_68_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_68 = {Walloc33bits_68_io_cout_group_14,Walloc33bits_68_io_cout_group_13,
    Walloc33bits_68_io_cout_group_12,Walloc33bits_68_io_cout_group_11,Walloc33bits_68_io_cout_group_10,
    Walloc33bits_68_io_cout_group_9,Walloc33bits_68_io_cout_group_8,Walloc33bits_68_io_cout_group_7,lo_lo_68}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_68 = {Walloc33bits_68_io_cout_group_21,Walloc33bits_68_io_cout_group_20,
    Walloc33bits_68_io_cout_group_19,Walloc33bits_68_io_cout_group_18,Walloc33bits_68_io_cout_group_17,
    Walloc33bits_68_io_cout_group_16,Walloc33bits_68_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_68 = {Walloc33bits_68_io_cout_group_29,Walloc33bits_68_io_cout_group_28,
    Walloc33bits_68_io_cout_group_27,Walloc33bits_68_io_cout_group_26,Walloc33bits_68_io_cout_group_25,
    Walloc33bits_68_io_cout_group_24,Walloc33bits_68_io_cout_group_23,Walloc33bits_68_io_cout_group_22,hi_lo_68}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_69 = {Walloc33bits_69_io_cout_group_6,Walloc33bits_69_io_cout_group_5,Walloc33bits_69_io_cout_group_4
    ,Walloc33bits_69_io_cout_group_3,Walloc33bits_69_io_cout_group_2,Walloc33bits_69_io_cout_group_1,
    Walloc33bits_69_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_69 = {Walloc33bits_69_io_cout_group_14,Walloc33bits_69_io_cout_group_13,
    Walloc33bits_69_io_cout_group_12,Walloc33bits_69_io_cout_group_11,Walloc33bits_69_io_cout_group_10,
    Walloc33bits_69_io_cout_group_9,Walloc33bits_69_io_cout_group_8,Walloc33bits_69_io_cout_group_7,lo_lo_69}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_69 = {Walloc33bits_69_io_cout_group_21,Walloc33bits_69_io_cout_group_20,
    Walloc33bits_69_io_cout_group_19,Walloc33bits_69_io_cout_group_18,Walloc33bits_69_io_cout_group_17,
    Walloc33bits_69_io_cout_group_16,Walloc33bits_69_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_69 = {Walloc33bits_69_io_cout_group_29,Walloc33bits_69_io_cout_group_28,
    Walloc33bits_69_io_cout_group_27,Walloc33bits_69_io_cout_group_26,Walloc33bits_69_io_cout_group_25,
    Walloc33bits_69_io_cout_group_24,Walloc33bits_69_io_cout_group_23,Walloc33bits_69_io_cout_group_22,hi_lo_69}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_70 = {Walloc33bits_70_io_cout_group_6,Walloc33bits_70_io_cout_group_5,Walloc33bits_70_io_cout_group_4
    ,Walloc33bits_70_io_cout_group_3,Walloc33bits_70_io_cout_group_2,Walloc33bits_70_io_cout_group_1,
    Walloc33bits_70_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_70 = {Walloc33bits_70_io_cout_group_14,Walloc33bits_70_io_cout_group_13,
    Walloc33bits_70_io_cout_group_12,Walloc33bits_70_io_cout_group_11,Walloc33bits_70_io_cout_group_10,
    Walloc33bits_70_io_cout_group_9,Walloc33bits_70_io_cout_group_8,Walloc33bits_70_io_cout_group_7,lo_lo_70}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_70 = {Walloc33bits_70_io_cout_group_21,Walloc33bits_70_io_cout_group_20,
    Walloc33bits_70_io_cout_group_19,Walloc33bits_70_io_cout_group_18,Walloc33bits_70_io_cout_group_17,
    Walloc33bits_70_io_cout_group_16,Walloc33bits_70_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_70 = {Walloc33bits_70_io_cout_group_29,Walloc33bits_70_io_cout_group_28,
    Walloc33bits_70_io_cout_group_27,Walloc33bits_70_io_cout_group_26,Walloc33bits_70_io_cout_group_25,
    Walloc33bits_70_io_cout_group_24,Walloc33bits_70_io_cout_group_23,Walloc33bits_70_io_cout_group_22,hi_lo_70}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_71 = {Walloc33bits_71_io_cout_group_6,Walloc33bits_71_io_cout_group_5,Walloc33bits_71_io_cout_group_4
    ,Walloc33bits_71_io_cout_group_3,Walloc33bits_71_io_cout_group_2,Walloc33bits_71_io_cout_group_1,
    Walloc33bits_71_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_71 = {Walloc33bits_71_io_cout_group_14,Walloc33bits_71_io_cout_group_13,
    Walloc33bits_71_io_cout_group_12,Walloc33bits_71_io_cout_group_11,Walloc33bits_71_io_cout_group_10,
    Walloc33bits_71_io_cout_group_9,Walloc33bits_71_io_cout_group_8,Walloc33bits_71_io_cout_group_7,lo_lo_71}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_71 = {Walloc33bits_71_io_cout_group_21,Walloc33bits_71_io_cout_group_20,
    Walloc33bits_71_io_cout_group_19,Walloc33bits_71_io_cout_group_18,Walloc33bits_71_io_cout_group_17,
    Walloc33bits_71_io_cout_group_16,Walloc33bits_71_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_71 = {Walloc33bits_71_io_cout_group_29,Walloc33bits_71_io_cout_group_28,
    Walloc33bits_71_io_cout_group_27,Walloc33bits_71_io_cout_group_26,Walloc33bits_71_io_cout_group_25,
    Walloc33bits_71_io_cout_group_24,Walloc33bits_71_io_cout_group_23,Walloc33bits_71_io_cout_group_22,hi_lo_71}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_72 = {Walloc33bits_72_io_cout_group_6,Walloc33bits_72_io_cout_group_5,Walloc33bits_72_io_cout_group_4
    ,Walloc33bits_72_io_cout_group_3,Walloc33bits_72_io_cout_group_2,Walloc33bits_72_io_cout_group_1,
    Walloc33bits_72_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_72 = {Walloc33bits_72_io_cout_group_14,Walloc33bits_72_io_cout_group_13,
    Walloc33bits_72_io_cout_group_12,Walloc33bits_72_io_cout_group_11,Walloc33bits_72_io_cout_group_10,
    Walloc33bits_72_io_cout_group_9,Walloc33bits_72_io_cout_group_8,Walloc33bits_72_io_cout_group_7,lo_lo_72}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_72 = {Walloc33bits_72_io_cout_group_21,Walloc33bits_72_io_cout_group_20,
    Walloc33bits_72_io_cout_group_19,Walloc33bits_72_io_cout_group_18,Walloc33bits_72_io_cout_group_17,
    Walloc33bits_72_io_cout_group_16,Walloc33bits_72_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_72 = {Walloc33bits_72_io_cout_group_29,Walloc33bits_72_io_cout_group_28,
    Walloc33bits_72_io_cout_group_27,Walloc33bits_72_io_cout_group_26,Walloc33bits_72_io_cout_group_25,
    Walloc33bits_72_io_cout_group_24,Walloc33bits_72_io_cout_group_23,Walloc33bits_72_io_cout_group_22,hi_lo_72}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_73 = {Walloc33bits_73_io_cout_group_6,Walloc33bits_73_io_cout_group_5,Walloc33bits_73_io_cout_group_4
    ,Walloc33bits_73_io_cout_group_3,Walloc33bits_73_io_cout_group_2,Walloc33bits_73_io_cout_group_1,
    Walloc33bits_73_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_73 = {Walloc33bits_73_io_cout_group_14,Walloc33bits_73_io_cout_group_13,
    Walloc33bits_73_io_cout_group_12,Walloc33bits_73_io_cout_group_11,Walloc33bits_73_io_cout_group_10,
    Walloc33bits_73_io_cout_group_9,Walloc33bits_73_io_cout_group_8,Walloc33bits_73_io_cout_group_7,lo_lo_73}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_73 = {Walloc33bits_73_io_cout_group_21,Walloc33bits_73_io_cout_group_20,
    Walloc33bits_73_io_cout_group_19,Walloc33bits_73_io_cout_group_18,Walloc33bits_73_io_cout_group_17,
    Walloc33bits_73_io_cout_group_16,Walloc33bits_73_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_73 = {Walloc33bits_73_io_cout_group_29,Walloc33bits_73_io_cout_group_28,
    Walloc33bits_73_io_cout_group_27,Walloc33bits_73_io_cout_group_26,Walloc33bits_73_io_cout_group_25,
    Walloc33bits_73_io_cout_group_24,Walloc33bits_73_io_cout_group_23,Walloc33bits_73_io_cout_group_22,hi_lo_73}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_74 = {Walloc33bits_74_io_cout_group_6,Walloc33bits_74_io_cout_group_5,Walloc33bits_74_io_cout_group_4
    ,Walloc33bits_74_io_cout_group_3,Walloc33bits_74_io_cout_group_2,Walloc33bits_74_io_cout_group_1,
    Walloc33bits_74_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_74 = {Walloc33bits_74_io_cout_group_14,Walloc33bits_74_io_cout_group_13,
    Walloc33bits_74_io_cout_group_12,Walloc33bits_74_io_cout_group_11,Walloc33bits_74_io_cout_group_10,
    Walloc33bits_74_io_cout_group_9,Walloc33bits_74_io_cout_group_8,Walloc33bits_74_io_cout_group_7,lo_lo_74}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_74 = {Walloc33bits_74_io_cout_group_21,Walloc33bits_74_io_cout_group_20,
    Walloc33bits_74_io_cout_group_19,Walloc33bits_74_io_cout_group_18,Walloc33bits_74_io_cout_group_17,
    Walloc33bits_74_io_cout_group_16,Walloc33bits_74_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_74 = {Walloc33bits_74_io_cout_group_29,Walloc33bits_74_io_cout_group_28,
    Walloc33bits_74_io_cout_group_27,Walloc33bits_74_io_cout_group_26,Walloc33bits_74_io_cout_group_25,
    Walloc33bits_74_io_cout_group_24,Walloc33bits_74_io_cout_group_23,Walloc33bits_74_io_cout_group_22,hi_lo_74}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_75 = {Walloc33bits_75_io_cout_group_6,Walloc33bits_75_io_cout_group_5,Walloc33bits_75_io_cout_group_4
    ,Walloc33bits_75_io_cout_group_3,Walloc33bits_75_io_cout_group_2,Walloc33bits_75_io_cout_group_1,
    Walloc33bits_75_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_75 = {Walloc33bits_75_io_cout_group_14,Walloc33bits_75_io_cout_group_13,
    Walloc33bits_75_io_cout_group_12,Walloc33bits_75_io_cout_group_11,Walloc33bits_75_io_cout_group_10,
    Walloc33bits_75_io_cout_group_9,Walloc33bits_75_io_cout_group_8,Walloc33bits_75_io_cout_group_7,lo_lo_75}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_75 = {Walloc33bits_75_io_cout_group_21,Walloc33bits_75_io_cout_group_20,
    Walloc33bits_75_io_cout_group_19,Walloc33bits_75_io_cout_group_18,Walloc33bits_75_io_cout_group_17,
    Walloc33bits_75_io_cout_group_16,Walloc33bits_75_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_75 = {Walloc33bits_75_io_cout_group_29,Walloc33bits_75_io_cout_group_28,
    Walloc33bits_75_io_cout_group_27,Walloc33bits_75_io_cout_group_26,Walloc33bits_75_io_cout_group_25,
    Walloc33bits_75_io_cout_group_24,Walloc33bits_75_io_cout_group_23,Walloc33bits_75_io_cout_group_22,hi_lo_75}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_76 = {Walloc33bits_76_io_cout_group_6,Walloc33bits_76_io_cout_group_5,Walloc33bits_76_io_cout_group_4
    ,Walloc33bits_76_io_cout_group_3,Walloc33bits_76_io_cout_group_2,Walloc33bits_76_io_cout_group_1,
    Walloc33bits_76_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_76 = {Walloc33bits_76_io_cout_group_14,Walloc33bits_76_io_cout_group_13,
    Walloc33bits_76_io_cout_group_12,Walloc33bits_76_io_cout_group_11,Walloc33bits_76_io_cout_group_10,
    Walloc33bits_76_io_cout_group_9,Walloc33bits_76_io_cout_group_8,Walloc33bits_76_io_cout_group_7,lo_lo_76}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_76 = {Walloc33bits_76_io_cout_group_21,Walloc33bits_76_io_cout_group_20,
    Walloc33bits_76_io_cout_group_19,Walloc33bits_76_io_cout_group_18,Walloc33bits_76_io_cout_group_17,
    Walloc33bits_76_io_cout_group_16,Walloc33bits_76_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_76 = {Walloc33bits_76_io_cout_group_29,Walloc33bits_76_io_cout_group_28,
    Walloc33bits_76_io_cout_group_27,Walloc33bits_76_io_cout_group_26,Walloc33bits_76_io_cout_group_25,
    Walloc33bits_76_io_cout_group_24,Walloc33bits_76_io_cout_group_23,Walloc33bits_76_io_cout_group_22,hi_lo_76}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_77 = {Walloc33bits_77_io_cout_group_6,Walloc33bits_77_io_cout_group_5,Walloc33bits_77_io_cout_group_4
    ,Walloc33bits_77_io_cout_group_3,Walloc33bits_77_io_cout_group_2,Walloc33bits_77_io_cout_group_1,
    Walloc33bits_77_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_77 = {Walloc33bits_77_io_cout_group_14,Walloc33bits_77_io_cout_group_13,
    Walloc33bits_77_io_cout_group_12,Walloc33bits_77_io_cout_group_11,Walloc33bits_77_io_cout_group_10,
    Walloc33bits_77_io_cout_group_9,Walloc33bits_77_io_cout_group_8,Walloc33bits_77_io_cout_group_7,lo_lo_77}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_77 = {Walloc33bits_77_io_cout_group_21,Walloc33bits_77_io_cout_group_20,
    Walloc33bits_77_io_cout_group_19,Walloc33bits_77_io_cout_group_18,Walloc33bits_77_io_cout_group_17,
    Walloc33bits_77_io_cout_group_16,Walloc33bits_77_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_77 = {Walloc33bits_77_io_cout_group_29,Walloc33bits_77_io_cout_group_28,
    Walloc33bits_77_io_cout_group_27,Walloc33bits_77_io_cout_group_26,Walloc33bits_77_io_cout_group_25,
    Walloc33bits_77_io_cout_group_24,Walloc33bits_77_io_cout_group_23,Walloc33bits_77_io_cout_group_22,hi_lo_77}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_78 = {Walloc33bits_78_io_cout_group_6,Walloc33bits_78_io_cout_group_5,Walloc33bits_78_io_cout_group_4
    ,Walloc33bits_78_io_cout_group_3,Walloc33bits_78_io_cout_group_2,Walloc33bits_78_io_cout_group_1,
    Walloc33bits_78_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_78 = {Walloc33bits_78_io_cout_group_14,Walloc33bits_78_io_cout_group_13,
    Walloc33bits_78_io_cout_group_12,Walloc33bits_78_io_cout_group_11,Walloc33bits_78_io_cout_group_10,
    Walloc33bits_78_io_cout_group_9,Walloc33bits_78_io_cout_group_8,Walloc33bits_78_io_cout_group_7,lo_lo_78}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_78 = {Walloc33bits_78_io_cout_group_21,Walloc33bits_78_io_cout_group_20,
    Walloc33bits_78_io_cout_group_19,Walloc33bits_78_io_cout_group_18,Walloc33bits_78_io_cout_group_17,
    Walloc33bits_78_io_cout_group_16,Walloc33bits_78_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_78 = {Walloc33bits_78_io_cout_group_29,Walloc33bits_78_io_cout_group_28,
    Walloc33bits_78_io_cout_group_27,Walloc33bits_78_io_cout_group_26,Walloc33bits_78_io_cout_group_25,
    Walloc33bits_78_io_cout_group_24,Walloc33bits_78_io_cout_group_23,Walloc33bits_78_io_cout_group_22,hi_lo_78}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_79 = {Walloc33bits_79_io_cout_group_6,Walloc33bits_79_io_cout_group_5,Walloc33bits_79_io_cout_group_4
    ,Walloc33bits_79_io_cout_group_3,Walloc33bits_79_io_cout_group_2,Walloc33bits_79_io_cout_group_1,
    Walloc33bits_79_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_79 = {Walloc33bits_79_io_cout_group_14,Walloc33bits_79_io_cout_group_13,
    Walloc33bits_79_io_cout_group_12,Walloc33bits_79_io_cout_group_11,Walloc33bits_79_io_cout_group_10,
    Walloc33bits_79_io_cout_group_9,Walloc33bits_79_io_cout_group_8,Walloc33bits_79_io_cout_group_7,lo_lo_79}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_79 = {Walloc33bits_79_io_cout_group_21,Walloc33bits_79_io_cout_group_20,
    Walloc33bits_79_io_cout_group_19,Walloc33bits_79_io_cout_group_18,Walloc33bits_79_io_cout_group_17,
    Walloc33bits_79_io_cout_group_16,Walloc33bits_79_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_79 = {Walloc33bits_79_io_cout_group_29,Walloc33bits_79_io_cout_group_28,
    Walloc33bits_79_io_cout_group_27,Walloc33bits_79_io_cout_group_26,Walloc33bits_79_io_cout_group_25,
    Walloc33bits_79_io_cout_group_24,Walloc33bits_79_io_cout_group_23,Walloc33bits_79_io_cout_group_22,hi_lo_79}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_80 = {Walloc33bits_80_io_cout_group_6,Walloc33bits_80_io_cout_group_5,Walloc33bits_80_io_cout_group_4
    ,Walloc33bits_80_io_cout_group_3,Walloc33bits_80_io_cout_group_2,Walloc33bits_80_io_cout_group_1,
    Walloc33bits_80_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_80 = {Walloc33bits_80_io_cout_group_14,Walloc33bits_80_io_cout_group_13,
    Walloc33bits_80_io_cout_group_12,Walloc33bits_80_io_cout_group_11,Walloc33bits_80_io_cout_group_10,
    Walloc33bits_80_io_cout_group_9,Walloc33bits_80_io_cout_group_8,Walloc33bits_80_io_cout_group_7,lo_lo_80}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_80 = {Walloc33bits_80_io_cout_group_21,Walloc33bits_80_io_cout_group_20,
    Walloc33bits_80_io_cout_group_19,Walloc33bits_80_io_cout_group_18,Walloc33bits_80_io_cout_group_17,
    Walloc33bits_80_io_cout_group_16,Walloc33bits_80_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_80 = {Walloc33bits_80_io_cout_group_29,Walloc33bits_80_io_cout_group_28,
    Walloc33bits_80_io_cout_group_27,Walloc33bits_80_io_cout_group_26,Walloc33bits_80_io_cout_group_25,
    Walloc33bits_80_io_cout_group_24,Walloc33bits_80_io_cout_group_23,Walloc33bits_80_io_cout_group_22,hi_lo_80}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_81 = {Walloc33bits_81_io_cout_group_6,Walloc33bits_81_io_cout_group_5,Walloc33bits_81_io_cout_group_4
    ,Walloc33bits_81_io_cout_group_3,Walloc33bits_81_io_cout_group_2,Walloc33bits_81_io_cout_group_1,
    Walloc33bits_81_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_81 = {Walloc33bits_81_io_cout_group_14,Walloc33bits_81_io_cout_group_13,
    Walloc33bits_81_io_cout_group_12,Walloc33bits_81_io_cout_group_11,Walloc33bits_81_io_cout_group_10,
    Walloc33bits_81_io_cout_group_9,Walloc33bits_81_io_cout_group_8,Walloc33bits_81_io_cout_group_7,lo_lo_81}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_81 = {Walloc33bits_81_io_cout_group_21,Walloc33bits_81_io_cout_group_20,
    Walloc33bits_81_io_cout_group_19,Walloc33bits_81_io_cout_group_18,Walloc33bits_81_io_cout_group_17,
    Walloc33bits_81_io_cout_group_16,Walloc33bits_81_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_81 = {Walloc33bits_81_io_cout_group_29,Walloc33bits_81_io_cout_group_28,
    Walloc33bits_81_io_cout_group_27,Walloc33bits_81_io_cout_group_26,Walloc33bits_81_io_cout_group_25,
    Walloc33bits_81_io_cout_group_24,Walloc33bits_81_io_cout_group_23,Walloc33bits_81_io_cout_group_22,hi_lo_81}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_82 = {Walloc33bits_82_io_cout_group_6,Walloc33bits_82_io_cout_group_5,Walloc33bits_82_io_cout_group_4
    ,Walloc33bits_82_io_cout_group_3,Walloc33bits_82_io_cout_group_2,Walloc33bits_82_io_cout_group_1,
    Walloc33bits_82_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_82 = {Walloc33bits_82_io_cout_group_14,Walloc33bits_82_io_cout_group_13,
    Walloc33bits_82_io_cout_group_12,Walloc33bits_82_io_cout_group_11,Walloc33bits_82_io_cout_group_10,
    Walloc33bits_82_io_cout_group_9,Walloc33bits_82_io_cout_group_8,Walloc33bits_82_io_cout_group_7,lo_lo_82}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_82 = {Walloc33bits_82_io_cout_group_21,Walloc33bits_82_io_cout_group_20,
    Walloc33bits_82_io_cout_group_19,Walloc33bits_82_io_cout_group_18,Walloc33bits_82_io_cout_group_17,
    Walloc33bits_82_io_cout_group_16,Walloc33bits_82_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_82 = {Walloc33bits_82_io_cout_group_29,Walloc33bits_82_io_cout_group_28,
    Walloc33bits_82_io_cout_group_27,Walloc33bits_82_io_cout_group_26,Walloc33bits_82_io_cout_group_25,
    Walloc33bits_82_io_cout_group_24,Walloc33bits_82_io_cout_group_23,Walloc33bits_82_io_cout_group_22,hi_lo_82}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_83 = {Walloc33bits_83_io_cout_group_6,Walloc33bits_83_io_cout_group_5,Walloc33bits_83_io_cout_group_4
    ,Walloc33bits_83_io_cout_group_3,Walloc33bits_83_io_cout_group_2,Walloc33bits_83_io_cout_group_1,
    Walloc33bits_83_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_83 = {Walloc33bits_83_io_cout_group_14,Walloc33bits_83_io_cout_group_13,
    Walloc33bits_83_io_cout_group_12,Walloc33bits_83_io_cout_group_11,Walloc33bits_83_io_cout_group_10,
    Walloc33bits_83_io_cout_group_9,Walloc33bits_83_io_cout_group_8,Walloc33bits_83_io_cout_group_7,lo_lo_83}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_83 = {Walloc33bits_83_io_cout_group_21,Walloc33bits_83_io_cout_group_20,
    Walloc33bits_83_io_cout_group_19,Walloc33bits_83_io_cout_group_18,Walloc33bits_83_io_cout_group_17,
    Walloc33bits_83_io_cout_group_16,Walloc33bits_83_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_83 = {Walloc33bits_83_io_cout_group_29,Walloc33bits_83_io_cout_group_28,
    Walloc33bits_83_io_cout_group_27,Walloc33bits_83_io_cout_group_26,Walloc33bits_83_io_cout_group_25,
    Walloc33bits_83_io_cout_group_24,Walloc33bits_83_io_cout_group_23,Walloc33bits_83_io_cout_group_22,hi_lo_83}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_84 = {Walloc33bits_84_io_cout_group_6,Walloc33bits_84_io_cout_group_5,Walloc33bits_84_io_cout_group_4
    ,Walloc33bits_84_io_cout_group_3,Walloc33bits_84_io_cout_group_2,Walloc33bits_84_io_cout_group_1,
    Walloc33bits_84_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_84 = {Walloc33bits_84_io_cout_group_14,Walloc33bits_84_io_cout_group_13,
    Walloc33bits_84_io_cout_group_12,Walloc33bits_84_io_cout_group_11,Walloc33bits_84_io_cout_group_10,
    Walloc33bits_84_io_cout_group_9,Walloc33bits_84_io_cout_group_8,Walloc33bits_84_io_cout_group_7,lo_lo_84}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_84 = {Walloc33bits_84_io_cout_group_21,Walloc33bits_84_io_cout_group_20,
    Walloc33bits_84_io_cout_group_19,Walloc33bits_84_io_cout_group_18,Walloc33bits_84_io_cout_group_17,
    Walloc33bits_84_io_cout_group_16,Walloc33bits_84_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_84 = {Walloc33bits_84_io_cout_group_29,Walloc33bits_84_io_cout_group_28,
    Walloc33bits_84_io_cout_group_27,Walloc33bits_84_io_cout_group_26,Walloc33bits_84_io_cout_group_25,
    Walloc33bits_84_io_cout_group_24,Walloc33bits_84_io_cout_group_23,Walloc33bits_84_io_cout_group_22,hi_lo_84}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_85 = {Walloc33bits_85_io_cout_group_6,Walloc33bits_85_io_cout_group_5,Walloc33bits_85_io_cout_group_4
    ,Walloc33bits_85_io_cout_group_3,Walloc33bits_85_io_cout_group_2,Walloc33bits_85_io_cout_group_1,
    Walloc33bits_85_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_85 = {Walloc33bits_85_io_cout_group_14,Walloc33bits_85_io_cout_group_13,
    Walloc33bits_85_io_cout_group_12,Walloc33bits_85_io_cout_group_11,Walloc33bits_85_io_cout_group_10,
    Walloc33bits_85_io_cout_group_9,Walloc33bits_85_io_cout_group_8,Walloc33bits_85_io_cout_group_7,lo_lo_85}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_85 = {Walloc33bits_85_io_cout_group_21,Walloc33bits_85_io_cout_group_20,
    Walloc33bits_85_io_cout_group_19,Walloc33bits_85_io_cout_group_18,Walloc33bits_85_io_cout_group_17,
    Walloc33bits_85_io_cout_group_16,Walloc33bits_85_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_85 = {Walloc33bits_85_io_cout_group_29,Walloc33bits_85_io_cout_group_28,
    Walloc33bits_85_io_cout_group_27,Walloc33bits_85_io_cout_group_26,Walloc33bits_85_io_cout_group_25,
    Walloc33bits_85_io_cout_group_24,Walloc33bits_85_io_cout_group_23,Walloc33bits_85_io_cout_group_22,hi_lo_85}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_86 = {Walloc33bits_86_io_cout_group_6,Walloc33bits_86_io_cout_group_5,Walloc33bits_86_io_cout_group_4
    ,Walloc33bits_86_io_cout_group_3,Walloc33bits_86_io_cout_group_2,Walloc33bits_86_io_cout_group_1,
    Walloc33bits_86_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_86 = {Walloc33bits_86_io_cout_group_14,Walloc33bits_86_io_cout_group_13,
    Walloc33bits_86_io_cout_group_12,Walloc33bits_86_io_cout_group_11,Walloc33bits_86_io_cout_group_10,
    Walloc33bits_86_io_cout_group_9,Walloc33bits_86_io_cout_group_8,Walloc33bits_86_io_cout_group_7,lo_lo_86}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_86 = {Walloc33bits_86_io_cout_group_21,Walloc33bits_86_io_cout_group_20,
    Walloc33bits_86_io_cout_group_19,Walloc33bits_86_io_cout_group_18,Walloc33bits_86_io_cout_group_17,
    Walloc33bits_86_io_cout_group_16,Walloc33bits_86_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_86 = {Walloc33bits_86_io_cout_group_29,Walloc33bits_86_io_cout_group_28,
    Walloc33bits_86_io_cout_group_27,Walloc33bits_86_io_cout_group_26,Walloc33bits_86_io_cout_group_25,
    Walloc33bits_86_io_cout_group_24,Walloc33bits_86_io_cout_group_23,Walloc33bits_86_io_cout_group_22,hi_lo_86}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_87 = {Walloc33bits_87_io_cout_group_6,Walloc33bits_87_io_cout_group_5,Walloc33bits_87_io_cout_group_4
    ,Walloc33bits_87_io_cout_group_3,Walloc33bits_87_io_cout_group_2,Walloc33bits_87_io_cout_group_1,
    Walloc33bits_87_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_87 = {Walloc33bits_87_io_cout_group_14,Walloc33bits_87_io_cout_group_13,
    Walloc33bits_87_io_cout_group_12,Walloc33bits_87_io_cout_group_11,Walloc33bits_87_io_cout_group_10,
    Walloc33bits_87_io_cout_group_9,Walloc33bits_87_io_cout_group_8,Walloc33bits_87_io_cout_group_7,lo_lo_87}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_87 = {Walloc33bits_87_io_cout_group_21,Walloc33bits_87_io_cout_group_20,
    Walloc33bits_87_io_cout_group_19,Walloc33bits_87_io_cout_group_18,Walloc33bits_87_io_cout_group_17,
    Walloc33bits_87_io_cout_group_16,Walloc33bits_87_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_87 = {Walloc33bits_87_io_cout_group_29,Walloc33bits_87_io_cout_group_28,
    Walloc33bits_87_io_cout_group_27,Walloc33bits_87_io_cout_group_26,Walloc33bits_87_io_cout_group_25,
    Walloc33bits_87_io_cout_group_24,Walloc33bits_87_io_cout_group_23,Walloc33bits_87_io_cout_group_22,hi_lo_87}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_88 = {Walloc33bits_88_io_cout_group_6,Walloc33bits_88_io_cout_group_5,Walloc33bits_88_io_cout_group_4
    ,Walloc33bits_88_io_cout_group_3,Walloc33bits_88_io_cout_group_2,Walloc33bits_88_io_cout_group_1,
    Walloc33bits_88_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_88 = {Walloc33bits_88_io_cout_group_14,Walloc33bits_88_io_cout_group_13,
    Walloc33bits_88_io_cout_group_12,Walloc33bits_88_io_cout_group_11,Walloc33bits_88_io_cout_group_10,
    Walloc33bits_88_io_cout_group_9,Walloc33bits_88_io_cout_group_8,Walloc33bits_88_io_cout_group_7,lo_lo_88}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_88 = {Walloc33bits_88_io_cout_group_21,Walloc33bits_88_io_cout_group_20,
    Walloc33bits_88_io_cout_group_19,Walloc33bits_88_io_cout_group_18,Walloc33bits_88_io_cout_group_17,
    Walloc33bits_88_io_cout_group_16,Walloc33bits_88_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_88 = {Walloc33bits_88_io_cout_group_29,Walloc33bits_88_io_cout_group_28,
    Walloc33bits_88_io_cout_group_27,Walloc33bits_88_io_cout_group_26,Walloc33bits_88_io_cout_group_25,
    Walloc33bits_88_io_cout_group_24,Walloc33bits_88_io_cout_group_23,Walloc33bits_88_io_cout_group_22,hi_lo_88}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_89 = {Walloc33bits_89_io_cout_group_6,Walloc33bits_89_io_cout_group_5,Walloc33bits_89_io_cout_group_4
    ,Walloc33bits_89_io_cout_group_3,Walloc33bits_89_io_cout_group_2,Walloc33bits_89_io_cout_group_1,
    Walloc33bits_89_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_89 = {Walloc33bits_89_io_cout_group_14,Walloc33bits_89_io_cout_group_13,
    Walloc33bits_89_io_cout_group_12,Walloc33bits_89_io_cout_group_11,Walloc33bits_89_io_cout_group_10,
    Walloc33bits_89_io_cout_group_9,Walloc33bits_89_io_cout_group_8,Walloc33bits_89_io_cout_group_7,lo_lo_89}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_89 = {Walloc33bits_89_io_cout_group_21,Walloc33bits_89_io_cout_group_20,
    Walloc33bits_89_io_cout_group_19,Walloc33bits_89_io_cout_group_18,Walloc33bits_89_io_cout_group_17,
    Walloc33bits_89_io_cout_group_16,Walloc33bits_89_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_89 = {Walloc33bits_89_io_cout_group_29,Walloc33bits_89_io_cout_group_28,
    Walloc33bits_89_io_cout_group_27,Walloc33bits_89_io_cout_group_26,Walloc33bits_89_io_cout_group_25,
    Walloc33bits_89_io_cout_group_24,Walloc33bits_89_io_cout_group_23,Walloc33bits_89_io_cout_group_22,hi_lo_89}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_90 = {Walloc33bits_90_io_cout_group_6,Walloc33bits_90_io_cout_group_5,Walloc33bits_90_io_cout_group_4
    ,Walloc33bits_90_io_cout_group_3,Walloc33bits_90_io_cout_group_2,Walloc33bits_90_io_cout_group_1,
    Walloc33bits_90_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_90 = {Walloc33bits_90_io_cout_group_14,Walloc33bits_90_io_cout_group_13,
    Walloc33bits_90_io_cout_group_12,Walloc33bits_90_io_cout_group_11,Walloc33bits_90_io_cout_group_10,
    Walloc33bits_90_io_cout_group_9,Walloc33bits_90_io_cout_group_8,Walloc33bits_90_io_cout_group_7,lo_lo_90}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_90 = {Walloc33bits_90_io_cout_group_21,Walloc33bits_90_io_cout_group_20,
    Walloc33bits_90_io_cout_group_19,Walloc33bits_90_io_cout_group_18,Walloc33bits_90_io_cout_group_17,
    Walloc33bits_90_io_cout_group_16,Walloc33bits_90_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_90 = {Walloc33bits_90_io_cout_group_29,Walloc33bits_90_io_cout_group_28,
    Walloc33bits_90_io_cout_group_27,Walloc33bits_90_io_cout_group_26,Walloc33bits_90_io_cout_group_25,
    Walloc33bits_90_io_cout_group_24,Walloc33bits_90_io_cout_group_23,Walloc33bits_90_io_cout_group_22,hi_lo_90}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_91 = {Walloc33bits_91_io_cout_group_6,Walloc33bits_91_io_cout_group_5,Walloc33bits_91_io_cout_group_4
    ,Walloc33bits_91_io_cout_group_3,Walloc33bits_91_io_cout_group_2,Walloc33bits_91_io_cout_group_1,
    Walloc33bits_91_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_91 = {Walloc33bits_91_io_cout_group_14,Walloc33bits_91_io_cout_group_13,
    Walloc33bits_91_io_cout_group_12,Walloc33bits_91_io_cout_group_11,Walloc33bits_91_io_cout_group_10,
    Walloc33bits_91_io_cout_group_9,Walloc33bits_91_io_cout_group_8,Walloc33bits_91_io_cout_group_7,lo_lo_91}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_91 = {Walloc33bits_91_io_cout_group_21,Walloc33bits_91_io_cout_group_20,
    Walloc33bits_91_io_cout_group_19,Walloc33bits_91_io_cout_group_18,Walloc33bits_91_io_cout_group_17,
    Walloc33bits_91_io_cout_group_16,Walloc33bits_91_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_91 = {Walloc33bits_91_io_cout_group_29,Walloc33bits_91_io_cout_group_28,
    Walloc33bits_91_io_cout_group_27,Walloc33bits_91_io_cout_group_26,Walloc33bits_91_io_cout_group_25,
    Walloc33bits_91_io_cout_group_24,Walloc33bits_91_io_cout_group_23,Walloc33bits_91_io_cout_group_22,hi_lo_91}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_92 = {Walloc33bits_92_io_cout_group_6,Walloc33bits_92_io_cout_group_5,Walloc33bits_92_io_cout_group_4
    ,Walloc33bits_92_io_cout_group_3,Walloc33bits_92_io_cout_group_2,Walloc33bits_92_io_cout_group_1,
    Walloc33bits_92_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_92 = {Walloc33bits_92_io_cout_group_14,Walloc33bits_92_io_cout_group_13,
    Walloc33bits_92_io_cout_group_12,Walloc33bits_92_io_cout_group_11,Walloc33bits_92_io_cout_group_10,
    Walloc33bits_92_io_cout_group_9,Walloc33bits_92_io_cout_group_8,Walloc33bits_92_io_cout_group_7,lo_lo_92}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_92 = {Walloc33bits_92_io_cout_group_21,Walloc33bits_92_io_cout_group_20,
    Walloc33bits_92_io_cout_group_19,Walloc33bits_92_io_cout_group_18,Walloc33bits_92_io_cout_group_17,
    Walloc33bits_92_io_cout_group_16,Walloc33bits_92_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_92 = {Walloc33bits_92_io_cout_group_29,Walloc33bits_92_io_cout_group_28,
    Walloc33bits_92_io_cout_group_27,Walloc33bits_92_io_cout_group_26,Walloc33bits_92_io_cout_group_25,
    Walloc33bits_92_io_cout_group_24,Walloc33bits_92_io_cout_group_23,Walloc33bits_92_io_cout_group_22,hi_lo_92}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_93 = {Walloc33bits_93_io_cout_group_6,Walloc33bits_93_io_cout_group_5,Walloc33bits_93_io_cout_group_4
    ,Walloc33bits_93_io_cout_group_3,Walloc33bits_93_io_cout_group_2,Walloc33bits_93_io_cout_group_1,
    Walloc33bits_93_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_93 = {Walloc33bits_93_io_cout_group_14,Walloc33bits_93_io_cout_group_13,
    Walloc33bits_93_io_cout_group_12,Walloc33bits_93_io_cout_group_11,Walloc33bits_93_io_cout_group_10,
    Walloc33bits_93_io_cout_group_9,Walloc33bits_93_io_cout_group_8,Walloc33bits_93_io_cout_group_7,lo_lo_93}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_93 = {Walloc33bits_93_io_cout_group_21,Walloc33bits_93_io_cout_group_20,
    Walloc33bits_93_io_cout_group_19,Walloc33bits_93_io_cout_group_18,Walloc33bits_93_io_cout_group_17,
    Walloc33bits_93_io_cout_group_16,Walloc33bits_93_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_93 = {Walloc33bits_93_io_cout_group_29,Walloc33bits_93_io_cout_group_28,
    Walloc33bits_93_io_cout_group_27,Walloc33bits_93_io_cout_group_26,Walloc33bits_93_io_cout_group_25,
    Walloc33bits_93_io_cout_group_24,Walloc33bits_93_io_cout_group_23,Walloc33bits_93_io_cout_group_22,hi_lo_93}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_94 = {Walloc33bits_94_io_cout_group_6,Walloc33bits_94_io_cout_group_5,Walloc33bits_94_io_cout_group_4
    ,Walloc33bits_94_io_cout_group_3,Walloc33bits_94_io_cout_group_2,Walloc33bits_94_io_cout_group_1,
    Walloc33bits_94_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_94 = {Walloc33bits_94_io_cout_group_14,Walloc33bits_94_io_cout_group_13,
    Walloc33bits_94_io_cout_group_12,Walloc33bits_94_io_cout_group_11,Walloc33bits_94_io_cout_group_10,
    Walloc33bits_94_io_cout_group_9,Walloc33bits_94_io_cout_group_8,Walloc33bits_94_io_cout_group_7,lo_lo_94}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_94 = {Walloc33bits_94_io_cout_group_21,Walloc33bits_94_io_cout_group_20,
    Walloc33bits_94_io_cout_group_19,Walloc33bits_94_io_cout_group_18,Walloc33bits_94_io_cout_group_17,
    Walloc33bits_94_io_cout_group_16,Walloc33bits_94_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_94 = {Walloc33bits_94_io_cout_group_29,Walloc33bits_94_io_cout_group_28,
    Walloc33bits_94_io_cout_group_27,Walloc33bits_94_io_cout_group_26,Walloc33bits_94_io_cout_group_25,
    Walloc33bits_94_io_cout_group_24,Walloc33bits_94_io_cout_group_23,Walloc33bits_94_io_cout_group_22,hi_lo_94}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_95 = {Walloc33bits_95_io_cout_group_6,Walloc33bits_95_io_cout_group_5,Walloc33bits_95_io_cout_group_4
    ,Walloc33bits_95_io_cout_group_3,Walloc33bits_95_io_cout_group_2,Walloc33bits_95_io_cout_group_1,
    Walloc33bits_95_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_95 = {Walloc33bits_95_io_cout_group_14,Walloc33bits_95_io_cout_group_13,
    Walloc33bits_95_io_cout_group_12,Walloc33bits_95_io_cout_group_11,Walloc33bits_95_io_cout_group_10,
    Walloc33bits_95_io_cout_group_9,Walloc33bits_95_io_cout_group_8,Walloc33bits_95_io_cout_group_7,lo_lo_95}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_95 = {Walloc33bits_95_io_cout_group_21,Walloc33bits_95_io_cout_group_20,
    Walloc33bits_95_io_cout_group_19,Walloc33bits_95_io_cout_group_18,Walloc33bits_95_io_cout_group_17,
    Walloc33bits_95_io_cout_group_16,Walloc33bits_95_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_95 = {Walloc33bits_95_io_cout_group_29,Walloc33bits_95_io_cout_group_28,
    Walloc33bits_95_io_cout_group_27,Walloc33bits_95_io_cout_group_26,Walloc33bits_95_io_cout_group_25,
    Walloc33bits_95_io_cout_group_24,Walloc33bits_95_io_cout_group_23,Walloc33bits_95_io_cout_group_22,hi_lo_95}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_96 = {Walloc33bits_96_io_cout_group_6,Walloc33bits_96_io_cout_group_5,Walloc33bits_96_io_cout_group_4
    ,Walloc33bits_96_io_cout_group_3,Walloc33bits_96_io_cout_group_2,Walloc33bits_96_io_cout_group_1,
    Walloc33bits_96_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_96 = {Walloc33bits_96_io_cout_group_14,Walloc33bits_96_io_cout_group_13,
    Walloc33bits_96_io_cout_group_12,Walloc33bits_96_io_cout_group_11,Walloc33bits_96_io_cout_group_10,
    Walloc33bits_96_io_cout_group_9,Walloc33bits_96_io_cout_group_8,Walloc33bits_96_io_cout_group_7,lo_lo_96}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_96 = {Walloc33bits_96_io_cout_group_21,Walloc33bits_96_io_cout_group_20,
    Walloc33bits_96_io_cout_group_19,Walloc33bits_96_io_cout_group_18,Walloc33bits_96_io_cout_group_17,
    Walloc33bits_96_io_cout_group_16,Walloc33bits_96_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_96 = {Walloc33bits_96_io_cout_group_29,Walloc33bits_96_io_cout_group_28,
    Walloc33bits_96_io_cout_group_27,Walloc33bits_96_io_cout_group_26,Walloc33bits_96_io_cout_group_25,
    Walloc33bits_96_io_cout_group_24,Walloc33bits_96_io_cout_group_23,Walloc33bits_96_io_cout_group_22,hi_lo_96}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_97 = {Walloc33bits_97_io_cout_group_6,Walloc33bits_97_io_cout_group_5,Walloc33bits_97_io_cout_group_4
    ,Walloc33bits_97_io_cout_group_3,Walloc33bits_97_io_cout_group_2,Walloc33bits_97_io_cout_group_1,
    Walloc33bits_97_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_97 = {Walloc33bits_97_io_cout_group_14,Walloc33bits_97_io_cout_group_13,
    Walloc33bits_97_io_cout_group_12,Walloc33bits_97_io_cout_group_11,Walloc33bits_97_io_cout_group_10,
    Walloc33bits_97_io_cout_group_9,Walloc33bits_97_io_cout_group_8,Walloc33bits_97_io_cout_group_7,lo_lo_97}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_97 = {Walloc33bits_97_io_cout_group_21,Walloc33bits_97_io_cout_group_20,
    Walloc33bits_97_io_cout_group_19,Walloc33bits_97_io_cout_group_18,Walloc33bits_97_io_cout_group_17,
    Walloc33bits_97_io_cout_group_16,Walloc33bits_97_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_97 = {Walloc33bits_97_io_cout_group_29,Walloc33bits_97_io_cout_group_28,
    Walloc33bits_97_io_cout_group_27,Walloc33bits_97_io_cout_group_26,Walloc33bits_97_io_cout_group_25,
    Walloc33bits_97_io_cout_group_24,Walloc33bits_97_io_cout_group_23,Walloc33bits_97_io_cout_group_22,hi_lo_97}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_98 = {Walloc33bits_98_io_cout_group_6,Walloc33bits_98_io_cout_group_5,Walloc33bits_98_io_cout_group_4
    ,Walloc33bits_98_io_cout_group_3,Walloc33bits_98_io_cout_group_2,Walloc33bits_98_io_cout_group_1,
    Walloc33bits_98_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_98 = {Walloc33bits_98_io_cout_group_14,Walloc33bits_98_io_cout_group_13,
    Walloc33bits_98_io_cout_group_12,Walloc33bits_98_io_cout_group_11,Walloc33bits_98_io_cout_group_10,
    Walloc33bits_98_io_cout_group_9,Walloc33bits_98_io_cout_group_8,Walloc33bits_98_io_cout_group_7,lo_lo_98}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_98 = {Walloc33bits_98_io_cout_group_21,Walloc33bits_98_io_cout_group_20,
    Walloc33bits_98_io_cout_group_19,Walloc33bits_98_io_cout_group_18,Walloc33bits_98_io_cout_group_17,
    Walloc33bits_98_io_cout_group_16,Walloc33bits_98_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_98 = {Walloc33bits_98_io_cout_group_29,Walloc33bits_98_io_cout_group_28,
    Walloc33bits_98_io_cout_group_27,Walloc33bits_98_io_cout_group_26,Walloc33bits_98_io_cout_group_25,
    Walloc33bits_98_io_cout_group_24,Walloc33bits_98_io_cout_group_23,Walloc33bits_98_io_cout_group_22,hi_lo_98}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_99 = {Walloc33bits_99_io_cout_group_6,Walloc33bits_99_io_cout_group_5,Walloc33bits_99_io_cout_group_4
    ,Walloc33bits_99_io_cout_group_3,Walloc33bits_99_io_cout_group_2,Walloc33bits_99_io_cout_group_1,
    Walloc33bits_99_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_99 = {Walloc33bits_99_io_cout_group_14,Walloc33bits_99_io_cout_group_13,
    Walloc33bits_99_io_cout_group_12,Walloc33bits_99_io_cout_group_11,Walloc33bits_99_io_cout_group_10,
    Walloc33bits_99_io_cout_group_9,Walloc33bits_99_io_cout_group_8,Walloc33bits_99_io_cout_group_7,lo_lo_99}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_99 = {Walloc33bits_99_io_cout_group_21,Walloc33bits_99_io_cout_group_20,
    Walloc33bits_99_io_cout_group_19,Walloc33bits_99_io_cout_group_18,Walloc33bits_99_io_cout_group_17,
    Walloc33bits_99_io_cout_group_16,Walloc33bits_99_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_99 = {Walloc33bits_99_io_cout_group_29,Walloc33bits_99_io_cout_group_28,
    Walloc33bits_99_io_cout_group_27,Walloc33bits_99_io_cout_group_26,Walloc33bits_99_io_cout_group_25,
    Walloc33bits_99_io_cout_group_24,Walloc33bits_99_io_cout_group_23,Walloc33bits_99_io_cout_group_22,hi_lo_99}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_100 = {Walloc33bits_100_io_cout_group_6,Walloc33bits_100_io_cout_group_5,
    Walloc33bits_100_io_cout_group_4,Walloc33bits_100_io_cout_group_3,Walloc33bits_100_io_cout_group_2,
    Walloc33bits_100_io_cout_group_1,Walloc33bits_100_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_100 = {Walloc33bits_100_io_cout_group_14,Walloc33bits_100_io_cout_group_13,
    Walloc33bits_100_io_cout_group_12,Walloc33bits_100_io_cout_group_11,Walloc33bits_100_io_cout_group_10,
    Walloc33bits_100_io_cout_group_9,Walloc33bits_100_io_cout_group_8,Walloc33bits_100_io_cout_group_7,lo_lo_100}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_100 = {Walloc33bits_100_io_cout_group_21,Walloc33bits_100_io_cout_group_20,
    Walloc33bits_100_io_cout_group_19,Walloc33bits_100_io_cout_group_18,Walloc33bits_100_io_cout_group_17,
    Walloc33bits_100_io_cout_group_16,Walloc33bits_100_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_100 = {Walloc33bits_100_io_cout_group_29,Walloc33bits_100_io_cout_group_28,
    Walloc33bits_100_io_cout_group_27,Walloc33bits_100_io_cout_group_26,Walloc33bits_100_io_cout_group_25,
    Walloc33bits_100_io_cout_group_24,Walloc33bits_100_io_cout_group_23,Walloc33bits_100_io_cout_group_22,hi_lo_100}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_101 = {Walloc33bits_101_io_cout_group_6,Walloc33bits_101_io_cout_group_5,
    Walloc33bits_101_io_cout_group_4,Walloc33bits_101_io_cout_group_3,Walloc33bits_101_io_cout_group_2,
    Walloc33bits_101_io_cout_group_1,Walloc33bits_101_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_101 = {Walloc33bits_101_io_cout_group_14,Walloc33bits_101_io_cout_group_13,
    Walloc33bits_101_io_cout_group_12,Walloc33bits_101_io_cout_group_11,Walloc33bits_101_io_cout_group_10,
    Walloc33bits_101_io_cout_group_9,Walloc33bits_101_io_cout_group_8,Walloc33bits_101_io_cout_group_7,lo_lo_101}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_101 = {Walloc33bits_101_io_cout_group_21,Walloc33bits_101_io_cout_group_20,
    Walloc33bits_101_io_cout_group_19,Walloc33bits_101_io_cout_group_18,Walloc33bits_101_io_cout_group_17,
    Walloc33bits_101_io_cout_group_16,Walloc33bits_101_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_101 = {Walloc33bits_101_io_cout_group_29,Walloc33bits_101_io_cout_group_28,
    Walloc33bits_101_io_cout_group_27,Walloc33bits_101_io_cout_group_26,Walloc33bits_101_io_cout_group_25,
    Walloc33bits_101_io_cout_group_24,Walloc33bits_101_io_cout_group_23,Walloc33bits_101_io_cout_group_22,hi_lo_101}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_102 = {Walloc33bits_102_io_cout_group_6,Walloc33bits_102_io_cout_group_5,
    Walloc33bits_102_io_cout_group_4,Walloc33bits_102_io_cout_group_3,Walloc33bits_102_io_cout_group_2,
    Walloc33bits_102_io_cout_group_1,Walloc33bits_102_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_102 = {Walloc33bits_102_io_cout_group_14,Walloc33bits_102_io_cout_group_13,
    Walloc33bits_102_io_cout_group_12,Walloc33bits_102_io_cout_group_11,Walloc33bits_102_io_cout_group_10,
    Walloc33bits_102_io_cout_group_9,Walloc33bits_102_io_cout_group_8,Walloc33bits_102_io_cout_group_7,lo_lo_102}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_102 = {Walloc33bits_102_io_cout_group_21,Walloc33bits_102_io_cout_group_20,
    Walloc33bits_102_io_cout_group_19,Walloc33bits_102_io_cout_group_18,Walloc33bits_102_io_cout_group_17,
    Walloc33bits_102_io_cout_group_16,Walloc33bits_102_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_102 = {Walloc33bits_102_io_cout_group_29,Walloc33bits_102_io_cout_group_28,
    Walloc33bits_102_io_cout_group_27,Walloc33bits_102_io_cout_group_26,Walloc33bits_102_io_cout_group_25,
    Walloc33bits_102_io_cout_group_24,Walloc33bits_102_io_cout_group_23,Walloc33bits_102_io_cout_group_22,hi_lo_102}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_103 = {Walloc33bits_103_io_cout_group_6,Walloc33bits_103_io_cout_group_5,
    Walloc33bits_103_io_cout_group_4,Walloc33bits_103_io_cout_group_3,Walloc33bits_103_io_cout_group_2,
    Walloc33bits_103_io_cout_group_1,Walloc33bits_103_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_103 = {Walloc33bits_103_io_cout_group_14,Walloc33bits_103_io_cout_group_13,
    Walloc33bits_103_io_cout_group_12,Walloc33bits_103_io_cout_group_11,Walloc33bits_103_io_cout_group_10,
    Walloc33bits_103_io_cout_group_9,Walloc33bits_103_io_cout_group_8,Walloc33bits_103_io_cout_group_7,lo_lo_103}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_103 = {Walloc33bits_103_io_cout_group_21,Walloc33bits_103_io_cout_group_20,
    Walloc33bits_103_io_cout_group_19,Walloc33bits_103_io_cout_group_18,Walloc33bits_103_io_cout_group_17,
    Walloc33bits_103_io_cout_group_16,Walloc33bits_103_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_103 = {Walloc33bits_103_io_cout_group_29,Walloc33bits_103_io_cout_group_28,
    Walloc33bits_103_io_cout_group_27,Walloc33bits_103_io_cout_group_26,Walloc33bits_103_io_cout_group_25,
    Walloc33bits_103_io_cout_group_24,Walloc33bits_103_io_cout_group_23,Walloc33bits_103_io_cout_group_22,hi_lo_103}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_104 = {Walloc33bits_104_io_cout_group_6,Walloc33bits_104_io_cout_group_5,
    Walloc33bits_104_io_cout_group_4,Walloc33bits_104_io_cout_group_3,Walloc33bits_104_io_cout_group_2,
    Walloc33bits_104_io_cout_group_1,Walloc33bits_104_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_104 = {Walloc33bits_104_io_cout_group_14,Walloc33bits_104_io_cout_group_13,
    Walloc33bits_104_io_cout_group_12,Walloc33bits_104_io_cout_group_11,Walloc33bits_104_io_cout_group_10,
    Walloc33bits_104_io_cout_group_9,Walloc33bits_104_io_cout_group_8,Walloc33bits_104_io_cout_group_7,lo_lo_104}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_104 = {Walloc33bits_104_io_cout_group_21,Walloc33bits_104_io_cout_group_20,
    Walloc33bits_104_io_cout_group_19,Walloc33bits_104_io_cout_group_18,Walloc33bits_104_io_cout_group_17,
    Walloc33bits_104_io_cout_group_16,Walloc33bits_104_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_104 = {Walloc33bits_104_io_cout_group_29,Walloc33bits_104_io_cout_group_28,
    Walloc33bits_104_io_cout_group_27,Walloc33bits_104_io_cout_group_26,Walloc33bits_104_io_cout_group_25,
    Walloc33bits_104_io_cout_group_24,Walloc33bits_104_io_cout_group_23,Walloc33bits_104_io_cout_group_22,hi_lo_104}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_105 = {Walloc33bits_105_io_cout_group_6,Walloc33bits_105_io_cout_group_5,
    Walloc33bits_105_io_cout_group_4,Walloc33bits_105_io_cout_group_3,Walloc33bits_105_io_cout_group_2,
    Walloc33bits_105_io_cout_group_1,Walloc33bits_105_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_105 = {Walloc33bits_105_io_cout_group_14,Walloc33bits_105_io_cout_group_13,
    Walloc33bits_105_io_cout_group_12,Walloc33bits_105_io_cout_group_11,Walloc33bits_105_io_cout_group_10,
    Walloc33bits_105_io_cout_group_9,Walloc33bits_105_io_cout_group_8,Walloc33bits_105_io_cout_group_7,lo_lo_105}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_105 = {Walloc33bits_105_io_cout_group_21,Walloc33bits_105_io_cout_group_20,
    Walloc33bits_105_io_cout_group_19,Walloc33bits_105_io_cout_group_18,Walloc33bits_105_io_cout_group_17,
    Walloc33bits_105_io_cout_group_16,Walloc33bits_105_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_105 = {Walloc33bits_105_io_cout_group_29,Walloc33bits_105_io_cout_group_28,
    Walloc33bits_105_io_cout_group_27,Walloc33bits_105_io_cout_group_26,Walloc33bits_105_io_cout_group_25,
    Walloc33bits_105_io_cout_group_24,Walloc33bits_105_io_cout_group_23,Walloc33bits_105_io_cout_group_22,hi_lo_105}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_106 = {Walloc33bits_106_io_cout_group_6,Walloc33bits_106_io_cout_group_5,
    Walloc33bits_106_io_cout_group_4,Walloc33bits_106_io_cout_group_3,Walloc33bits_106_io_cout_group_2,
    Walloc33bits_106_io_cout_group_1,Walloc33bits_106_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_106 = {Walloc33bits_106_io_cout_group_14,Walloc33bits_106_io_cout_group_13,
    Walloc33bits_106_io_cout_group_12,Walloc33bits_106_io_cout_group_11,Walloc33bits_106_io_cout_group_10,
    Walloc33bits_106_io_cout_group_9,Walloc33bits_106_io_cout_group_8,Walloc33bits_106_io_cout_group_7,lo_lo_106}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_106 = {Walloc33bits_106_io_cout_group_21,Walloc33bits_106_io_cout_group_20,
    Walloc33bits_106_io_cout_group_19,Walloc33bits_106_io_cout_group_18,Walloc33bits_106_io_cout_group_17,
    Walloc33bits_106_io_cout_group_16,Walloc33bits_106_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_106 = {Walloc33bits_106_io_cout_group_29,Walloc33bits_106_io_cout_group_28,
    Walloc33bits_106_io_cout_group_27,Walloc33bits_106_io_cout_group_26,Walloc33bits_106_io_cout_group_25,
    Walloc33bits_106_io_cout_group_24,Walloc33bits_106_io_cout_group_23,Walloc33bits_106_io_cout_group_22,hi_lo_106}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_107 = {Walloc33bits_107_io_cout_group_6,Walloc33bits_107_io_cout_group_5,
    Walloc33bits_107_io_cout_group_4,Walloc33bits_107_io_cout_group_3,Walloc33bits_107_io_cout_group_2,
    Walloc33bits_107_io_cout_group_1,Walloc33bits_107_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_107 = {Walloc33bits_107_io_cout_group_14,Walloc33bits_107_io_cout_group_13,
    Walloc33bits_107_io_cout_group_12,Walloc33bits_107_io_cout_group_11,Walloc33bits_107_io_cout_group_10,
    Walloc33bits_107_io_cout_group_9,Walloc33bits_107_io_cout_group_8,Walloc33bits_107_io_cout_group_7,lo_lo_107}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_107 = {Walloc33bits_107_io_cout_group_21,Walloc33bits_107_io_cout_group_20,
    Walloc33bits_107_io_cout_group_19,Walloc33bits_107_io_cout_group_18,Walloc33bits_107_io_cout_group_17,
    Walloc33bits_107_io_cout_group_16,Walloc33bits_107_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_107 = {Walloc33bits_107_io_cout_group_29,Walloc33bits_107_io_cout_group_28,
    Walloc33bits_107_io_cout_group_27,Walloc33bits_107_io_cout_group_26,Walloc33bits_107_io_cout_group_25,
    Walloc33bits_107_io_cout_group_24,Walloc33bits_107_io_cout_group_23,Walloc33bits_107_io_cout_group_22,hi_lo_107}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_108 = {Walloc33bits_108_io_cout_group_6,Walloc33bits_108_io_cout_group_5,
    Walloc33bits_108_io_cout_group_4,Walloc33bits_108_io_cout_group_3,Walloc33bits_108_io_cout_group_2,
    Walloc33bits_108_io_cout_group_1,Walloc33bits_108_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_108 = {Walloc33bits_108_io_cout_group_14,Walloc33bits_108_io_cout_group_13,
    Walloc33bits_108_io_cout_group_12,Walloc33bits_108_io_cout_group_11,Walloc33bits_108_io_cout_group_10,
    Walloc33bits_108_io_cout_group_9,Walloc33bits_108_io_cout_group_8,Walloc33bits_108_io_cout_group_7,lo_lo_108}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_108 = {Walloc33bits_108_io_cout_group_21,Walloc33bits_108_io_cout_group_20,
    Walloc33bits_108_io_cout_group_19,Walloc33bits_108_io_cout_group_18,Walloc33bits_108_io_cout_group_17,
    Walloc33bits_108_io_cout_group_16,Walloc33bits_108_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_108 = {Walloc33bits_108_io_cout_group_29,Walloc33bits_108_io_cout_group_28,
    Walloc33bits_108_io_cout_group_27,Walloc33bits_108_io_cout_group_26,Walloc33bits_108_io_cout_group_25,
    Walloc33bits_108_io_cout_group_24,Walloc33bits_108_io_cout_group_23,Walloc33bits_108_io_cout_group_22,hi_lo_108}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_109 = {Walloc33bits_109_io_cout_group_6,Walloc33bits_109_io_cout_group_5,
    Walloc33bits_109_io_cout_group_4,Walloc33bits_109_io_cout_group_3,Walloc33bits_109_io_cout_group_2,
    Walloc33bits_109_io_cout_group_1,Walloc33bits_109_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_109 = {Walloc33bits_109_io_cout_group_14,Walloc33bits_109_io_cout_group_13,
    Walloc33bits_109_io_cout_group_12,Walloc33bits_109_io_cout_group_11,Walloc33bits_109_io_cout_group_10,
    Walloc33bits_109_io_cout_group_9,Walloc33bits_109_io_cout_group_8,Walloc33bits_109_io_cout_group_7,lo_lo_109}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_109 = {Walloc33bits_109_io_cout_group_21,Walloc33bits_109_io_cout_group_20,
    Walloc33bits_109_io_cout_group_19,Walloc33bits_109_io_cout_group_18,Walloc33bits_109_io_cout_group_17,
    Walloc33bits_109_io_cout_group_16,Walloc33bits_109_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_109 = {Walloc33bits_109_io_cout_group_29,Walloc33bits_109_io_cout_group_28,
    Walloc33bits_109_io_cout_group_27,Walloc33bits_109_io_cout_group_26,Walloc33bits_109_io_cout_group_25,
    Walloc33bits_109_io_cout_group_24,Walloc33bits_109_io_cout_group_23,Walloc33bits_109_io_cout_group_22,hi_lo_109}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_110 = {Walloc33bits_110_io_cout_group_6,Walloc33bits_110_io_cout_group_5,
    Walloc33bits_110_io_cout_group_4,Walloc33bits_110_io_cout_group_3,Walloc33bits_110_io_cout_group_2,
    Walloc33bits_110_io_cout_group_1,Walloc33bits_110_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_110 = {Walloc33bits_110_io_cout_group_14,Walloc33bits_110_io_cout_group_13,
    Walloc33bits_110_io_cout_group_12,Walloc33bits_110_io_cout_group_11,Walloc33bits_110_io_cout_group_10,
    Walloc33bits_110_io_cout_group_9,Walloc33bits_110_io_cout_group_8,Walloc33bits_110_io_cout_group_7,lo_lo_110}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_110 = {Walloc33bits_110_io_cout_group_21,Walloc33bits_110_io_cout_group_20,
    Walloc33bits_110_io_cout_group_19,Walloc33bits_110_io_cout_group_18,Walloc33bits_110_io_cout_group_17,
    Walloc33bits_110_io_cout_group_16,Walloc33bits_110_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_110 = {Walloc33bits_110_io_cout_group_29,Walloc33bits_110_io_cout_group_28,
    Walloc33bits_110_io_cout_group_27,Walloc33bits_110_io_cout_group_26,Walloc33bits_110_io_cout_group_25,
    Walloc33bits_110_io_cout_group_24,Walloc33bits_110_io_cout_group_23,Walloc33bits_110_io_cout_group_22,hi_lo_110}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_111 = {Walloc33bits_111_io_cout_group_6,Walloc33bits_111_io_cout_group_5,
    Walloc33bits_111_io_cout_group_4,Walloc33bits_111_io_cout_group_3,Walloc33bits_111_io_cout_group_2,
    Walloc33bits_111_io_cout_group_1,Walloc33bits_111_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_111 = {Walloc33bits_111_io_cout_group_14,Walloc33bits_111_io_cout_group_13,
    Walloc33bits_111_io_cout_group_12,Walloc33bits_111_io_cout_group_11,Walloc33bits_111_io_cout_group_10,
    Walloc33bits_111_io_cout_group_9,Walloc33bits_111_io_cout_group_8,Walloc33bits_111_io_cout_group_7,lo_lo_111}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_111 = {Walloc33bits_111_io_cout_group_21,Walloc33bits_111_io_cout_group_20,
    Walloc33bits_111_io_cout_group_19,Walloc33bits_111_io_cout_group_18,Walloc33bits_111_io_cout_group_17,
    Walloc33bits_111_io_cout_group_16,Walloc33bits_111_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_111 = {Walloc33bits_111_io_cout_group_29,Walloc33bits_111_io_cout_group_28,
    Walloc33bits_111_io_cout_group_27,Walloc33bits_111_io_cout_group_26,Walloc33bits_111_io_cout_group_25,
    Walloc33bits_111_io_cout_group_24,Walloc33bits_111_io_cout_group_23,Walloc33bits_111_io_cout_group_22,hi_lo_111}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_112 = {Walloc33bits_112_io_cout_group_6,Walloc33bits_112_io_cout_group_5,
    Walloc33bits_112_io_cout_group_4,Walloc33bits_112_io_cout_group_3,Walloc33bits_112_io_cout_group_2,
    Walloc33bits_112_io_cout_group_1,Walloc33bits_112_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_112 = {Walloc33bits_112_io_cout_group_14,Walloc33bits_112_io_cout_group_13,
    Walloc33bits_112_io_cout_group_12,Walloc33bits_112_io_cout_group_11,Walloc33bits_112_io_cout_group_10,
    Walloc33bits_112_io_cout_group_9,Walloc33bits_112_io_cout_group_8,Walloc33bits_112_io_cout_group_7,lo_lo_112}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_112 = {Walloc33bits_112_io_cout_group_21,Walloc33bits_112_io_cout_group_20,
    Walloc33bits_112_io_cout_group_19,Walloc33bits_112_io_cout_group_18,Walloc33bits_112_io_cout_group_17,
    Walloc33bits_112_io_cout_group_16,Walloc33bits_112_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_112 = {Walloc33bits_112_io_cout_group_29,Walloc33bits_112_io_cout_group_28,
    Walloc33bits_112_io_cout_group_27,Walloc33bits_112_io_cout_group_26,Walloc33bits_112_io_cout_group_25,
    Walloc33bits_112_io_cout_group_24,Walloc33bits_112_io_cout_group_23,Walloc33bits_112_io_cout_group_22,hi_lo_112}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_113 = {Walloc33bits_113_io_cout_group_6,Walloc33bits_113_io_cout_group_5,
    Walloc33bits_113_io_cout_group_4,Walloc33bits_113_io_cout_group_3,Walloc33bits_113_io_cout_group_2,
    Walloc33bits_113_io_cout_group_1,Walloc33bits_113_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_113 = {Walloc33bits_113_io_cout_group_14,Walloc33bits_113_io_cout_group_13,
    Walloc33bits_113_io_cout_group_12,Walloc33bits_113_io_cout_group_11,Walloc33bits_113_io_cout_group_10,
    Walloc33bits_113_io_cout_group_9,Walloc33bits_113_io_cout_group_8,Walloc33bits_113_io_cout_group_7,lo_lo_113}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_113 = {Walloc33bits_113_io_cout_group_21,Walloc33bits_113_io_cout_group_20,
    Walloc33bits_113_io_cout_group_19,Walloc33bits_113_io_cout_group_18,Walloc33bits_113_io_cout_group_17,
    Walloc33bits_113_io_cout_group_16,Walloc33bits_113_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_113 = {Walloc33bits_113_io_cout_group_29,Walloc33bits_113_io_cout_group_28,
    Walloc33bits_113_io_cout_group_27,Walloc33bits_113_io_cout_group_26,Walloc33bits_113_io_cout_group_25,
    Walloc33bits_113_io_cout_group_24,Walloc33bits_113_io_cout_group_23,Walloc33bits_113_io_cout_group_22,hi_lo_113}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_114 = {Walloc33bits_114_io_cout_group_6,Walloc33bits_114_io_cout_group_5,
    Walloc33bits_114_io_cout_group_4,Walloc33bits_114_io_cout_group_3,Walloc33bits_114_io_cout_group_2,
    Walloc33bits_114_io_cout_group_1,Walloc33bits_114_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_114 = {Walloc33bits_114_io_cout_group_14,Walloc33bits_114_io_cout_group_13,
    Walloc33bits_114_io_cout_group_12,Walloc33bits_114_io_cout_group_11,Walloc33bits_114_io_cout_group_10,
    Walloc33bits_114_io_cout_group_9,Walloc33bits_114_io_cout_group_8,Walloc33bits_114_io_cout_group_7,lo_lo_114}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_114 = {Walloc33bits_114_io_cout_group_21,Walloc33bits_114_io_cout_group_20,
    Walloc33bits_114_io_cout_group_19,Walloc33bits_114_io_cout_group_18,Walloc33bits_114_io_cout_group_17,
    Walloc33bits_114_io_cout_group_16,Walloc33bits_114_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_114 = {Walloc33bits_114_io_cout_group_29,Walloc33bits_114_io_cout_group_28,
    Walloc33bits_114_io_cout_group_27,Walloc33bits_114_io_cout_group_26,Walloc33bits_114_io_cout_group_25,
    Walloc33bits_114_io_cout_group_24,Walloc33bits_114_io_cout_group_23,Walloc33bits_114_io_cout_group_22,hi_lo_114}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_115 = {Walloc33bits_115_io_cout_group_6,Walloc33bits_115_io_cout_group_5,
    Walloc33bits_115_io_cout_group_4,Walloc33bits_115_io_cout_group_3,Walloc33bits_115_io_cout_group_2,
    Walloc33bits_115_io_cout_group_1,Walloc33bits_115_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_115 = {Walloc33bits_115_io_cout_group_14,Walloc33bits_115_io_cout_group_13,
    Walloc33bits_115_io_cout_group_12,Walloc33bits_115_io_cout_group_11,Walloc33bits_115_io_cout_group_10,
    Walloc33bits_115_io_cout_group_9,Walloc33bits_115_io_cout_group_8,Walloc33bits_115_io_cout_group_7,lo_lo_115}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_115 = {Walloc33bits_115_io_cout_group_21,Walloc33bits_115_io_cout_group_20,
    Walloc33bits_115_io_cout_group_19,Walloc33bits_115_io_cout_group_18,Walloc33bits_115_io_cout_group_17,
    Walloc33bits_115_io_cout_group_16,Walloc33bits_115_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_115 = {Walloc33bits_115_io_cout_group_29,Walloc33bits_115_io_cout_group_28,
    Walloc33bits_115_io_cout_group_27,Walloc33bits_115_io_cout_group_26,Walloc33bits_115_io_cout_group_25,
    Walloc33bits_115_io_cout_group_24,Walloc33bits_115_io_cout_group_23,Walloc33bits_115_io_cout_group_22,hi_lo_115}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_116 = {Walloc33bits_116_io_cout_group_6,Walloc33bits_116_io_cout_group_5,
    Walloc33bits_116_io_cout_group_4,Walloc33bits_116_io_cout_group_3,Walloc33bits_116_io_cout_group_2,
    Walloc33bits_116_io_cout_group_1,Walloc33bits_116_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_116 = {Walloc33bits_116_io_cout_group_14,Walloc33bits_116_io_cout_group_13,
    Walloc33bits_116_io_cout_group_12,Walloc33bits_116_io_cout_group_11,Walloc33bits_116_io_cout_group_10,
    Walloc33bits_116_io_cout_group_9,Walloc33bits_116_io_cout_group_8,Walloc33bits_116_io_cout_group_7,lo_lo_116}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_116 = {Walloc33bits_116_io_cout_group_21,Walloc33bits_116_io_cout_group_20,
    Walloc33bits_116_io_cout_group_19,Walloc33bits_116_io_cout_group_18,Walloc33bits_116_io_cout_group_17,
    Walloc33bits_116_io_cout_group_16,Walloc33bits_116_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_116 = {Walloc33bits_116_io_cout_group_29,Walloc33bits_116_io_cout_group_28,
    Walloc33bits_116_io_cout_group_27,Walloc33bits_116_io_cout_group_26,Walloc33bits_116_io_cout_group_25,
    Walloc33bits_116_io_cout_group_24,Walloc33bits_116_io_cout_group_23,Walloc33bits_116_io_cout_group_22,hi_lo_116}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_117 = {Walloc33bits_117_io_cout_group_6,Walloc33bits_117_io_cout_group_5,
    Walloc33bits_117_io_cout_group_4,Walloc33bits_117_io_cout_group_3,Walloc33bits_117_io_cout_group_2,
    Walloc33bits_117_io_cout_group_1,Walloc33bits_117_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_117 = {Walloc33bits_117_io_cout_group_14,Walloc33bits_117_io_cout_group_13,
    Walloc33bits_117_io_cout_group_12,Walloc33bits_117_io_cout_group_11,Walloc33bits_117_io_cout_group_10,
    Walloc33bits_117_io_cout_group_9,Walloc33bits_117_io_cout_group_8,Walloc33bits_117_io_cout_group_7,lo_lo_117}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_117 = {Walloc33bits_117_io_cout_group_21,Walloc33bits_117_io_cout_group_20,
    Walloc33bits_117_io_cout_group_19,Walloc33bits_117_io_cout_group_18,Walloc33bits_117_io_cout_group_17,
    Walloc33bits_117_io_cout_group_16,Walloc33bits_117_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_117 = {Walloc33bits_117_io_cout_group_29,Walloc33bits_117_io_cout_group_28,
    Walloc33bits_117_io_cout_group_27,Walloc33bits_117_io_cout_group_26,Walloc33bits_117_io_cout_group_25,
    Walloc33bits_117_io_cout_group_24,Walloc33bits_117_io_cout_group_23,Walloc33bits_117_io_cout_group_22,hi_lo_117}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_118 = {Walloc33bits_118_io_cout_group_6,Walloc33bits_118_io_cout_group_5,
    Walloc33bits_118_io_cout_group_4,Walloc33bits_118_io_cout_group_3,Walloc33bits_118_io_cout_group_2,
    Walloc33bits_118_io_cout_group_1,Walloc33bits_118_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_118 = {Walloc33bits_118_io_cout_group_14,Walloc33bits_118_io_cout_group_13,
    Walloc33bits_118_io_cout_group_12,Walloc33bits_118_io_cout_group_11,Walloc33bits_118_io_cout_group_10,
    Walloc33bits_118_io_cout_group_9,Walloc33bits_118_io_cout_group_8,Walloc33bits_118_io_cout_group_7,lo_lo_118}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_118 = {Walloc33bits_118_io_cout_group_21,Walloc33bits_118_io_cout_group_20,
    Walloc33bits_118_io_cout_group_19,Walloc33bits_118_io_cout_group_18,Walloc33bits_118_io_cout_group_17,
    Walloc33bits_118_io_cout_group_16,Walloc33bits_118_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_118 = {Walloc33bits_118_io_cout_group_29,Walloc33bits_118_io_cout_group_28,
    Walloc33bits_118_io_cout_group_27,Walloc33bits_118_io_cout_group_26,Walloc33bits_118_io_cout_group_25,
    Walloc33bits_118_io_cout_group_24,Walloc33bits_118_io_cout_group_23,Walloc33bits_118_io_cout_group_22,hi_lo_118}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_119 = {Walloc33bits_119_io_cout_group_6,Walloc33bits_119_io_cout_group_5,
    Walloc33bits_119_io_cout_group_4,Walloc33bits_119_io_cout_group_3,Walloc33bits_119_io_cout_group_2,
    Walloc33bits_119_io_cout_group_1,Walloc33bits_119_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_119 = {Walloc33bits_119_io_cout_group_14,Walloc33bits_119_io_cout_group_13,
    Walloc33bits_119_io_cout_group_12,Walloc33bits_119_io_cout_group_11,Walloc33bits_119_io_cout_group_10,
    Walloc33bits_119_io_cout_group_9,Walloc33bits_119_io_cout_group_8,Walloc33bits_119_io_cout_group_7,lo_lo_119}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_119 = {Walloc33bits_119_io_cout_group_21,Walloc33bits_119_io_cout_group_20,
    Walloc33bits_119_io_cout_group_19,Walloc33bits_119_io_cout_group_18,Walloc33bits_119_io_cout_group_17,
    Walloc33bits_119_io_cout_group_16,Walloc33bits_119_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_119 = {Walloc33bits_119_io_cout_group_29,Walloc33bits_119_io_cout_group_28,
    Walloc33bits_119_io_cout_group_27,Walloc33bits_119_io_cout_group_26,Walloc33bits_119_io_cout_group_25,
    Walloc33bits_119_io_cout_group_24,Walloc33bits_119_io_cout_group_23,Walloc33bits_119_io_cout_group_22,hi_lo_119}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_120 = {Walloc33bits_120_io_cout_group_6,Walloc33bits_120_io_cout_group_5,
    Walloc33bits_120_io_cout_group_4,Walloc33bits_120_io_cout_group_3,Walloc33bits_120_io_cout_group_2,
    Walloc33bits_120_io_cout_group_1,Walloc33bits_120_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_120 = {Walloc33bits_120_io_cout_group_14,Walloc33bits_120_io_cout_group_13,
    Walloc33bits_120_io_cout_group_12,Walloc33bits_120_io_cout_group_11,Walloc33bits_120_io_cout_group_10,
    Walloc33bits_120_io_cout_group_9,Walloc33bits_120_io_cout_group_8,Walloc33bits_120_io_cout_group_7,lo_lo_120}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_120 = {Walloc33bits_120_io_cout_group_21,Walloc33bits_120_io_cout_group_20,
    Walloc33bits_120_io_cout_group_19,Walloc33bits_120_io_cout_group_18,Walloc33bits_120_io_cout_group_17,
    Walloc33bits_120_io_cout_group_16,Walloc33bits_120_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_120 = {Walloc33bits_120_io_cout_group_29,Walloc33bits_120_io_cout_group_28,
    Walloc33bits_120_io_cout_group_27,Walloc33bits_120_io_cout_group_26,Walloc33bits_120_io_cout_group_25,
    Walloc33bits_120_io_cout_group_24,Walloc33bits_120_io_cout_group_23,Walloc33bits_120_io_cout_group_22,hi_lo_120}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_121 = {Walloc33bits_121_io_cout_group_6,Walloc33bits_121_io_cout_group_5,
    Walloc33bits_121_io_cout_group_4,Walloc33bits_121_io_cout_group_3,Walloc33bits_121_io_cout_group_2,
    Walloc33bits_121_io_cout_group_1,Walloc33bits_121_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_121 = {Walloc33bits_121_io_cout_group_14,Walloc33bits_121_io_cout_group_13,
    Walloc33bits_121_io_cout_group_12,Walloc33bits_121_io_cout_group_11,Walloc33bits_121_io_cout_group_10,
    Walloc33bits_121_io_cout_group_9,Walloc33bits_121_io_cout_group_8,Walloc33bits_121_io_cout_group_7,lo_lo_121}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_121 = {Walloc33bits_121_io_cout_group_21,Walloc33bits_121_io_cout_group_20,
    Walloc33bits_121_io_cout_group_19,Walloc33bits_121_io_cout_group_18,Walloc33bits_121_io_cout_group_17,
    Walloc33bits_121_io_cout_group_16,Walloc33bits_121_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_121 = {Walloc33bits_121_io_cout_group_29,Walloc33bits_121_io_cout_group_28,
    Walloc33bits_121_io_cout_group_27,Walloc33bits_121_io_cout_group_26,Walloc33bits_121_io_cout_group_25,
    Walloc33bits_121_io_cout_group_24,Walloc33bits_121_io_cout_group_23,Walloc33bits_121_io_cout_group_22,hi_lo_121}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_122 = {Walloc33bits_122_io_cout_group_6,Walloc33bits_122_io_cout_group_5,
    Walloc33bits_122_io_cout_group_4,Walloc33bits_122_io_cout_group_3,Walloc33bits_122_io_cout_group_2,
    Walloc33bits_122_io_cout_group_1,Walloc33bits_122_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_122 = {Walloc33bits_122_io_cout_group_14,Walloc33bits_122_io_cout_group_13,
    Walloc33bits_122_io_cout_group_12,Walloc33bits_122_io_cout_group_11,Walloc33bits_122_io_cout_group_10,
    Walloc33bits_122_io_cout_group_9,Walloc33bits_122_io_cout_group_8,Walloc33bits_122_io_cout_group_7,lo_lo_122}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_122 = {Walloc33bits_122_io_cout_group_21,Walloc33bits_122_io_cout_group_20,
    Walloc33bits_122_io_cout_group_19,Walloc33bits_122_io_cout_group_18,Walloc33bits_122_io_cout_group_17,
    Walloc33bits_122_io_cout_group_16,Walloc33bits_122_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_122 = {Walloc33bits_122_io_cout_group_29,Walloc33bits_122_io_cout_group_28,
    Walloc33bits_122_io_cout_group_27,Walloc33bits_122_io_cout_group_26,Walloc33bits_122_io_cout_group_25,
    Walloc33bits_122_io_cout_group_24,Walloc33bits_122_io_cout_group_23,Walloc33bits_122_io_cout_group_22,hi_lo_122}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_123 = {Walloc33bits_123_io_cout_group_6,Walloc33bits_123_io_cout_group_5,
    Walloc33bits_123_io_cout_group_4,Walloc33bits_123_io_cout_group_3,Walloc33bits_123_io_cout_group_2,
    Walloc33bits_123_io_cout_group_1,Walloc33bits_123_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_123 = {Walloc33bits_123_io_cout_group_14,Walloc33bits_123_io_cout_group_13,
    Walloc33bits_123_io_cout_group_12,Walloc33bits_123_io_cout_group_11,Walloc33bits_123_io_cout_group_10,
    Walloc33bits_123_io_cout_group_9,Walloc33bits_123_io_cout_group_8,Walloc33bits_123_io_cout_group_7,lo_lo_123}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_123 = {Walloc33bits_123_io_cout_group_21,Walloc33bits_123_io_cout_group_20,
    Walloc33bits_123_io_cout_group_19,Walloc33bits_123_io_cout_group_18,Walloc33bits_123_io_cout_group_17,
    Walloc33bits_123_io_cout_group_16,Walloc33bits_123_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_123 = {Walloc33bits_123_io_cout_group_29,Walloc33bits_123_io_cout_group_28,
    Walloc33bits_123_io_cout_group_27,Walloc33bits_123_io_cout_group_26,Walloc33bits_123_io_cout_group_25,
    Walloc33bits_123_io_cout_group_24,Walloc33bits_123_io_cout_group_23,Walloc33bits_123_io_cout_group_22,hi_lo_123}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_124 = {Walloc33bits_124_io_cout_group_6,Walloc33bits_124_io_cout_group_5,
    Walloc33bits_124_io_cout_group_4,Walloc33bits_124_io_cout_group_3,Walloc33bits_124_io_cout_group_2,
    Walloc33bits_124_io_cout_group_1,Walloc33bits_124_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_124 = {Walloc33bits_124_io_cout_group_14,Walloc33bits_124_io_cout_group_13,
    Walloc33bits_124_io_cout_group_12,Walloc33bits_124_io_cout_group_11,Walloc33bits_124_io_cout_group_10,
    Walloc33bits_124_io_cout_group_9,Walloc33bits_124_io_cout_group_8,Walloc33bits_124_io_cout_group_7,lo_lo_124}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_124 = {Walloc33bits_124_io_cout_group_21,Walloc33bits_124_io_cout_group_20,
    Walloc33bits_124_io_cout_group_19,Walloc33bits_124_io_cout_group_18,Walloc33bits_124_io_cout_group_17,
    Walloc33bits_124_io_cout_group_16,Walloc33bits_124_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_124 = {Walloc33bits_124_io_cout_group_29,Walloc33bits_124_io_cout_group_28,
    Walloc33bits_124_io_cout_group_27,Walloc33bits_124_io_cout_group_26,Walloc33bits_124_io_cout_group_25,
    Walloc33bits_124_io_cout_group_24,Walloc33bits_124_io_cout_group_23,Walloc33bits_124_io_cout_group_22,hi_lo_124}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_125 = {Walloc33bits_125_io_cout_group_6,Walloc33bits_125_io_cout_group_5,
    Walloc33bits_125_io_cout_group_4,Walloc33bits_125_io_cout_group_3,Walloc33bits_125_io_cout_group_2,
    Walloc33bits_125_io_cout_group_1,Walloc33bits_125_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_125 = {Walloc33bits_125_io_cout_group_14,Walloc33bits_125_io_cout_group_13,
    Walloc33bits_125_io_cout_group_12,Walloc33bits_125_io_cout_group_11,Walloc33bits_125_io_cout_group_10,
    Walloc33bits_125_io_cout_group_9,Walloc33bits_125_io_cout_group_8,Walloc33bits_125_io_cout_group_7,lo_lo_125}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_125 = {Walloc33bits_125_io_cout_group_21,Walloc33bits_125_io_cout_group_20,
    Walloc33bits_125_io_cout_group_19,Walloc33bits_125_io_cout_group_18,Walloc33bits_125_io_cout_group_17,
    Walloc33bits_125_io_cout_group_16,Walloc33bits_125_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_125 = {Walloc33bits_125_io_cout_group_29,Walloc33bits_125_io_cout_group_28,
    Walloc33bits_125_io_cout_group_27,Walloc33bits_125_io_cout_group_26,Walloc33bits_125_io_cout_group_25,
    Walloc33bits_125_io_cout_group_24,Walloc33bits_125_io_cout_group_23,Walloc33bits_125_io_cout_group_22,hi_lo_125}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_126 = {Walloc33bits_126_io_cout_group_6,Walloc33bits_126_io_cout_group_5,
    Walloc33bits_126_io_cout_group_4,Walloc33bits_126_io_cout_group_3,Walloc33bits_126_io_cout_group_2,
    Walloc33bits_126_io_cout_group_1,Walloc33bits_126_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_126 = {Walloc33bits_126_io_cout_group_14,Walloc33bits_126_io_cout_group_13,
    Walloc33bits_126_io_cout_group_12,Walloc33bits_126_io_cout_group_11,Walloc33bits_126_io_cout_group_10,
    Walloc33bits_126_io_cout_group_9,Walloc33bits_126_io_cout_group_8,Walloc33bits_126_io_cout_group_7,lo_lo_126}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_126 = {Walloc33bits_126_io_cout_group_21,Walloc33bits_126_io_cout_group_20,
    Walloc33bits_126_io_cout_group_19,Walloc33bits_126_io_cout_group_18,Walloc33bits_126_io_cout_group_17,
    Walloc33bits_126_io_cout_group_16,Walloc33bits_126_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_126 = {Walloc33bits_126_io_cout_group_29,Walloc33bits_126_io_cout_group_28,
    Walloc33bits_126_io_cout_group_27,Walloc33bits_126_io_cout_group_26,Walloc33bits_126_io_cout_group_25,
    Walloc33bits_126_io_cout_group_24,Walloc33bits_126_io_cout_group_23,Walloc33bits_126_io_cout_group_22,hi_lo_126}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_127 = {Walloc33bits_127_io_cout_group_6,Walloc33bits_127_io_cout_group_5,
    Walloc33bits_127_io_cout_group_4,Walloc33bits_127_io_cout_group_3,Walloc33bits_127_io_cout_group_2,
    Walloc33bits_127_io_cout_group_1,Walloc33bits_127_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_127 = {Walloc33bits_127_io_cout_group_14,Walloc33bits_127_io_cout_group_13,
    Walloc33bits_127_io_cout_group_12,Walloc33bits_127_io_cout_group_11,Walloc33bits_127_io_cout_group_10,
    Walloc33bits_127_io_cout_group_9,Walloc33bits_127_io_cout_group_8,Walloc33bits_127_io_cout_group_7,lo_lo_127}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_127 = {Walloc33bits_127_io_cout_group_21,Walloc33bits_127_io_cout_group_20,
    Walloc33bits_127_io_cout_group_19,Walloc33bits_127_io_cout_group_18,Walloc33bits_127_io_cout_group_17,
    Walloc33bits_127_io_cout_group_16,Walloc33bits_127_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_127 = {Walloc33bits_127_io_cout_group_29,Walloc33bits_127_io_cout_group_28,
    Walloc33bits_127_io_cout_group_27,Walloc33bits_127_io_cout_group_26,Walloc33bits_127_io_cout_group_25,
    Walloc33bits_127_io_cout_group_24,Walloc33bits_127_io_cout_group_23,Walloc33bits_127_io_cout_group_22,hi_lo_127}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_128 = {Walloc33bits_128_io_cout_group_6,Walloc33bits_128_io_cout_group_5,
    Walloc33bits_128_io_cout_group_4,Walloc33bits_128_io_cout_group_3,Walloc33bits_128_io_cout_group_2,
    Walloc33bits_128_io_cout_group_1,Walloc33bits_128_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_128 = {Walloc33bits_128_io_cout_group_14,Walloc33bits_128_io_cout_group_13,
    Walloc33bits_128_io_cout_group_12,Walloc33bits_128_io_cout_group_11,Walloc33bits_128_io_cout_group_10,
    Walloc33bits_128_io_cout_group_9,Walloc33bits_128_io_cout_group_8,Walloc33bits_128_io_cout_group_7,lo_lo_128}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_128 = {Walloc33bits_128_io_cout_group_21,Walloc33bits_128_io_cout_group_20,
    Walloc33bits_128_io_cout_group_19,Walloc33bits_128_io_cout_group_18,Walloc33bits_128_io_cout_group_17,
    Walloc33bits_128_io_cout_group_16,Walloc33bits_128_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_128 = {Walloc33bits_128_io_cout_group_29,Walloc33bits_128_io_cout_group_28,
    Walloc33bits_128_io_cout_group_27,Walloc33bits_128_io_cout_group_26,Walloc33bits_128_io_cout_group_25,
    Walloc33bits_128_io_cout_group_24,Walloc33bits_128_io_cout_group_23,Walloc33bits_128_io_cout_group_22,hi_lo_128}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_129 = {Walloc33bits_129_io_cout_group_6,Walloc33bits_129_io_cout_group_5,
    Walloc33bits_129_io_cout_group_4,Walloc33bits_129_io_cout_group_3,Walloc33bits_129_io_cout_group_2,
    Walloc33bits_129_io_cout_group_1,Walloc33bits_129_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_129 = {Walloc33bits_129_io_cout_group_14,Walloc33bits_129_io_cout_group_13,
    Walloc33bits_129_io_cout_group_12,Walloc33bits_129_io_cout_group_11,Walloc33bits_129_io_cout_group_10,
    Walloc33bits_129_io_cout_group_9,Walloc33bits_129_io_cout_group_8,Walloc33bits_129_io_cout_group_7,lo_lo_129}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_129 = {Walloc33bits_129_io_cout_group_21,Walloc33bits_129_io_cout_group_20,
    Walloc33bits_129_io_cout_group_19,Walloc33bits_129_io_cout_group_18,Walloc33bits_129_io_cout_group_17,
    Walloc33bits_129_io_cout_group_16,Walloc33bits_129_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_129 = {Walloc33bits_129_io_cout_group_29,Walloc33bits_129_io_cout_group_28,
    Walloc33bits_129_io_cout_group_27,Walloc33bits_129_io_cout_group_26,Walloc33bits_129_io_cout_group_25,
    Walloc33bits_129_io_cout_group_24,Walloc33bits_129_io_cout_group_23,Walloc33bits_129_io_cout_group_22,hi_lo_129}; // @[WallaceTest.scala 224:37]
  wire [6:0] lo_lo_130 = {Walloc33bits_130_io_cout_group_6,Walloc33bits_130_io_cout_group_5,
    Walloc33bits_130_io_cout_group_4,Walloc33bits_130_io_cout_group_3,Walloc33bits_130_io_cout_group_2,
    Walloc33bits_130_io_cout_group_1,Walloc33bits_130_io_cout_group_0}; // @[WallaceTest.scala 224:37]
  wire [14:0] lo_130 = {Walloc33bits_130_io_cout_group_14,Walloc33bits_130_io_cout_group_13,
    Walloc33bits_130_io_cout_group_12,Walloc33bits_130_io_cout_group_11,Walloc33bits_130_io_cout_group_10,
    Walloc33bits_130_io_cout_group_9,Walloc33bits_130_io_cout_group_8,Walloc33bits_130_io_cout_group_7,lo_lo_130}; // @[WallaceTest.scala 224:37]
  wire [6:0] hi_lo_130 = {Walloc33bits_130_io_cout_group_21,Walloc33bits_130_io_cout_group_20,
    Walloc33bits_130_io_cout_group_19,Walloc33bits_130_io_cout_group_18,Walloc33bits_130_io_cout_group_17,
    Walloc33bits_130_io_cout_group_16,Walloc33bits_130_io_cout_group_15}; // @[WallaceTest.scala 224:37]
  wire [14:0] hi_130 = {Walloc33bits_130_io_cout_group_29,Walloc33bits_130_io_cout_group_28,
    Walloc33bits_130_io_cout_group_27,Walloc33bits_130_io_cout_group_26,Walloc33bits_130_io_cout_group_25,
    Walloc33bits_130_io_cout_group_24,Walloc33bits_130_io_cout_group_23,Walloc33bits_130_io_cout_group_22,hi_lo_130}; // @[WallaceTest.scala 224:37]
  wire  adder_b_0 = switch_io_cout[1]; // @[WallaceTest.scala 229:22]
  wire  adder_a_1 = Walloc33bits_1_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_0 = Walloc33bits_io_cout; // @[WallaceTest.scala 207:21 220:13]
  wire  adder_a_3 = Walloc33bits_3_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_2 = Walloc33bits_2_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_5 = Walloc33bits_5_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_4 = Walloc33bits_4_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_7 = Walloc33bits_7_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_6 = Walloc33bits_6_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_lo_lo_lo_lo = {adder_a_7,adder_a_6,adder_a_5,adder_a_4,adder_a_3,adder_a_2,adder_a_1,adder_a_0}; // @[WallaceTest.scala 231:22]
  wire  adder_a_9 = Walloc33bits_9_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_8 = Walloc33bits_8_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_11 = Walloc33bits_11_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_10 = Walloc33bits_10_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_13 = Walloc33bits_13_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_12 = Walloc33bits_12_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_15 = Walloc33bits_15_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_14 = Walloc33bits_14_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_17 = Walloc33bits_17_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_16 = Walloc33bits_16_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_19 = Walloc33bits_19_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_18 = Walloc33bits_18_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_21 = Walloc33bits_21_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_20 = Walloc33bits_20_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_23 = Walloc33bits_23_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_22 = Walloc33bits_22_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_lo_lo_hi_lo = {adder_a_23,adder_a_22,adder_a_21,adder_a_20,adder_a_19,adder_a_18,adder_a_17,
    adder_a_16}; // @[WallaceTest.scala 231:22]
  wire  adder_a_25 = Walloc33bits_25_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_24 = Walloc33bits_24_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_27 = Walloc33bits_27_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_26 = Walloc33bits_26_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_29 = Walloc33bits_29_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_28 = Walloc33bits_28_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_32 = Walloc33bits_32_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_31 = Walloc33bits_31_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_30 = Walloc33bits_30_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [16:0] result_lo_lo_hi = {adder_a_32,adder_a_31,adder_a_30,adder_a_29,adder_a_28,adder_a_27,adder_a_26,adder_a_25
    ,adder_a_24,result_lo_lo_hi_lo}; // @[WallaceTest.scala 231:22]
  wire [32:0] result_lo_lo = {result_lo_lo_hi,adder_a_15,adder_a_14,adder_a_13,adder_a_12,adder_a_11,adder_a_10,
    adder_a_9,adder_a_8,result_lo_lo_lo_lo}; // @[WallaceTest.scala 231:22]
  wire  adder_a_34 = Walloc33bits_34_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_33 = Walloc33bits_33_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_36 = Walloc33bits_36_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_35 = Walloc33bits_35_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_38 = Walloc33bits_38_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_37 = Walloc33bits_37_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_40 = Walloc33bits_40_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_39 = Walloc33bits_39_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_lo_hi_lo_lo = {adder_a_40,adder_a_39,adder_a_38,adder_a_37,adder_a_36,adder_a_35,adder_a_34,
    adder_a_33}; // @[WallaceTest.scala 231:22]
  wire  adder_a_42 = Walloc33bits_42_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_41 = Walloc33bits_41_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_44 = Walloc33bits_44_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_43 = Walloc33bits_43_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_46 = Walloc33bits_46_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_45 = Walloc33bits_45_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_48 = Walloc33bits_48_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_47 = Walloc33bits_47_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_50 = Walloc33bits_50_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_49 = Walloc33bits_49_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_52 = Walloc33bits_52_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_51 = Walloc33bits_51_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_54 = Walloc33bits_54_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_53 = Walloc33bits_53_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_56 = Walloc33bits_56_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_55 = Walloc33bits_55_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_lo_hi_hi_lo = {adder_a_56,adder_a_55,adder_a_54,adder_a_53,adder_a_52,adder_a_51,adder_a_50,
    adder_a_49}; // @[WallaceTest.scala 231:22]
  wire  adder_a_58 = Walloc33bits_58_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_57 = Walloc33bits_57_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_60 = Walloc33bits_60_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_59 = Walloc33bits_59_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_62 = Walloc33bits_62_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_61 = Walloc33bits_61_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_65 = Walloc33bits_65_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_64 = Walloc33bits_64_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_63 = Walloc33bits_63_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [16:0] result_lo_hi_hi = {adder_a_65,adder_a_64,adder_a_63,adder_a_62,adder_a_61,adder_a_60,adder_a_59,adder_a_58
    ,adder_a_57,result_lo_hi_hi_lo}; // @[WallaceTest.scala 231:22]
  wire [32:0] result_lo_hi = {result_lo_hi_hi,adder_a_48,adder_a_47,adder_a_46,adder_a_45,adder_a_44,adder_a_43,
    adder_a_42,adder_a_41,result_lo_hi_lo_lo}; // @[WallaceTest.scala 231:22]
  wire  adder_a_67 = Walloc33bits_67_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_66 = Walloc33bits_66_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_69 = Walloc33bits_69_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_68 = Walloc33bits_68_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_71 = Walloc33bits_71_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_70 = Walloc33bits_70_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_73 = Walloc33bits_73_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_72 = Walloc33bits_72_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_hi_lo_lo_lo = {adder_a_73,adder_a_72,adder_a_71,adder_a_70,adder_a_69,adder_a_68,adder_a_67,
    adder_a_66}; // @[WallaceTest.scala 231:22]
  wire  adder_a_75 = Walloc33bits_75_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_74 = Walloc33bits_74_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_77 = Walloc33bits_77_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_76 = Walloc33bits_76_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_79 = Walloc33bits_79_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_78 = Walloc33bits_78_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_81 = Walloc33bits_81_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_80 = Walloc33bits_80_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_83 = Walloc33bits_83_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_82 = Walloc33bits_82_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_85 = Walloc33bits_85_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_84 = Walloc33bits_84_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_87 = Walloc33bits_87_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_86 = Walloc33bits_86_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_89 = Walloc33bits_89_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_88 = Walloc33bits_88_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_hi_lo_hi_lo = {adder_a_89,adder_a_88,adder_a_87,adder_a_86,adder_a_85,adder_a_84,adder_a_83,
    adder_a_82}; // @[WallaceTest.scala 231:22]
  wire  adder_a_91 = Walloc33bits_91_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_90 = Walloc33bits_90_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_93 = Walloc33bits_93_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_92 = Walloc33bits_92_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_95 = Walloc33bits_95_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_94 = Walloc33bits_94_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_98 = Walloc33bits_98_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_97 = Walloc33bits_97_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_96 = Walloc33bits_96_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [16:0] result_hi_lo_hi = {adder_a_98,adder_a_97,adder_a_96,adder_a_95,adder_a_94,adder_a_93,adder_a_92,adder_a_91
    ,adder_a_90,result_hi_lo_hi_lo}; // @[WallaceTest.scala 231:22]
  wire [32:0] result_hi_lo = {result_hi_lo_hi,adder_a_81,adder_a_80,adder_a_79,adder_a_78,adder_a_77,adder_a_76,
    adder_a_75,adder_a_74,result_hi_lo_lo_lo}; // @[WallaceTest.scala 231:22]
  wire  adder_a_100 = Walloc33bits_100_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_99 = Walloc33bits_99_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_102 = Walloc33bits_102_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_101 = Walloc33bits_101_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_104 = Walloc33bits_104_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_103 = Walloc33bits_103_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_106 = Walloc33bits_106_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_105 = Walloc33bits_105_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_hi_hi_lo_lo = {adder_a_106,adder_a_105,adder_a_104,adder_a_103,adder_a_102,adder_a_101,adder_a_100,
    adder_a_99}; // @[WallaceTest.scala 231:22]
  wire  adder_a_108 = Walloc33bits_108_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_107 = Walloc33bits_107_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_110 = Walloc33bits_110_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_109 = Walloc33bits_109_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_112 = Walloc33bits_112_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_111 = Walloc33bits_111_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_114 = Walloc33bits_114_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_113 = Walloc33bits_113_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_116 = Walloc33bits_116_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_115 = Walloc33bits_115_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_118 = Walloc33bits_118_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_117 = Walloc33bits_117_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_120 = Walloc33bits_120_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_119 = Walloc33bits_119_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_122 = Walloc33bits_122_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_121 = Walloc33bits_121_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [7:0] result_hi_hi_hi_lo = {adder_a_122,adder_a_121,adder_a_120,adder_a_119,adder_a_118,adder_a_117,adder_a_116,
    adder_a_115}; // @[WallaceTest.scala 231:22]
  wire  adder_a_124 = Walloc33bits_124_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_123 = Walloc33bits_123_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_126 = Walloc33bits_126_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_125 = Walloc33bits_125_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_128 = Walloc33bits_128_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_127 = Walloc33bits_127_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_131 = Walloc33bits_131_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_130 = Walloc33bits_130_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire  adder_a_129 = Walloc33bits_129_io_cout; // @[WallaceTest.scala 207:21 225:15]
  wire [16:0] result_hi_hi_hi = {adder_a_131,adder_a_130,adder_a_129,adder_a_128,adder_a_127,adder_a_126,adder_a_125,
    adder_a_124,adder_a_123,result_hi_hi_hi_lo}; // @[WallaceTest.scala 231:22]
  wire [32:0] result_hi_hi = {result_hi_hi_hi,adder_a_114,adder_a_113,adder_a_112,adder_a_111,adder_a_110,adder_a_109,
    adder_a_108,adder_a_107,result_hi_hi_lo_lo}; // @[WallaceTest.scala 231:22]
  wire [131:0] _result_T = {result_hi_hi,result_hi_lo,result_lo_hi,result_lo_lo}; // @[WallaceTest.scala 231:22]
  wire  adder_b_1 = Walloc33bits_io_s; // @[WallaceTest.scala 208:21 221:13]
  wire  adder_b_3 = Walloc33bits_2_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_2 = Walloc33bits_1_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_5 = Walloc33bits_4_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_4 = Walloc33bits_3_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_7 = Walloc33bits_6_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_6 = Walloc33bits_5_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_lo_lo_lo_lo_1 = {adder_b_7,adder_b_6,adder_b_5,adder_b_4,adder_b_3,adder_b_2,adder_b_1,adder_b_0}; // @[WallaceTest.scala 231:39]
  wire  adder_b_9 = Walloc33bits_8_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_8 = Walloc33bits_7_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_11 = Walloc33bits_10_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_10 = Walloc33bits_9_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_13 = Walloc33bits_12_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_12 = Walloc33bits_11_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_15 = Walloc33bits_14_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_14 = Walloc33bits_13_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_17 = Walloc33bits_16_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_16 = Walloc33bits_15_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_19 = Walloc33bits_18_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_18 = Walloc33bits_17_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_21 = Walloc33bits_20_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_20 = Walloc33bits_19_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_23 = Walloc33bits_22_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_22 = Walloc33bits_21_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_lo_lo_hi_lo_1 = {adder_b_23,adder_b_22,adder_b_21,adder_b_20,adder_b_19,adder_b_18,adder_b_17,
    adder_b_16}; // @[WallaceTest.scala 231:39]
  wire  adder_b_25 = Walloc33bits_24_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_24 = Walloc33bits_23_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_27 = Walloc33bits_26_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_26 = Walloc33bits_25_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_29 = Walloc33bits_28_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_28 = Walloc33bits_27_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_32 = Walloc33bits_31_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_31 = Walloc33bits_30_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_30 = Walloc33bits_29_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [16:0] result_lo_lo_hi_1 = {adder_b_32,adder_b_31,adder_b_30,adder_b_29,adder_b_28,adder_b_27,adder_b_26,
    adder_b_25,adder_b_24,result_lo_lo_hi_lo_1}; // @[WallaceTest.scala 231:39]
  wire [32:0] result_lo_lo_1 = {result_lo_lo_hi_1,adder_b_15,adder_b_14,adder_b_13,adder_b_12,adder_b_11,adder_b_10,
    adder_b_9,adder_b_8,result_lo_lo_lo_lo_1}; // @[WallaceTest.scala 231:39]
  wire  adder_b_34 = Walloc33bits_33_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_33 = Walloc33bits_32_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_36 = Walloc33bits_35_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_35 = Walloc33bits_34_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_38 = Walloc33bits_37_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_37 = Walloc33bits_36_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_40 = Walloc33bits_39_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_39 = Walloc33bits_38_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_lo_hi_lo_lo_1 = {adder_b_40,adder_b_39,adder_b_38,adder_b_37,adder_b_36,adder_b_35,adder_b_34,
    adder_b_33}; // @[WallaceTest.scala 231:39]
  wire  adder_b_42 = Walloc33bits_41_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_41 = Walloc33bits_40_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_44 = Walloc33bits_43_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_43 = Walloc33bits_42_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_46 = Walloc33bits_45_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_45 = Walloc33bits_44_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_48 = Walloc33bits_47_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_47 = Walloc33bits_46_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_50 = Walloc33bits_49_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_49 = Walloc33bits_48_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_52 = Walloc33bits_51_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_51 = Walloc33bits_50_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_54 = Walloc33bits_53_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_53 = Walloc33bits_52_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_56 = Walloc33bits_55_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_55 = Walloc33bits_54_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_lo_hi_hi_lo_1 = {adder_b_56,adder_b_55,adder_b_54,adder_b_53,adder_b_52,adder_b_51,adder_b_50,
    adder_b_49}; // @[WallaceTest.scala 231:39]
  wire  adder_b_58 = Walloc33bits_57_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_57 = Walloc33bits_56_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_60 = Walloc33bits_59_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_59 = Walloc33bits_58_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_62 = Walloc33bits_61_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_61 = Walloc33bits_60_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_65 = Walloc33bits_64_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_64 = Walloc33bits_63_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_63 = Walloc33bits_62_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [16:0] result_lo_hi_hi_1 = {adder_b_65,adder_b_64,adder_b_63,adder_b_62,adder_b_61,adder_b_60,adder_b_59,
    adder_b_58,adder_b_57,result_lo_hi_hi_lo_1}; // @[WallaceTest.scala 231:39]
  wire [32:0] result_lo_hi_1 = {result_lo_hi_hi_1,adder_b_48,adder_b_47,adder_b_46,adder_b_45,adder_b_44,adder_b_43,
    adder_b_42,adder_b_41,result_lo_hi_lo_lo_1}; // @[WallaceTest.scala 231:39]
  wire  adder_b_67 = Walloc33bits_66_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_66 = Walloc33bits_65_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_69 = Walloc33bits_68_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_68 = Walloc33bits_67_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_71 = Walloc33bits_70_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_70 = Walloc33bits_69_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_73 = Walloc33bits_72_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_72 = Walloc33bits_71_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_hi_lo_lo_lo_1 = {adder_b_73,adder_b_72,adder_b_71,adder_b_70,adder_b_69,adder_b_68,adder_b_67,
    adder_b_66}; // @[WallaceTest.scala 231:39]
  wire  adder_b_75 = Walloc33bits_74_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_74 = Walloc33bits_73_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_77 = Walloc33bits_76_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_76 = Walloc33bits_75_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_79 = Walloc33bits_78_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_78 = Walloc33bits_77_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_81 = Walloc33bits_80_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_80 = Walloc33bits_79_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_83 = Walloc33bits_82_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_82 = Walloc33bits_81_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_85 = Walloc33bits_84_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_84 = Walloc33bits_83_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_87 = Walloc33bits_86_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_86 = Walloc33bits_85_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_89 = Walloc33bits_88_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_88 = Walloc33bits_87_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_hi_lo_hi_lo_1 = {adder_b_89,adder_b_88,adder_b_87,adder_b_86,adder_b_85,adder_b_84,adder_b_83,
    adder_b_82}; // @[WallaceTest.scala 231:39]
  wire  adder_b_91 = Walloc33bits_90_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_90 = Walloc33bits_89_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_93 = Walloc33bits_92_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_92 = Walloc33bits_91_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_95 = Walloc33bits_94_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_94 = Walloc33bits_93_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_98 = Walloc33bits_97_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_97 = Walloc33bits_96_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_96 = Walloc33bits_95_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [16:0] result_hi_lo_hi_1 = {adder_b_98,adder_b_97,adder_b_96,adder_b_95,adder_b_94,adder_b_93,adder_b_92,
    adder_b_91,adder_b_90,result_hi_lo_hi_lo_1}; // @[WallaceTest.scala 231:39]
  wire [32:0] result_hi_lo_1 = {result_hi_lo_hi_1,adder_b_81,adder_b_80,adder_b_79,adder_b_78,adder_b_77,adder_b_76,
    adder_b_75,adder_b_74,result_hi_lo_lo_lo_1}; // @[WallaceTest.scala 231:39]
  wire  adder_b_100 = Walloc33bits_99_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_99 = Walloc33bits_98_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_102 = Walloc33bits_101_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_101 = Walloc33bits_100_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_104 = Walloc33bits_103_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_103 = Walloc33bits_102_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_106 = Walloc33bits_105_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_105 = Walloc33bits_104_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_hi_hi_lo_lo_1 = {adder_b_106,adder_b_105,adder_b_104,adder_b_103,adder_b_102,adder_b_101,adder_b_100
    ,adder_b_99}; // @[WallaceTest.scala 231:39]
  wire  adder_b_108 = Walloc33bits_107_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_107 = Walloc33bits_106_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_110 = Walloc33bits_109_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_109 = Walloc33bits_108_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_112 = Walloc33bits_111_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_111 = Walloc33bits_110_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_115 = Walloc33bits_114_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_114 = Walloc33bits_113_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_113 = Walloc33bits_112_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [16:0] result_hi_hi_lo_1 = {adder_b_115,adder_b_114,adder_b_113,adder_b_112,adder_b_111,adder_b_110,adder_b_109,
    adder_b_108,adder_b_107,result_hi_hi_lo_lo_1}; // @[WallaceTest.scala 231:39]
  wire  adder_b_117 = Walloc33bits_116_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_116 = Walloc33bits_115_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_119 = Walloc33bits_118_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_118 = Walloc33bits_117_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_121 = Walloc33bits_120_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_120 = Walloc33bits_119_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_123 = Walloc33bits_122_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_122 = Walloc33bits_121_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [7:0] result_hi_hi_hi_lo_1 = {adder_b_123,adder_b_122,adder_b_121,adder_b_120,adder_b_119,adder_b_118,adder_b_117
    ,adder_b_116}; // @[WallaceTest.scala 231:39]
  wire  adder_b_125 = Walloc33bits_124_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_124 = Walloc33bits_123_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_127 = Walloc33bits_126_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_126 = Walloc33bits_125_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_129 = Walloc33bits_128_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_128 = Walloc33bits_127_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_132 = Walloc33bits_131_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_131 = Walloc33bits_130_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire  adder_b_130 = Walloc33bits_129_io_s; // @[WallaceTest.scala 208:21 226:17]
  wire [16:0] result_hi_hi_hi_1 = {adder_b_132,adder_b_131,adder_b_130,adder_b_129,adder_b_128,adder_b_127,adder_b_126,
    adder_b_125,adder_b_124,result_hi_hi_hi_lo_1}; // @[WallaceTest.scala 231:39]
  wire [132:0] _result_T_1 = {result_hi_hi_hi_1,result_hi_hi_lo_1,result_hi_lo_1,result_lo_hi_1,result_lo_lo_1}; // @[WallaceTest.scala 231:39]
  wire [132:0] _GEN_0 = {{1'd0}, _result_T}; // @[WallaceTest.scala 231:29]
  wire [132:0] _result_T_4 = _GEN_0 + _result_T_1; // @[WallaceTest.scala 231:29]
  wire [132:0] _GEN_1 = {{132'd0}, switch_io_cout[0]}; // @[WallaceTest.scala 231:53]
  wire [132:0] _result_T_7 = _result_T_4 + _GEN_1; // @[WallaceTest.scala 231:53]
  wire [127:0] result = _result_T_7[127:0]; // @[WallaceTest.scala 231:66]
  gen_p gen_p ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_io_src),
    .io_x(gen_p_io_x),
    .io_p(gen_p_io_p),
    .io_c(gen_p_io_c)
  );
  gen_p gen_p_1 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_1_io_src),
    .io_x(gen_p_1_io_x),
    .io_p(gen_p_1_io_p),
    .io_c(gen_p_1_io_c)
  );
  gen_p gen_p_2 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_2_io_src),
    .io_x(gen_p_2_io_x),
    .io_p(gen_p_2_io_p),
    .io_c(gen_p_2_io_c)
  );
  gen_p gen_p_3 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_3_io_src),
    .io_x(gen_p_3_io_x),
    .io_p(gen_p_3_io_p),
    .io_c(gen_p_3_io_c)
  );
  gen_p gen_p_4 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_4_io_src),
    .io_x(gen_p_4_io_x),
    .io_p(gen_p_4_io_p),
    .io_c(gen_p_4_io_c)
  );
  gen_p gen_p_5 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_5_io_src),
    .io_x(gen_p_5_io_x),
    .io_p(gen_p_5_io_p),
    .io_c(gen_p_5_io_c)
  );
  gen_p gen_p_6 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_6_io_src),
    .io_x(gen_p_6_io_x),
    .io_p(gen_p_6_io_p),
    .io_c(gen_p_6_io_c)
  );
  gen_p gen_p_7 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_7_io_src),
    .io_x(gen_p_7_io_x),
    .io_p(gen_p_7_io_p),
    .io_c(gen_p_7_io_c)
  );
  gen_p gen_p_8 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_8_io_src),
    .io_x(gen_p_8_io_x),
    .io_p(gen_p_8_io_p),
    .io_c(gen_p_8_io_c)
  );
  gen_p gen_p_9 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_9_io_src),
    .io_x(gen_p_9_io_x),
    .io_p(gen_p_9_io_p),
    .io_c(gen_p_9_io_c)
  );
  gen_p gen_p_10 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_10_io_src),
    .io_x(gen_p_10_io_x),
    .io_p(gen_p_10_io_p),
    .io_c(gen_p_10_io_c)
  );
  gen_p gen_p_11 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_11_io_src),
    .io_x(gen_p_11_io_x),
    .io_p(gen_p_11_io_p),
    .io_c(gen_p_11_io_c)
  );
  gen_p gen_p_12 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_12_io_src),
    .io_x(gen_p_12_io_x),
    .io_p(gen_p_12_io_p),
    .io_c(gen_p_12_io_c)
  );
  gen_p gen_p_13 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_13_io_src),
    .io_x(gen_p_13_io_x),
    .io_p(gen_p_13_io_p),
    .io_c(gen_p_13_io_c)
  );
  gen_p gen_p_14 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_14_io_src),
    .io_x(gen_p_14_io_x),
    .io_p(gen_p_14_io_p),
    .io_c(gen_p_14_io_c)
  );
  gen_p gen_p_15 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_15_io_src),
    .io_x(gen_p_15_io_x),
    .io_p(gen_p_15_io_p),
    .io_c(gen_p_15_io_c)
  );
  gen_p gen_p_16 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_16_io_src),
    .io_x(gen_p_16_io_x),
    .io_p(gen_p_16_io_p),
    .io_c(gen_p_16_io_c)
  );
  gen_p gen_p_17 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_17_io_src),
    .io_x(gen_p_17_io_x),
    .io_p(gen_p_17_io_p),
    .io_c(gen_p_17_io_c)
  );
  gen_p gen_p_18 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_18_io_src),
    .io_x(gen_p_18_io_x),
    .io_p(gen_p_18_io_p),
    .io_c(gen_p_18_io_c)
  );
  gen_p gen_p_19 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_19_io_src),
    .io_x(gen_p_19_io_x),
    .io_p(gen_p_19_io_p),
    .io_c(gen_p_19_io_c)
  );
  gen_p gen_p_20 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_20_io_src),
    .io_x(gen_p_20_io_x),
    .io_p(gen_p_20_io_p),
    .io_c(gen_p_20_io_c)
  );
  gen_p gen_p_21 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_21_io_src),
    .io_x(gen_p_21_io_x),
    .io_p(gen_p_21_io_p),
    .io_c(gen_p_21_io_c)
  );
  gen_p gen_p_22 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_22_io_src),
    .io_x(gen_p_22_io_x),
    .io_p(gen_p_22_io_p),
    .io_c(gen_p_22_io_c)
  );
  gen_p gen_p_23 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_23_io_src),
    .io_x(gen_p_23_io_x),
    .io_p(gen_p_23_io_p),
    .io_c(gen_p_23_io_c)
  );
  gen_p gen_p_24 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_24_io_src),
    .io_x(gen_p_24_io_x),
    .io_p(gen_p_24_io_p),
    .io_c(gen_p_24_io_c)
  );
  gen_p gen_p_25 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_25_io_src),
    .io_x(gen_p_25_io_x),
    .io_p(gen_p_25_io_p),
    .io_c(gen_p_25_io_c)
  );
  gen_p gen_p_26 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_26_io_src),
    .io_x(gen_p_26_io_x),
    .io_p(gen_p_26_io_p),
    .io_c(gen_p_26_io_c)
  );
  gen_p gen_p_27 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_27_io_src),
    .io_x(gen_p_27_io_x),
    .io_p(gen_p_27_io_p),
    .io_c(gen_p_27_io_c)
  );
  gen_p gen_p_28 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_28_io_src),
    .io_x(gen_p_28_io_x),
    .io_p(gen_p_28_io_p),
    .io_c(gen_p_28_io_c)
  );
  gen_p gen_p_29 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_29_io_src),
    .io_x(gen_p_29_io_x),
    .io_p(gen_p_29_io_p),
    .io_c(gen_p_29_io_c)
  );
  gen_p gen_p_30 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_30_io_src),
    .io_x(gen_p_30_io_x),
    .io_p(gen_p_30_io_p),
    .io_c(gen_p_30_io_c)
  );
  gen_p gen_p_31 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_31_io_src),
    .io_x(gen_p_31_io_x),
    .io_p(gen_p_31_io_p),
    .io_c(gen_p_31_io_c)
  );
  gen_p gen_p_32 ( // @[WallaceTest.scala 204:30]
    .io_src(gen_p_32_io_src),
    .io_x(gen_p_32_io_x),
    .io_p(gen_p_32_io_p),
    .io_c(gen_p_32_io_c)
  );
  switch switch ( // @[WallaceTest.scala 205:16]
    .clock(switch_clock),
    .reset(switch_reset),
    .io_in_0(switch_io_in_0),
    .io_in_1(switch_io_in_1),
    .io_in_2(switch_io_in_2),
    .io_in_3(switch_io_in_3),
    .io_in_4(switch_io_in_4),
    .io_in_5(switch_io_in_5),
    .io_in_6(switch_io_in_6),
    .io_in_7(switch_io_in_7),
    .io_in_8(switch_io_in_8),
    .io_in_9(switch_io_in_9),
    .io_in_10(switch_io_in_10),
    .io_in_11(switch_io_in_11),
    .io_in_12(switch_io_in_12),
    .io_in_13(switch_io_in_13),
    .io_in_14(switch_io_in_14),
    .io_in_15(switch_io_in_15),
    .io_in_16(switch_io_in_16),
    .io_in_17(switch_io_in_17),
    .io_in_18(switch_io_in_18),
    .io_in_19(switch_io_in_19),
    .io_in_20(switch_io_in_20),
    .io_in_21(switch_io_in_21),
    .io_in_22(switch_io_in_22),
    .io_in_23(switch_io_in_23),
    .io_in_24(switch_io_in_24),
    .io_in_25(switch_io_in_25),
    .io_in_26(switch_io_in_26),
    .io_in_27(switch_io_in_27),
    .io_in_28(switch_io_in_28),
    .io_in_29(switch_io_in_29),
    .io_in_30(switch_io_in_30),
    .io_in_31(switch_io_in_31),
    .io_in_32(switch_io_in_32),
    .io_out_0(switch_io_out_0),
    .io_out_1(switch_io_out_1),
    .io_out_2(switch_io_out_2),
    .io_out_3(switch_io_out_3),
    .io_out_4(switch_io_out_4),
    .io_out_5(switch_io_out_5),
    .io_out_6(switch_io_out_6),
    .io_out_7(switch_io_out_7),
    .io_out_8(switch_io_out_8),
    .io_out_9(switch_io_out_9),
    .io_out_10(switch_io_out_10),
    .io_out_11(switch_io_out_11),
    .io_out_12(switch_io_out_12),
    .io_out_13(switch_io_out_13),
    .io_out_14(switch_io_out_14),
    .io_out_15(switch_io_out_15),
    .io_out_16(switch_io_out_16),
    .io_out_17(switch_io_out_17),
    .io_out_18(switch_io_out_18),
    .io_out_19(switch_io_out_19),
    .io_out_20(switch_io_out_20),
    .io_out_21(switch_io_out_21),
    .io_out_22(switch_io_out_22),
    .io_out_23(switch_io_out_23),
    .io_out_24(switch_io_out_24),
    .io_out_25(switch_io_out_25),
    .io_out_26(switch_io_out_26),
    .io_out_27(switch_io_out_27),
    .io_out_28(switch_io_out_28),
    .io_out_29(switch_io_out_29),
    .io_out_30(switch_io_out_30),
    .io_out_31(switch_io_out_31),
    .io_out_32(switch_io_out_32),
    .io_out_33(switch_io_out_33),
    .io_out_34(switch_io_out_34),
    .io_out_35(switch_io_out_35),
    .io_out_36(switch_io_out_36),
    .io_out_37(switch_io_out_37),
    .io_out_38(switch_io_out_38),
    .io_out_39(switch_io_out_39),
    .io_out_40(switch_io_out_40),
    .io_out_41(switch_io_out_41),
    .io_out_42(switch_io_out_42),
    .io_out_43(switch_io_out_43),
    .io_out_44(switch_io_out_44),
    .io_out_45(switch_io_out_45),
    .io_out_46(switch_io_out_46),
    .io_out_47(switch_io_out_47),
    .io_out_48(switch_io_out_48),
    .io_out_49(switch_io_out_49),
    .io_out_50(switch_io_out_50),
    .io_out_51(switch_io_out_51),
    .io_out_52(switch_io_out_52),
    .io_out_53(switch_io_out_53),
    .io_out_54(switch_io_out_54),
    .io_out_55(switch_io_out_55),
    .io_out_56(switch_io_out_56),
    .io_out_57(switch_io_out_57),
    .io_out_58(switch_io_out_58),
    .io_out_59(switch_io_out_59),
    .io_out_60(switch_io_out_60),
    .io_out_61(switch_io_out_61),
    .io_out_62(switch_io_out_62),
    .io_out_63(switch_io_out_63),
    .io_out_64(switch_io_out_64),
    .io_out_65(switch_io_out_65),
    .io_out_66(switch_io_out_66),
    .io_out_67(switch_io_out_67),
    .io_out_68(switch_io_out_68),
    .io_out_69(switch_io_out_69),
    .io_out_70(switch_io_out_70),
    .io_out_71(switch_io_out_71),
    .io_out_72(switch_io_out_72),
    .io_out_73(switch_io_out_73),
    .io_out_74(switch_io_out_74),
    .io_out_75(switch_io_out_75),
    .io_out_76(switch_io_out_76),
    .io_out_77(switch_io_out_77),
    .io_out_78(switch_io_out_78),
    .io_out_79(switch_io_out_79),
    .io_out_80(switch_io_out_80),
    .io_out_81(switch_io_out_81),
    .io_out_82(switch_io_out_82),
    .io_out_83(switch_io_out_83),
    .io_out_84(switch_io_out_84),
    .io_out_85(switch_io_out_85),
    .io_out_86(switch_io_out_86),
    .io_out_87(switch_io_out_87),
    .io_out_88(switch_io_out_88),
    .io_out_89(switch_io_out_89),
    .io_out_90(switch_io_out_90),
    .io_out_91(switch_io_out_91),
    .io_out_92(switch_io_out_92),
    .io_out_93(switch_io_out_93),
    .io_out_94(switch_io_out_94),
    .io_out_95(switch_io_out_95),
    .io_out_96(switch_io_out_96),
    .io_out_97(switch_io_out_97),
    .io_out_98(switch_io_out_98),
    .io_out_99(switch_io_out_99),
    .io_out_100(switch_io_out_100),
    .io_out_101(switch_io_out_101),
    .io_out_102(switch_io_out_102),
    .io_out_103(switch_io_out_103),
    .io_out_104(switch_io_out_104),
    .io_out_105(switch_io_out_105),
    .io_out_106(switch_io_out_106),
    .io_out_107(switch_io_out_107),
    .io_out_108(switch_io_out_108),
    .io_out_109(switch_io_out_109),
    .io_out_110(switch_io_out_110),
    .io_out_111(switch_io_out_111),
    .io_out_112(switch_io_out_112),
    .io_out_113(switch_io_out_113),
    .io_out_114(switch_io_out_114),
    .io_out_115(switch_io_out_115),
    .io_out_116(switch_io_out_116),
    .io_out_117(switch_io_out_117),
    .io_out_118(switch_io_out_118),
    .io_out_119(switch_io_out_119),
    .io_out_120(switch_io_out_120),
    .io_out_121(switch_io_out_121),
    .io_out_122(switch_io_out_122),
    .io_out_123(switch_io_out_123),
    .io_out_124(switch_io_out_124),
    .io_out_125(switch_io_out_125),
    .io_out_126(switch_io_out_126),
    .io_out_127(switch_io_out_127),
    .io_out_128(switch_io_out_128),
    .io_out_129(switch_io_out_129),
    .io_out_130(switch_io_out_130),
    .io_out_131(switch_io_out_131),
    .io_cin_0(switch_io_cin_0),
    .io_cin_1(switch_io_cin_1),
    .io_cin_2(switch_io_cin_2),
    .io_cin_3(switch_io_cin_3),
    .io_cin_4(switch_io_cin_4),
    .io_cin_5(switch_io_cin_5),
    .io_cin_6(switch_io_cin_6),
    .io_cin_7(switch_io_cin_7),
    .io_cin_8(switch_io_cin_8),
    .io_cin_9(switch_io_cin_9),
    .io_cin_10(switch_io_cin_10),
    .io_cin_11(switch_io_cin_11),
    .io_cin_12(switch_io_cin_12),
    .io_cin_13(switch_io_cin_13),
    .io_cin_14(switch_io_cin_14),
    .io_cin_15(switch_io_cin_15),
    .io_cin_16(switch_io_cin_16),
    .io_cin_17(switch_io_cin_17),
    .io_cin_18(switch_io_cin_18),
    .io_cin_19(switch_io_cin_19),
    .io_cin_20(switch_io_cin_20),
    .io_cin_21(switch_io_cin_21),
    .io_cin_22(switch_io_cin_22),
    .io_cin_23(switch_io_cin_23),
    .io_cin_24(switch_io_cin_24),
    .io_cin_25(switch_io_cin_25),
    .io_cin_26(switch_io_cin_26),
    .io_cin_27(switch_io_cin_27),
    .io_cin_28(switch_io_cin_28),
    .io_cin_29(switch_io_cin_29),
    .io_cin_30(switch_io_cin_30),
    .io_cin_31(switch_io_cin_31),
    .io_cin_32(switch_io_cin_32),
    .io_cout(switch_io_cout)
  );
  Walloc33bits Walloc33bits ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_io_src_in),
    .io_cin(Walloc33bits_io_cin),
    .io_cout_group_0(Walloc33bits_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_io_cout_group_29),
    .io_cout(Walloc33bits_io_cout),
    .io_s(Walloc33bits_io_s)
  );
  Walloc33bits Walloc33bits_1 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_1_io_src_in),
    .io_cin(Walloc33bits_1_io_cin),
    .io_cout_group_0(Walloc33bits_1_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_1_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_1_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_1_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_1_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_1_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_1_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_1_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_1_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_1_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_1_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_1_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_1_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_1_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_1_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_1_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_1_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_1_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_1_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_1_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_1_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_1_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_1_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_1_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_1_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_1_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_1_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_1_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_1_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_1_io_cout_group_29),
    .io_cout(Walloc33bits_1_io_cout),
    .io_s(Walloc33bits_1_io_s)
  );
  Walloc33bits Walloc33bits_2 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_2_io_src_in),
    .io_cin(Walloc33bits_2_io_cin),
    .io_cout_group_0(Walloc33bits_2_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_2_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_2_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_2_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_2_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_2_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_2_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_2_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_2_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_2_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_2_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_2_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_2_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_2_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_2_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_2_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_2_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_2_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_2_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_2_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_2_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_2_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_2_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_2_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_2_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_2_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_2_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_2_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_2_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_2_io_cout_group_29),
    .io_cout(Walloc33bits_2_io_cout),
    .io_s(Walloc33bits_2_io_s)
  );
  Walloc33bits Walloc33bits_3 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_3_io_src_in),
    .io_cin(Walloc33bits_3_io_cin),
    .io_cout_group_0(Walloc33bits_3_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_3_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_3_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_3_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_3_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_3_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_3_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_3_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_3_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_3_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_3_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_3_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_3_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_3_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_3_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_3_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_3_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_3_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_3_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_3_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_3_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_3_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_3_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_3_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_3_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_3_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_3_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_3_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_3_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_3_io_cout_group_29),
    .io_cout(Walloc33bits_3_io_cout),
    .io_s(Walloc33bits_3_io_s)
  );
  Walloc33bits Walloc33bits_4 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_4_io_src_in),
    .io_cin(Walloc33bits_4_io_cin),
    .io_cout_group_0(Walloc33bits_4_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_4_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_4_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_4_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_4_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_4_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_4_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_4_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_4_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_4_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_4_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_4_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_4_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_4_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_4_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_4_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_4_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_4_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_4_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_4_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_4_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_4_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_4_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_4_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_4_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_4_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_4_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_4_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_4_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_4_io_cout_group_29),
    .io_cout(Walloc33bits_4_io_cout),
    .io_s(Walloc33bits_4_io_s)
  );
  Walloc33bits Walloc33bits_5 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_5_io_src_in),
    .io_cin(Walloc33bits_5_io_cin),
    .io_cout_group_0(Walloc33bits_5_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_5_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_5_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_5_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_5_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_5_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_5_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_5_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_5_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_5_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_5_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_5_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_5_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_5_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_5_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_5_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_5_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_5_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_5_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_5_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_5_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_5_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_5_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_5_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_5_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_5_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_5_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_5_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_5_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_5_io_cout_group_29),
    .io_cout(Walloc33bits_5_io_cout),
    .io_s(Walloc33bits_5_io_s)
  );
  Walloc33bits Walloc33bits_6 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_6_io_src_in),
    .io_cin(Walloc33bits_6_io_cin),
    .io_cout_group_0(Walloc33bits_6_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_6_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_6_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_6_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_6_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_6_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_6_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_6_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_6_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_6_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_6_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_6_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_6_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_6_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_6_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_6_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_6_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_6_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_6_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_6_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_6_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_6_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_6_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_6_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_6_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_6_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_6_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_6_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_6_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_6_io_cout_group_29),
    .io_cout(Walloc33bits_6_io_cout),
    .io_s(Walloc33bits_6_io_s)
  );
  Walloc33bits Walloc33bits_7 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_7_io_src_in),
    .io_cin(Walloc33bits_7_io_cin),
    .io_cout_group_0(Walloc33bits_7_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_7_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_7_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_7_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_7_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_7_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_7_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_7_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_7_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_7_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_7_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_7_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_7_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_7_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_7_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_7_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_7_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_7_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_7_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_7_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_7_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_7_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_7_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_7_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_7_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_7_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_7_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_7_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_7_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_7_io_cout_group_29),
    .io_cout(Walloc33bits_7_io_cout),
    .io_s(Walloc33bits_7_io_s)
  );
  Walloc33bits Walloc33bits_8 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_8_io_src_in),
    .io_cin(Walloc33bits_8_io_cin),
    .io_cout_group_0(Walloc33bits_8_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_8_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_8_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_8_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_8_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_8_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_8_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_8_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_8_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_8_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_8_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_8_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_8_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_8_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_8_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_8_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_8_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_8_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_8_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_8_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_8_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_8_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_8_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_8_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_8_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_8_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_8_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_8_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_8_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_8_io_cout_group_29),
    .io_cout(Walloc33bits_8_io_cout),
    .io_s(Walloc33bits_8_io_s)
  );
  Walloc33bits Walloc33bits_9 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_9_io_src_in),
    .io_cin(Walloc33bits_9_io_cin),
    .io_cout_group_0(Walloc33bits_9_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_9_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_9_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_9_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_9_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_9_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_9_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_9_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_9_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_9_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_9_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_9_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_9_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_9_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_9_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_9_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_9_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_9_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_9_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_9_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_9_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_9_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_9_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_9_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_9_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_9_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_9_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_9_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_9_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_9_io_cout_group_29),
    .io_cout(Walloc33bits_9_io_cout),
    .io_s(Walloc33bits_9_io_s)
  );
  Walloc33bits Walloc33bits_10 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_10_io_src_in),
    .io_cin(Walloc33bits_10_io_cin),
    .io_cout_group_0(Walloc33bits_10_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_10_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_10_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_10_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_10_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_10_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_10_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_10_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_10_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_10_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_10_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_10_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_10_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_10_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_10_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_10_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_10_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_10_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_10_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_10_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_10_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_10_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_10_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_10_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_10_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_10_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_10_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_10_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_10_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_10_io_cout_group_29),
    .io_cout(Walloc33bits_10_io_cout),
    .io_s(Walloc33bits_10_io_s)
  );
  Walloc33bits Walloc33bits_11 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_11_io_src_in),
    .io_cin(Walloc33bits_11_io_cin),
    .io_cout_group_0(Walloc33bits_11_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_11_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_11_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_11_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_11_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_11_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_11_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_11_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_11_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_11_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_11_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_11_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_11_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_11_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_11_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_11_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_11_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_11_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_11_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_11_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_11_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_11_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_11_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_11_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_11_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_11_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_11_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_11_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_11_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_11_io_cout_group_29),
    .io_cout(Walloc33bits_11_io_cout),
    .io_s(Walloc33bits_11_io_s)
  );
  Walloc33bits Walloc33bits_12 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_12_io_src_in),
    .io_cin(Walloc33bits_12_io_cin),
    .io_cout_group_0(Walloc33bits_12_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_12_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_12_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_12_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_12_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_12_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_12_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_12_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_12_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_12_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_12_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_12_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_12_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_12_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_12_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_12_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_12_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_12_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_12_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_12_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_12_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_12_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_12_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_12_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_12_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_12_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_12_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_12_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_12_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_12_io_cout_group_29),
    .io_cout(Walloc33bits_12_io_cout),
    .io_s(Walloc33bits_12_io_s)
  );
  Walloc33bits Walloc33bits_13 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_13_io_src_in),
    .io_cin(Walloc33bits_13_io_cin),
    .io_cout_group_0(Walloc33bits_13_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_13_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_13_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_13_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_13_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_13_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_13_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_13_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_13_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_13_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_13_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_13_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_13_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_13_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_13_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_13_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_13_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_13_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_13_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_13_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_13_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_13_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_13_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_13_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_13_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_13_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_13_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_13_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_13_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_13_io_cout_group_29),
    .io_cout(Walloc33bits_13_io_cout),
    .io_s(Walloc33bits_13_io_s)
  );
  Walloc33bits Walloc33bits_14 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_14_io_src_in),
    .io_cin(Walloc33bits_14_io_cin),
    .io_cout_group_0(Walloc33bits_14_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_14_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_14_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_14_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_14_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_14_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_14_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_14_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_14_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_14_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_14_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_14_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_14_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_14_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_14_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_14_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_14_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_14_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_14_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_14_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_14_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_14_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_14_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_14_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_14_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_14_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_14_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_14_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_14_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_14_io_cout_group_29),
    .io_cout(Walloc33bits_14_io_cout),
    .io_s(Walloc33bits_14_io_s)
  );
  Walloc33bits Walloc33bits_15 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_15_io_src_in),
    .io_cin(Walloc33bits_15_io_cin),
    .io_cout_group_0(Walloc33bits_15_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_15_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_15_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_15_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_15_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_15_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_15_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_15_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_15_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_15_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_15_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_15_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_15_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_15_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_15_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_15_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_15_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_15_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_15_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_15_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_15_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_15_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_15_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_15_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_15_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_15_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_15_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_15_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_15_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_15_io_cout_group_29),
    .io_cout(Walloc33bits_15_io_cout),
    .io_s(Walloc33bits_15_io_s)
  );
  Walloc33bits Walloc33bits_16 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_16_io_src_in),
    .io_cin(Walloc33bits_16_io_cin),
    .io_cout_group_0(Walloc33bits_16_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_16_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_16_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_16_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_16_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_16_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_16_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_16_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_16_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_16_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_16_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_16_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_16_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_16_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_16_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_16_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_16_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_16_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_16_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_16_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_16_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_16_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_16_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_16_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_16_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_16_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_16_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_16_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_16_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_16_io_cout_group_29),
    .io_cout(Walloc33bits_16_io_cout),
    .io_s(Walloc33bits_16_io_s)
  );
  Walloc33bits Walloc33bits_17 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_17_io_src_in),
    .io_cin(Walloc33bits_17_io_cin),
    .io_cout_group_0(Walloc33bits_17_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_17_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_17_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_17_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_17_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_17_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_17_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_17_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_17_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_17_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_17_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_17_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_17_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_17_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_17_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_17_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_17_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_17_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_17_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_17_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_17_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_17_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_17_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_17_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_17_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_17_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_17_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_17_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_17_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_17_io_cout_group_29),
    .io_cout(Walloc33bits_17_io_cout),
    .io_s(Walloc33bits_17_io_s)
  );
  Walloc33bits Walloc33bits_18 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_18_io_src_in),
    .io_cin(Walloc33bits_18_io_cin),
    .io_cout_group_0(Walloc33bits_18_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_18_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_18_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_18_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_18_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_18_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_18_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_18_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_18_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_18_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_18_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_18_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_18_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_18_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_18_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_18_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_18_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_18_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_18_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_18_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_18_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_18_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_18_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_18_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_18_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_18_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_18_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_18_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_18_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_18_io_cout_group_29),
    .io_cout(Walloc33bits_18_io_cout),
    .io_s(Walloc33bits_18_io_s)
  );
  Walloc33bits Walloc33bits_19 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_19_io_src_in),
    .io_cin(Walloc33bits_19_io_cin),
    .io_cout_group_0(Walloc33bits_19_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_19_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_19_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_19_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_19_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_19_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_19_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_19_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_19_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_19_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_19_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_19_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_19_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_19_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_19_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_19_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_19_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_19_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_19_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_19_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_19_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_19_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_19_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_19_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_19_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_19_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_19_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_19_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_19_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_19_io_cout_group_29),
    .io_cout(Walloc33bits_19_io_cout),
    .io_s(Walloc33bits_19_io_s)
  );
  Walloc33bits Walloc33bits_20 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_20_io_src_in),
    .io_cin(Walloc33bits_20_io_cin),
    .io_cout_group_0(Walloc33bits_20_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_20_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_20_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_20_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_20_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_20_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_20_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_20_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_20_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_20_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_20_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_20_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_20_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_20_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_20_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_20_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_20_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_20_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_20_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_20_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_20_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_20_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_20_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_20_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_20_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_20_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_20_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_20_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_20_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_20_io_cout_group_29),
    .io_cout(Walloc33bits_20_io_cout),
    .io_s(Walloc33bits_20_io_s)
  );
  Walloc33bits Walloc33bits_21 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_21_io_src_in),
    .io_cin(Walloc33bits_21_io_cin),
    .io_cout_group_0(Walloc33bits_21_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_21_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_21_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_21_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_21_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_21_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_21_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_21_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_21_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_21_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_21_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_21_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_21_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_21_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_21_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_21_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_21_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_21_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_21_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_21_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_21_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_21_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_21_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_21_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_21_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_21_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_21_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_21_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_21_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_21_io_cout_group_29),
    .io_cout(Walloc33bits_21_io_cout),
    .io_s(Walloc33bits_21_io_s)
  );
  Walloc33bits Walloc33bits_22 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_22_io_src_in),
    .io_cin(Walloc33bits_22_io_cin),
    .io_cout_group_0(Walloc33bits_22_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_22_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_22_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_22_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_22_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_22_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_22_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_22_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_22_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_22_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_22_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_22_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_22_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_22_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_22_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_22_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_22_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_22_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_22_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_22_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_22_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_22_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_22_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_22_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_22_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_22_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_22_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_22_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_22_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_22_io_cout_group_29),
    .io_cout(Walloc33bits_22_io_cout),
    .io_s(Walloc33bits_22_io_s)
  );
  Walloc33bits Walloc33bits_23 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_23_io_src_in),
    .io_cin(Walloc33bits_23_io_cin),
    .io_cout_group_0(Walloc33bits_23_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_23_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_23_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_23_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_23_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_23_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_23_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_23_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_23_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_23_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_23_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_23_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_23_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_23_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_23_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_23_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_23_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_23_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_23_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_23_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_23_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_23_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_23_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_23_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_23_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_23_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_23_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_23_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_23_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_23_io_cout_group_29),
    .io_cout(Walloc33bits_23_io_cout),
    .io_s(Walloc33bits_23_io_s)
  );
  Walloc33bits Walloc33bits_24 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_24_io_src_in),
    .io_cin(Walloc33bits_24_io_cin),
    .io_cout_group_0(Walloc33bits_24_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_24_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_24_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_24_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_24_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_24_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_24_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_24_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_24_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_24_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_24_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_24_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_24_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_24_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_24_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_24_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_24_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_24_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_24_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_24_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_24_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_24_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_24_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_24_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_24_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_24_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_24_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_24_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_24_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_24_io_cout_group_29),
    .io_cout(Walloc33bits_24_io_cout),
    .io_s(Walloc33bits_24_io_s)
  );
  Walloc33bits Walloc33bits_25 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_25_io_src_in),
    .io_cin(Walloc33bits_25_io_cin),
    .io_cout_group_0(Walloc33bits_25_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_25_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_25_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_25_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_25_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_25_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_25_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_25_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_25_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_25_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_25_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_25_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_25_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_25_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_25_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_25_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_25_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_25_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_25_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_25_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_25_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_25_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_25_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_25_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_25_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_25_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_25_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_25_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_25_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_25_io_cout_group_29),
    .io_cout(Walloc33bits_25_io_cout),
    .io_s(Walloc33bits_25_io_s)
  );
  Walloc33bits Walloc33bits_26 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_26_io_src_in),
    .io_cin(Walloc33bits_26_io_cin),
    .io_cout_group_0(Walloc33bits_26_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_26_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_26_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_26_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_26_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_26_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_26_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_26_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_26_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_26_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_26_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_26_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_26_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_26_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_26_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_26_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_26_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_26_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_26_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_26_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_26_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_26_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_26_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_26_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_26_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_26_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_26_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_26_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_26_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_26_io_cout_group_29),
    .io_cout(Walloc33bits_26_io_cout),
    .io_s(Walloc33bits_26_io_s)
  );
  Walloc33bits Walloc33bits_27 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_27_io_src_in),
    .io_cin(Walloc33bits_27_io_cin),
    .io_cout_group_0(Walloc33bits_27_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_27_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_27_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_27_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_27_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_27_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_27_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_27_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_27_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_27_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_27_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_27_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_27_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_27_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_27_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_27_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_27_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_27_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_27_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_27_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_27_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_27_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_27_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_27_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_27_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_27_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_27_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_27_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_27_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_27_io_cout_group_29),
    .io_cout(Walloc33bits_27_io_cout),
    .io_s(Walloc33bits_27_io_s)
  );
  Walloc33bits Walloc33bits_28 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_28_io_src_in),
    .io_cin(Walloc33bits_28_io_cin),
    .io_cout_group_0(Walloc33bits_28_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_28_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_28_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_28_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_28_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_28_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_28_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_28_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_28_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_28_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_28_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_28_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_28_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_28_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_28_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_28_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_28_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_28_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_28_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_28_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_28_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_28_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_28_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_28_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_28_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_28_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_28_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_28_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_28_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_28_io_cout_group_29),
    .io_cout(Walloc33bits_28_io_cout),
    .io_s(Walloc33bits_28_io_s)
  );
  Walloc33bits Walloc33bits_29 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_29_io_src_in),
    .io_cin(Walloc33bits_29_io_cin),
    .io_cout_group_0(Walloc33bits_29_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_29_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_29_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_29_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_29_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_29_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_29_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_29_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_29_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_29_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_29_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_29_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_29_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_29_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_29_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_29_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_29_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_29_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_29_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_29_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_29_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_29_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_29_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_29_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_29_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_29_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_29_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_29_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_29_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_29_io_cout_group_29),
    .io_cout(Walloc33bits_29_io_cout),
    .io_s(Walloc33bits_29_io_s)
  );
  Walloc33bits Walloc33bits_30 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_30_io_src_in),
    .io_cin(Walloc33bits_30_io_cin),
    .io_cout_group_0(Walloc33bits_30_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_30_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_30_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_30_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_30_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_30_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_30_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_30_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_30_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_30_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_30_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_30_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_30_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_30_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_30_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_30_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_30_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_30_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_30_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_30_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_30_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_30_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_30_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_30_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_30_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_30_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_30_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_30_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_30_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_30_io_cout_group_29),
    .io_cout(Walloc33bits_30_io_cout),
    .io_s(Walloc33bits_30_io_s)
  );
  Walloc33bits Walloc33bits_31 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_31_io_src_in),
    .io_cin(Walloc33bits_31_io_cin),
    .io_cout_group_0(Walloc33bits_31_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_31_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_31_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_31_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_31_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_31_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_31_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_31_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_31_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_31_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_31_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_31_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_31_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_31_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_31_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_31_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_31_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_31_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_31_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_31_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_31_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_31_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_31_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_31_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_31_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_31_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_31_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_31_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_31_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_31_io_cout_group_29),
    .io_cout(Walloc33bits_31_io_cout),
    .io_s(Walloc33bits_31_io_s)
  );
  Walloc33bits Walloc33bits_32 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_32_io_src_in),
    .io_cin(Walloc33bits_32_io_cin),
    .io_cout_group_0(Walloc33bits_32_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_32_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_32_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_32_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_32_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_32_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_32_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_32_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_32_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_32_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_32_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_32_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_32_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_32_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_32_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_32_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_32_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_32_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_32_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_32_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_32_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_32_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_32_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_32_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_32_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_32_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_32_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_32_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_32_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_32_io_cout_group_29),
    .io_cout(Walloc33bits_32_io_cout),
    .io_s(Walloc33bits_32_io_s)
  );
  Walloc33bits Walloc33bits_33 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_33_io_src_in),
    .io_cin(Walloc33bits_33_io_cin),
    .io_cout_group_0(Walloc33bits_33_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_33_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_33_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_33_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_33_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_33_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_33_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_33_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_33_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_33_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_33_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_33_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_33_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_33_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_33_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_33_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_33_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_33_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_33_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_33_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_33_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_33_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_33_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_33_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_33_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_33_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_33_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_33_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_33_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_33_io_cout_group_29),
    .io_cout(Walloc33bits_33_io_cout),
    .io_s(Walloc33bits_33_io_s)
  );
  Walloc33bits Walloc33bits_34 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_34_io_src_in),
    .io_cin(Walloc33bits_34_io_cin),
    .io_cout_group_0(Walloc33bits_34_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_34_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_34_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_34_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_34_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_34_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_34_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_34_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_34_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_34_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_34_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_34_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_34_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_34_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_34_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_34_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_34_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_34_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_34_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_34_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_34_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_34_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_34_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_34_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_34_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_34_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_34_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_34_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_34_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_34_io_cout_group_29),
    .io_cout(Walloc33bits_34_io_cout),
    .io_s(Walloc33bits_34_io_s)
  );
  Walloc33bits Walloc33bits_35 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_35_io_src_in),
    .io_cin(Walloc33bits_35_io_cin),
    .io_cout_group_0(Walloc33bits_35_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_35_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_35_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_35_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_35_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_35_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_35_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_35_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_35_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_35_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_35_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_35_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_35_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_35_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_35_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_35_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_35_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_35_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_35_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_35_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_35_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_35_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_35_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_35_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_35_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_35_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_35_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_35_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_35_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_35_io_cout_group_29),
    .io_cout(Walloc33bits_35_io_cout),
    .io_s(Walloc33bits_35_io_s)
  );
  Walloc33bits Walloc33bits_36 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_36_io_src_in),
    .io_cin(Walloc33bits_36_io_cin),
    .io_cout_group_0(Walloc33bits_36_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_36_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_36_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_36_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_36_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_36_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_36_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_36_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_36_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_36_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_36_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_36_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_36_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_36_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_36_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_36_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_36_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_36_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_36_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_36_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_36_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_36_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_36_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_36_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_36_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_36_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_36_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_36_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_36_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_36_io_cout_group_29),
    .io_cout(Walloc33bits_36_io_cout),
    .io_s(Walloc33bits_36_io_s)
  );
  Walloc33bits Walloc33bits_37 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_37_io_src_in),
    .io_cin(Walloc33bits_37_io_cin),
    .io_cout_group_0(Walloc33bits_37_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_37_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_37_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_37_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_37_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_37_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_37_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_37_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_37_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_37_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_37_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_37_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_37_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_37_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_37_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_37_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_37_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_37_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_37_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_37_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_37_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_37_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_37_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_37_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_37_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_37_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_37_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_37_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_37_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_37_io_cout_group_29),
    .io_cout(Walloc33bits_37_io_cout),
    .io_s(Walloc33bits_37_io_s)
  );
  Walloc33bits Walloc33bits_38 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_38_io_src_in),
    .io_cin(Walloc33bits_38_io_cin),
    .io_cout_group_0(Walloc33bits_38_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_38_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_38_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_38_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_38_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_38_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_38_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_38_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_38_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_38_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_38_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_38_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_38_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_38_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_38_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_38_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_38_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_38_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_38_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_38_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_38_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_38_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_38_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_38_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_38_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_38_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_38_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_38_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_38_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_38_io_cout_group_29),
    .io_cout(Walloc33bits_38_io_cout),
    .io_s(Walloc33bits_38_io_s)
  );
  Walloc33bits Walloc33bits_39 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_39_io_src_in),
    .io_cin(Walloc33bits_39_io_cin),
    .io_cout_group_0(Walloc33bits_39_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_39_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_39_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_39_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_39_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_39_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_39_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_39_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_39_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_39_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_39_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_39_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_39_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_39_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_39_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_39_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_39_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_39_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_39_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_39_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_39_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_39_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_39_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_39_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_39_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_39_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_39_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_39_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_39_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_39_io_cout_group_29),
    .io_cout(Walloc33bits_39_io_cout),
    .io_s(Walloc33bits_39_io_s)
  );
  Walloc33bits Walloc33bits_40 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_40_io_src_in),
    .io_cin(Walloc33bits_40_io_cin),
    .io_cout_group_0(Walloc33bits_40_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_40_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_40_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_40_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_40_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_40_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_40_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_40_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_40_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_40_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_40_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_40_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_40_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_40_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_40_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_40_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_40_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_40_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_40_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_40_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_40_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_40_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_40_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_40_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_40_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_40_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_40_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_40_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_40_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_40_io_cout_group_29),
    .io_cout(Walloc33bits_40_io_cout),
    .io_s(Walloc33bits_40_io_s)
  );
  Walloc33bits Walloc33bits_41 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_41_io_src_in),
    .io_cin(Walloc33bits_41_io_cin),
    .io_cout_group_0(Walloc33bits_41_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_41_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_41_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_41_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_41_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_41_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_41_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_41_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_41_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_41_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_41_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_41_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_41_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_41_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_41_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_41_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_41_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_41_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_41_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_41_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_41_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_41_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_41_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_41_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_41_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_41_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_41_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_41_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_41_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_41_io_cout_group_29),
    .io_cout(Walloc33bits_41_io_cout),
    .io_s(Walloc33bits_41_io_s)
  );
  Walloc33bits Walloc33bits_42 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_42_io_src_in),
    .io_cin(Walloc33bits_42_io_cin),
    .io_cout_group_0(Walloc33bits_42_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_42_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_42_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_42_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_42_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_42_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_42_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_42_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_42_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_42_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_42_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_42_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_42_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_42_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_42_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_42_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_42_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_42_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_42_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_42_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_42_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_42_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_42_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_42_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_42_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_42_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_42_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_42_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_42_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_42_io_cout_group_29),
    .io_cout(Walloc33bits_42_io_cout),
    .io_s(Walloc33bits_42_io_s)
  );
  Walloc33bits Walloc33bits_43 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_43_io_src_in),
    .io_cin(Walloc33bits_43_io_cin),
    .io_cout_group_0(Walloc33bits_43_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_43_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_43_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_43_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_43_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_43_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_43_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_43_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_43_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_43_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_43_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_43_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_43_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_43_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_43_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_43_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_43_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_43_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_43_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_43_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_43_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_43_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_43_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_43_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_43_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_43_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_43_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_43_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_43_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_43_io_cout_group_29),
    .io_cout(Walloc33bits_43_io_cout),
    .io_s(Walloc33bits_43_io_s)
  );
  Walloc33bits Walloc33bits_44 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_44_io_src_in),
    .io_cin(Walloc33bits_44_io_cin),
    .io_cout_group_0(Walloc33bits_44_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_44_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_44_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_44_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_44_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_44_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_44_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_44_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_44_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_44_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_44_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_44_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_44_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_44_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_44_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_44_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_44_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_44_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_44_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_44_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_44_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_44_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_44_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_44_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_44_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_44_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_44_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_44_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_44_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_44_io_cout_group_29),
    .io_cout(Walloc33bits_44_io_cout),
    .io_s(Walloc33bits_44_io_s)
  );
  Walloc33bits Walloc33bits_45 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_45_io_src_in),
    .io_cin(Walloc33bits_45_io_cin),
    .io_cout_group_0(Walloc33bits_45_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_45_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_45_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_45_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_45_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_45_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_45_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_45_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_45_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_45_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_45_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_45_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_45_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_45_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_45_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_45_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_45_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_45_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_45_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_45_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_45_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_45_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_45_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_45_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_45_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_45_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_45_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_45_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_45_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_45_io_cout_group_29),
    .io_cout(Walloc33bits_45_io_cout),
    .io_s(Walloc33bits_45_io_s)
  );
  Walloc33bits Walloc33bits_46 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_46_io_src_in),
    .io_cin(Walloc33bits_46_io_cin),
    .io_cout_group_0(Walloc33bits_46_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_46_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_46_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_46_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_46_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_46_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_46_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_46_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_46_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_46_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_46_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_46_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_46_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_46_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_46_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_46_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_46_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_46_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_46_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_46_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_46_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_46_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_46_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_46_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_46_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_46_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_46_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_46_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_46_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_46_io_cout_group_29),
    .io_cout(Walloc33bits_46_io_cout),
    .io_s(Walloc33bits_46_io_s)
  );
  Walloc33bits Walloc33bits_47 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_47_io_src_in),
    .io_cin(Walloc33bits_47_io_cin),
    .io_cout_group_0(Walloc33bits_47_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_47_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_47_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_47_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_47_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_47_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_47_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_47_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_47_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_47_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_47_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_47_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_47_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_47_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_47_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_47_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_47_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_47_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_47_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_47_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_47_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_47_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_47_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_47_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_47_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_47_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_47_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_47_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_47_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_47_io_cout_group_29),
    .io_cout(Walloc33bits_47_io_cout),
    .io_s(Walloc33bits_47_io_s)
  );
  Walloc33bits Walloc33bits_48 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_48_io_src_in),
    .io_cin(Walloc33bits_48_io_cin),
    .io_cout_group_0(Walloc33bits_48_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_48_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_48_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_48_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_48_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_48_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_48_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_48_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_48_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_48_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_48_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_48_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_48_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_48_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_48_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_48_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_48_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_48_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_48_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_48_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_48_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_48_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_48_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_48_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_48_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_48_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_48_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_48_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_48_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_48_io_cout_group_29),
    .io_cout(Walloc33bits_48_io_cout),
    .io_s(Walloc33bits_48_io_s)
  );
  Walloc33bits Walloc33bits_49 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_49_io_src_in),
    .io_cin(Walloc33bits_49_io_cin),
    .io_cout_group_0(Walloc33bits_49_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_49_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_49_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_49_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_49_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_49_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_49_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_49_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_49_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_49_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_49_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_49_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_49_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_49_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_49_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_49_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_49_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_49_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_49_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_49_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_49_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_49_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_49_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_49_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_49_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_49_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_49_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_49_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_49_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_49_io_cout_group_29),
    .io_cout(Walloc33bits_49_io_cout),
    .io_s(Walloc33bits_49_io_s)
  );
  Walloc33bits Walloc33bits_50 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_50_io_src_in),
    .io_cin(Walloc33bits_50_io_cin),
    .io_cout_group_0(Walloc33bits_50_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_50_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_50_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_50_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_50_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_50_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_50_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_50_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_50_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_50_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_50_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_50_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_50_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_50_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_50_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_50_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_50_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_50_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_50_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_50_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_50_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_50_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_50_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_50_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_50_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_50_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_50_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_50_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_50_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_50_io_cout_group_29),
    .io_cout(Walloc33bits_50_io_cout),
    .io_s(Walloc33bits_50_io_s)
  );
  Walloc33bits Walloc33bits_51 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_51_io_src_in),
    .io_cin(Walloc33bits_51_io_cin),
    .io_cout_group_0(Walloc33bits_51_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_51_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_51_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_51_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_51_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_51_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_51_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_51_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_51_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_51_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_51_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_51_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_51_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_51_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_51_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_51_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_51_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_51_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_51_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_51_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_51_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_51_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_51_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_51_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_51_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_51_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_51_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_51_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_51_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_51_io_cout_group_29),
    .io_cout(Walloc33bits_51_io_cout),
    .io_s(Walloc33bits_51_io_s)
  );
  Walloc33bits Walloc33bits_52 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_52_io_src_in),
    .io_cin(Walloc33bits_52_io_cin),
    .io_cout_group_0(Walloc33bits_52_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_52_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_52_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_52_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_52_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_52_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_52_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_52_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_52_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_52_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_52_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_52_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_52_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_52_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_52_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_52_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_52_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_52_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_52_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_52_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_52_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_52_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_52_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_52_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_52_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_52_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_52_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_52_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_52_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_52_io_cout_group_29),
    .io_cout(Walloc33bits_52_io_cout),
    .io_s(Walloc33bits_52_io_s)
  );
  Walloc33bits Walloc33bits_53 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_53_io_src_in),
    .io_cin(Walloc33bits_53_io_cin),
    .io_cout_group_0(Walloc33bits_53_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_53_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_53_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_53_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_53_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_53_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_53_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_53_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_53_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_53_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_53_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_53_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_53_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_53_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_53_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_53_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_53_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_53_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_53_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_53_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_53_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_53_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_53_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_53_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_53_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_53_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_53_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_53_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_53_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_53_io_cout_group_29),
    .io_cout(Walloc33bits_53_io_cout),
    .io_s(Walloc33bits_53_io_s)
  );
  Walloc33bits Walloc33bits_54 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_54_io_src_in),
    .io_cin(Walloc33bits_54_io_cin),
    .io_cout_group_0(Walloc33bits_54_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_54_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_54_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_54_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_54_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_54_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_54_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_54_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_54_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_54_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_54_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_54_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_54_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_54_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_54_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_54_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_54_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_54_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_54_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_54_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_54_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_54_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_54_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_54_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_54_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_54_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_54_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_54_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_54_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_54_io_cout_group_29),
    .io_cout(Walloc33bits_54_io_cout),
    .io_s(Walloc33bits_54_io_s)
  );
  Walloc33bits Walloc33bits_55 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_55_io_src_in),
    .io_cin(Walloc33bits_55_io_cin),
    .io_cout_group_0(Walloc33bits_55_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_55_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_55_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_55_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_55_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_55_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_55_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_55_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_55_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_55_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_55_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_55_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_55_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_55_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_55_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_55_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_55_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_55_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_55_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_55_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_55_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_55_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_55_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_55_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_55_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_55_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_55_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_55_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_55_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_55_io_cout_group_29),
    .io_cout(Walloc33bits_55_io_cout),
    .io_s(Walloc33bits_55_io_s)
  );
  Walloc33bits Walloc33bits_56 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_56_io_src_in),
    .io_cin(Walloc33bits_56_io_cin),
    .io_cout_group_0(Walloc33bits_56_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_56_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_56_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_56_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_56_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_56_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_56_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_56_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_56_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_56_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_56_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_56_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_56_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_56_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_56_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_56_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_56_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_56_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_56_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_56_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_56_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_56_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_56_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_56_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_56_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_56_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_56_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_56_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_56_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_56_io_cout_group_29),
    .io_cout(Walloc33bits_56_io_cout),
    .io_s(Walloc33bits_56_io_s)
  );
  Walloc33bits Walloc33bits_57 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_57_io_src_in),
    .io_cin(Walloc33bits_57_io_cin),
    .io_cout_group_0(Walloc33bits_57_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_57_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_57_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_57_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_57_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_57_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_57_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_57_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_57_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_57_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_57_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_57_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_57_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_57_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_57_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_57_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_57_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_57_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_57_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_57_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_57_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_57_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_57_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_57_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_57_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_57_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_57_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_57_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_57_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_57_io_cout_group_29),
    .io_cout(Walloc33bits_57_io_cout),
    .io_s(Walloc33bits_57_io_s)
  );
  Walloc33bits Walloc33bits_58 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_58_io_src_in),
    .io_cin(Walloc33bits_58_io_cin),
    .io_cout_group_0(Walloc33bits_58_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_58_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_58_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_58_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_58_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_58_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_58_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_58_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_58_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_58_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_58_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_58_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_58_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_58_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_58_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_58_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_58_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_58_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_58_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_58_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_58_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_58_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_58_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_58_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_58_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_58_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_58_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_58_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_58_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_58_io_cout_group_29),
    .io_cout(Walloc33bits_58_io_cout),
    .io_s(Walloc33bits_58_io_s)
  );
  Walloc33bits Walloc33bits_59 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_59_io_src_in),
    .io_cin(Walloc33bits_59_io_cin),
    .io_cout_group_0(Walloc33bits_59_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_59_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_59_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_59_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_59_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_59_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_59_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_59_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_59_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_59_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_59_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_59_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_59_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_59_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_59_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_59_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_59_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_59_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_59_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_59_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_59_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_59_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_59_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_59_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_59_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_59_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_59_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_59_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_59_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_59_io_cout_group_29),
    .io_cout(Walloc33bits_59_io_cout),
    .io_s(Walloc33bits_59_io_s)
  );
  Walloc33bits Walloc33bits_60 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_60_io_src_in),
    .io_cin(Walloc33bits_60_io_cin),
    .io_cout_group_0(Walloc33bits_60_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_60_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_60_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_60_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_60_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_60_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_60_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_60_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_60_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_60_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_60_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_60_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_60_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_60_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_60_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_60_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_60_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_60_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_60_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_60_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_60_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_60_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_60_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_60_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_60_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_60_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_60_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_60_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_60_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_60_io_cout_group_29),
    .io_cout(Walloc33bits_60_io_cout),
    .io_s(Walloc33bits_60_io_s)
  );
  Walloc33bits Walloc33bits_61 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_61_io_src_in),
    .io_cin(Walloc33bits_61_io_cin),
    .io_cout_group_0(Walloc33bits_61_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_61_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_61_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_61_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_61_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_61_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_61_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_61_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_61_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_61_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_61_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_61_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_61_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_61_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_61_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_61_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_61_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_61_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_61_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_61_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_61_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_61_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_61_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_61_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_61_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_61_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_61_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_61_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_61_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_61_io_cout_group_29),
    .io_cout(Walloc33bits_61_io_cout),
    .io_s(Walloc33bits_61_io_s)
  );
  Walloc33bits Walloc33bits_62 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_62_io_src_in),
    .io_cin(Walloc33bits_62_io_cin),
    .io_cout_group_0(Walloc33bits_62_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_62_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_62_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_62_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_62_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_62_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_62_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_62_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_62_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_62_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_62_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_62_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_62_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_62_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_62_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_62_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_62_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_62_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_62_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_62_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_62_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_62_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_62_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_62_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_62_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_62_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_62_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_62_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_62_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_62_io_cout_group_29),
    .io_cout(Walloc33bits_62_io_cout),
    .io_s(Walloc33bits_62_io_s)
  );
  Walloc33bits Walloc33bits_63 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_63_io_src_in),
    .io_cin(Walloc33bits_63_io_cin),
    .io_cout_group_0(Walloc33bits_63_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_63_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_63_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_63_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_63_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_63_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_63_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_63_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_63_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_63_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_63_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_63_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_63_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_63_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_63_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_63_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_63_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_63_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_63_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_63_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_63_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_63_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_63_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_63_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_63_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_63_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_63_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_63_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_63_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_63_io_cout_group_29),
    .io_cout(Walloc33bits_63_io_cout),
    .io_s(Walloc33bits_63_io_s)
  );
  Walloc33bits Walloc33bits_64 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_64_io_src_in),
    .io_cin(Walloc33bits_64_io_cin),
    .io_cout_group_0(Walloc33bits_64_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_64_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_64_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_64_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_64_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_64_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_64_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_64_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_64_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_64_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_64_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_64_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_64_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_64_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_64_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_64_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_64_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_64_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_64_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_64_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_64_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_64_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_64_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_64_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_64_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_64_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_64_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_64_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_64_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_64_io_cout_group_29),
    .io_cout(Walloc33bits_64_io_cout),
    .io_s(Walloc33bits_64_io_s)
  );
  Walloc33bits Walloc33bits_65 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_65_io_src_in),
    .io_cin(Walloc33bits_65_io_cin),
    .io_cout_group_0(Walloc33bits_65_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_65_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_65_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_65_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_65_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_65_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_65_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_65_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_65_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_65_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_65_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_65_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_65_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_65_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_65_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_65_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_65_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_65_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_65_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_65_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_65_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_65_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_65_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_65_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_65_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_65_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_65_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_65_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_65_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_65_io_cout_group_29),
    .io_cout(Walloc33bits_65_io_cout),
    .io_s(Walloc33bits_65_io_s)
  );
  Walloc33bits Walloc33bits_66 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_66_io_src_in),
    .io_cin(Walloc33bits_66_io_cin),
    .io_cout_group_0(Walloc33bits_66_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_66_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_66_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_66_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_66_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_66_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_66_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_66_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_66_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_66_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_66_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_66_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_66_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_66_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_66_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_66_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_66_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_66_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_66_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_66_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_66_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_66_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_66_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_66_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_66_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_66_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_66_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_66_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_66_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_66_io_cout_group_29),
    .io_cout(Walloc33bits_66_io_cout),
    .io_s(Walloc33bits_66_io_s)
  );
  Walloc33bits Walloc33bits_67 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_67_io_src_in),
    .io_cin(Walloc33bits_67_io_cin),
    .io_cout_group_0(Walloc33bits_67_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_67_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_67_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_67_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_67_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_67_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_67_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_67_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_67_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_67_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_67_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_67_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_67_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_67_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_67_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_67_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_67_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_67_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_67_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_67_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_67_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_67_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_67_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_67_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_67_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_67_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_67_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_67_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_67_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_67_io_cout_group_29),
    .io_cout(Walloc33bits_67_io_cout),
    .io_s(Walloc33bits_67_io_s)
  );
  Walloc33bits Walloc33bits_68 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_68_io_src_in),
    .io_cin(Walloc33bits_68_io_cin),
    .io_cout_group_0(Walloc33bits_68_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_68_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_68_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_68_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_68_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_68_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_68_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_68_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_68_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_68_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_68_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_68_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_68_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_68_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_68_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_68_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_68_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_68_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_68_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_68_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_68_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_68_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_68_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_68_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_68_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_68_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_68_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_68_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_68_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_68_io_cout_group_29),
    .io_cout(Walloc33bits_68_io_cout),
    .io_s(Walloc33bits_68_io_s)
  );
  Walloc33bits Walloc33bits_69 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_69_io_src_in),
    .io_cin(Walloc33bits_69_io_cin),
    .io_cout_group_0(Walloc33bits_69_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_69_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_69_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_69_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_69_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_69_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_69_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_69_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_69_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_69_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_69_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_69_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_69_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_69_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_69_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_69_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_69_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_69_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_69_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_69_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_69_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_69_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_69_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_69_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_69_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_69_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_69_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_69_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_69_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_69_io_cout_group_29),
    .io_cout(Walloc33bits_69_io_cout),
    .io_s(Walloc33bits_69_io_s)
  );
  Walloc33bits Walloc33bits_70 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_70_io_src_in),
    .io_cin(Walloc33bits_70_io_cin),
    .io_cout_group_0(Walloc33bits_70_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_70_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_70_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_70_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_70_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_70_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_70_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_70_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_70_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_70_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_70_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_70_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_70_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_70_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_70_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_70_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_70_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_70_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_70_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_70_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_70_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_70_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_70_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_70_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_70_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_70_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_70_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_70_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_70_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_70_io_cout_group_29),
    .io_cout(Walloc33bits_70_io_cout),
    .io_s(Walloc33bits_70_io_s)
  );
  Walloc33bits Walloc33bits_71 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_71_io_src_in),
    .io_cin(Walloc33bits_71_io_cin),
    .io_cout_group_0(Walloc33bits_71_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_71_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_71_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_71_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_71_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_71_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_71_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_71_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_71_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_71_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_71_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_71_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_71_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_71_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_71_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_71_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_71_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_71_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_71_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_71_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_71_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_71_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_71_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_71_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_71_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_71_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_71_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_71_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_71_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_71_io_cout_group_29),
    .io_cout(Walloc33bits_71_io_cout),
    .io_s(Walloc33bits_71_io_s)
  );
  Walloc33bits Walloc33bits_72 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_72_io_src_in),
    .io_cin(Walloc33bits_72_io_cin),
    .io_cout_group_0(Walloc33bits_72_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_72_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_72_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_72_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_72_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_72_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_72_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_72_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_72_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_72_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_72_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_72_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_72_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_72_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_72_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_72_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_72_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_72_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_72_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_72_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_72_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_72_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_72_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_72_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_72_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_72_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_72_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_72_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_72_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_72_io_cout_group_29),
    .io_cout(Walloc33bits_72_io_cout),
    .io_s(Walloc33bits_72_io_s)
  );
  Walloc33bits Walloc33bits_73 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_73_io_src_in),
    .io_cin(Walloc33bits_73_io_cin),
    .io_cout_group_0(Walloc33bits_73_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_73_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_73_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_73_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_73_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_73_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_73_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_73_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_73_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_73_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_73_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_73_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_73_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_73_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_73_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_73_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_73_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_73_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_73_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_73_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_73_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_73_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_73_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_73_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_73_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_73_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_73_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_73_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_73_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_73_io_cout_group_29),
    .io_cout(Walloc33bits_73_io_cout),
    .io_s(Walloc33bits_73_io_s)
  );
  Walloc33bits Walloc33bits_74 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_74_io_src_in),
    .io_cin(Walloc33bits_74_io_cin),
    .io_cout_group_0(Walloc33bits_74_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_74_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_74_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_74_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_74_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_74_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_74_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_74_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_74_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_74_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_74_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_74_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_74_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_74_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_74_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_74_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_74_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_74_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_74_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_74_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_74_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_74_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_74_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_74_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_74_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_74_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_74_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_74_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_74_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_74_io_cout_group_29),
    .io_cout(Walloc33bits_74_io_cout),
    .io_s(Walloc33bits_74_io_s)
  );
  Walloc33bits Walloc33bits_75 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_75_io_src_in),
    .io_cin(Walloc33bits_75_io_cin),
    .io_cout_group_0(Walloc33bits_75_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_75_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_75_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_75_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_75_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_75_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_75_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_75_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_75_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_75_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_75_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_75_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_75_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_75_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_75_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_75_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_75_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_75_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_75_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_75_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_75_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_75_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_75_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_75_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_75_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_75_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_75_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_75_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_75_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_75_io_cout_group_29),
    .io_cout(Walloc33bits_75_io_cout),
    .io_s(Walloc33bits_75_io_s)
  );
  Walloc33bits Walloc33bits_76 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_76_io_src_in),
    .io_cin(Walloc33bits_76_io_cin),
    .io_cout_group_0(Walloc33bits_76_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_76_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_76_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_76_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_76_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_76_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_76_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_76_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_76_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_76_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_76_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_76_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_76_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_76_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_76_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_76_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_76_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_76_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_76_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_76_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_76_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_76_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_76_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_76_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_76_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_76_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_76_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_76_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_76_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_76_io_cout_group_29),
    .io_cout(Walloc33bits_76_io_cout),
    .io_s(Walloc33bits_76_io_s)
  );
  Walloc33bits Walloc33bits_77 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_77_io_src_in),
    .io_cin(Walloc33bits_77_io_cin),
    .io_cout_group_0(Walloc33bits_77_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_77_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_77_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_77_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_77_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_77_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_77_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_77_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_77_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_77_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_77_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_77_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_77_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_77_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_77_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_77_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_77_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_77_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_77_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_77_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_77_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_77_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_77_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_77_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_77_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_77_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_77_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_77_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_77_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_77_io_cout_group_29),
    .io_cout(Walloc33bits_77_io_cout),
    .io_s(Walloc33bits_77_io_s)
  );
  Walloc33bits Walloc33bits_78 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_78_io_src_in),
    .io_cin(Walloc33bits_78_io_cin),
    .io_cout_group_0(Walloc33bits_78_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_78_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_78_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_78_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_78_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_78_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_78_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_78_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_78_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_78_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_78_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_78_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_78_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_78_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_78_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_78_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_78_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_78_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_78_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_78_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_78_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_78_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_78_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_78_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_78_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_78_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_78_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_78_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_78_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_78_io_cout_group_29),
    .io_cout(Walloc33bits_78_io_cout),
    .io_s(Walloc33bits_78_io_s)
  );
  Walloc33bits Walloc33bits_79 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_79_io_src_in),
    .io_cin(Walloc33bits_79_io_cin),
    .io_cout_group_0(Walloc33bits_79_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_79_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_79_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_79_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_79_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_79_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_79_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_79_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_79_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_79_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_79_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_79_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_79_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_79_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_79_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_79_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_79_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_79_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_79_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_79_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_79_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_79_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_79_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_79_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_79_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_79_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_79_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_79_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_79_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_79_io_cout_group_29),
    .io_cout(Walloc33bits_79_io_cout),
    .io_s(Walloc33bits_79_io_s)
  );
  Walloc33bits Walloc33bits_80 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_80_io_src_in),
    .io_cin(Walloc33bits_80_io_cin),
    .io_cout_group_0(Walloc33bits_80_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_80_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_80_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_80_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_80_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_80_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_80_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_80_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_80_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_80_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_80_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_80_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_80_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_80_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_80_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_80_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_80_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_80_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_80_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_80_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_80_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_80_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_80_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_80_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_80_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_80_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_80_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_80_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_80_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_80_io_cout_group_29),
    .io_cout(Walloc33bits_80_io_cout),
    .io_s(Walloc33bits_80_io_s)
  );
  Walloc33bits Walloc33bits_81 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_81_io_src_in),
    .io_cin(Walloc33bits_81_io_cin),
    .io_cout_group_0(Walloc33bits_81_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_81_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_81_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_81_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_81_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_81_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_81_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_81_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_81_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_81_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_81_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_81_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_81_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_81_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_81_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_81_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_81_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_81_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_81_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_81_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_81_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_81_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_81_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_81_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_81_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_81_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_81_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_81_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_81_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_81_io_cout_group_29),
    .io_cout(Walloc33bits_81_io_cout),
    .io_s(Walloc33bits_81_io_s)
  );
  Walloc33bits Walloc33bits_82 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_82_io_src_in),
    .io_cin(Walloc33bits_82_io_cin),
    .io_cout_group_0(Walloc33bits_82_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_82_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_82_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_82_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_82_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_82_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_82_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_82_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_82_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_82_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_82_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_82_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_82_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_82_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_82_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_82_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_82_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_82_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_82_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_82_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_82_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_82_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_82_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_82_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_82_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_82_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_82_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_82_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_82_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_82_io_cout_group_29),
    .io_cout(Walloc33bits_82_io_cout),
    .io_s(Walloc33bits_82_io_s)
  );
  Walloc33bits Walloc33bits_83 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_83_io_src_in),
    .io_cin(Walloc33bits_83_io_cin),
    .io_cout_group_0(Walloc33bits_83_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_83_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_83_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_83_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_83_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_83_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_83_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_83_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_83_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_83_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_83_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_83_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_83_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_83_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_83_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_83_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_83_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_83_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_83_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_83_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_83_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_83_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_83_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_83_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_83_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_83_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_83_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_83_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_83_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_83_io_cout_group_29),
    .io_cout(Walloc33bits_83_io_cout),
    .io_s(Walloc33bits_83_io_s)
  );
  Walloc33bits Walloc33bits_84 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_84_io_src_in),
    .io_cin(Walloc33bits_84_io_cin),
    .io_cout_group_0(Walloc33bits_84_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_84_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_84_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_84_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_84_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_84_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_84_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_84_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_84_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_84_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_84_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_84_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_84_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_84_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_84_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_84_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_84_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_84_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_84_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_84_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_84_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_84_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_84_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_84_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_84_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_84_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_84_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_84_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_84_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_84_io_cout_group_29),
    .io_cout(Walloc33bits_84_io_cout),
    .io_s(Walloc33bits_84_io_s)
  );
  Walloc33bits Walloc33bits_85 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_85_io_src_in),
    .io_cin(Walloc33bits_85_io_cin),
    .io_cout_group_0(Walloc33bits_85_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_85_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_85_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_85_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_85_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_85_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_85_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_85_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_85_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_85_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_85_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_85_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_85_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_85_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_85_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_85_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_85_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_85_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_85_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_85_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_85_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_85_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_85_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_85_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_85_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_85_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_85_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_85_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_85_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_85_io_cout_group_29),
    .io_cout(Walloc33bits_85_io_cout),
    .io_s(Walloc33bits_85_io_s)
  );
  Walloc33bits Walloc33bits_86 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_86_io_src_in),
    .io_cin(Walloc33bits_86_io_cin),
    .io_cout_group_0(Walloc33bits_86_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_86_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_86_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_86_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_86_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_86_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_86_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_86_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_86_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_86_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_86_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_86_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_86_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_86_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_86_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_86_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_86_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_86_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_86_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_86_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_86_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_86_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_86_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_86_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_86_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_86_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_86_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_86_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_86_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_86_io_cout_group_29),
    .io_cout(Walloc33bits_86_io_cout),
    .io_s(Walloc33bits_86_io_s)
  );
  Walloc33bits Walloc33bits_87 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_87_io_src_in),
    .io_cin(Walloc33bits_87_io_cin),
    .io_cout_group_0(Walloc33bits_87_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_87_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_87_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_87_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_87_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_87_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_87_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_87_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_87_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_87_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_87_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_87_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_87_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_87_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_87_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_87_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_87_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_87_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_87_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_87_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_87_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_87_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_87_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_87_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_87_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_87_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_87_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_87_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_87_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_87_io_cout_group_29),
    .io_cout(Walloc33bits_87_io_cout),
    .io_s(Walloc33bits_87_io_s)
  );
  Walloc33bits Walloc33bits_88 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_88_io_src_in),
    .io_cin(Walloc33bits_88_io_cin),
    .io_cout_group_0(Walloc33bits_88_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_88_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_88_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_88_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_88_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_88_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_88_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_88_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_88_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_88_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_88_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_88_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_88_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_88_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_88_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_88_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_88_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_88_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_88_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_88_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_88_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_88_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_88_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_88_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_88_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_88_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_88_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_88_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_88_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_88_io_cout_group_29),
    .io_cout(Walloc33bits_88_io_cout),
    .io_s(Walloc33bits_88_io_s)
  );
  Walloc33bits Walloc33bits_89 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_89_io_src_in),
    .io_cin(Walloc33bits_89_io_cin),
    .io_cout_group_0(Walloc33bits_89_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_89_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_89_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_89_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_89_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_89_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_89_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_89_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_89_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_89_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_89_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_89_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_89_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_89_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_89_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_89_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_89_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_89_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_89_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_89_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_89_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_89_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_89_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_89_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_89_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_89_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_89_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_89_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_89_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_89_io_cout_group_29),
    .io_cout(Walloc33bits_89_io_cout),
    .io_s(Walloc33bits_89_io_s)
  );
  Walloc33bits Walloc33bits_90 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_90_io_src_in),
    .io_cin(Walloc33bits_90_io_cin),
    .io_cout_group_0(Walloc33bits_90_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_90_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_90_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_90_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_90_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_90_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_90_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_90_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_90_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_90_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_90_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_90_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_90_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_90_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_90_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_90_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_90_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_90_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_90_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_90_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_90_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_90_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_90_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_90_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_90_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_90_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_90_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_90_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_90_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_90_io_cout_group_29),
    .io_cout(Walloc33bits_90_io_cout),
    .io_s(Walloc33bits_90_io_s)
  );
  Walloc33bits Walloc33bits_91 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_91_io_src_in),
    .io_cin(Walloc33bits_91_io_cin),
    .io_cout_group_0(Walloc33bits_91_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_91_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_91_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_91_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_91_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_91_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_91_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_91_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_91_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_91_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_91_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_91_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_91_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_91_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_91_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_91_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_91_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_91_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_91_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_91_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_91_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_91_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_91_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_91_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_91_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_91_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_91_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_91_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_91_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_91_io_cout_group_29),
    .io_cout(Walloc33bits_91_io_cout),
    .io_s(Walloc33bits_91_io_s)
  );
  Walloc33bits Walloc33bits_92 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_92_io_src_in),
    .io_cin(Walloc33bits_92_io_cin),
    .io_cout_group_0(Walloc33bits_92_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_92_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_92_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_92_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_92_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_92_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_92_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_92_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_92_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_92_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_92_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_92_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_92_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_92_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_92_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_92_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_92_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_92_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_92_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_92_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_92_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_92_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_92_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_92_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_92_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_92_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_92_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_92_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_92_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_92_io_cout_group_29),
    .io_cout(Walloc33bits_92_io_cout),
    .io_s(Walloc33bits_92_io_s)
  );
  Walloc33bits Walloc33bits_93 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_93_io_src_in),
    .io_cin(Walloc33bits_93_io_cin),
    .io_cout_group_0(Walloc33bits_93_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_93_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_93_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_93_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_93_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_93_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_93_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_93_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_93_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_93_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_93_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_93_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_93_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_93_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_93_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_93_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_93_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_93_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_93_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_93_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_93_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_93_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_93_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_93_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_93_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_93_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_93_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_93_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_93_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_93_io_cout_group_29),
    .io_cout(Walloc33bits_93_io_cout),
    .io_s(Walloc33bits_93_io_s)
  );
  Walloc33bits Walloc33bits_94 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_94_io_src_in),
    .io_cin(Walloc33bits_94_io_cin),
    .io_cout_group_0(Walloc33bits_94_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_94_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_94_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_94_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_94_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_94_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_94_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_94_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_94_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_94_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_94_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_94_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_94_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_94_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_94_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_94_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_94_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_94_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_94_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_94_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_94_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_94_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_94_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_94_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_94_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_94_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_94_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_94_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_94_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_94_io_cout_group_29),
    .io_cout(Walloc33bits_94_io_cout),
    .io_s(Walloc33bits_94_io_s)
  );
  Walloc33bits Walloc33bits_95 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_95_io_src_in),
    .io_cin(Walloc33bits_95_io_cin),
    .io_cout_group_0(Walloc33bits_95_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_95_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_95_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_95_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_95_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_95_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_95_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_95_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_95_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_95_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_95_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_95_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_95_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_95_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_95_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_95_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_95_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_95_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_95_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_95_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_95_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_95_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_95_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_95_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_95_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_95_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_95_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_95_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_95_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_95_io_cout_group_29),
    .io_cout(Walloc33bits_95_io_cout),
    .io_s(Walloc33bits_95_io_s)
  );
  Walloc33bits Walloc33bits_96 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_96_io_src_in),
    .io_cin(Walloc33bits_96_io_cin),
    .io_cout_group_0(Walloc33bits_96_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_96_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_96_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_96_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_96_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_96_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_96_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_96_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_96_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_96_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_96_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_96_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_96_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_96_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_96_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_96_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_96_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_96_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_96_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_96_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_96_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_96_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_96_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_96_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_96_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_96_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_96_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_96_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_96_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_96_io_cout_group_29),
    .io_cout(Walloc33bits_96_io_cout),
    .io_s(Walloc33bits_96_io_s)
  );
  Walloc33bits Walloc33bits_97 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_97_io_src_in),
    .io_cin(Walloc33bits_97_io_cin),
    .io_cout_group_0(Walloc33bits_97_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_97_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_97_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_97_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_97_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_97_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_97_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_97_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_97_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_97_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_97_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_97_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_97_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_97_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_97_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_97_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_97_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_97_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_97_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_97_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_97_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_97_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_97_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_97_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_97_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_97_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_97_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_97_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_97_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_97_io_cout_group_29),
    .io_cout(Walloc33bits_97_io_cout),
    .io_s(Walloc33bits_97_io_s)
  );
  Walloc33bits Walloc33bits_98 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_98_io_src_in),
    .io_cin(Walloc33bits_98_io_cin),
    .io_cout_group_0(Walloc33bits_98_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_98_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_98_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_98_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_98_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_98_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_98_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_98_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_98_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_98_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_98_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_98_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_98_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_98_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_98_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_98_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_98_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_98_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_98_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_98_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_98_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_98_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_98_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_98_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_98_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_98_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_98_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_98_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_98_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_98_io_cout_group_29),
    .io_cout(Walloc33bits_98_io_cout),
    .io_s(Walloc33bits_98_io_s)
  );
  Walloc33bits Walloc33bits_99 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_99_io_src_in),
    .io_cin(Walloc33bits_99_io_cin),
    .io_cout_group_0(Walloc33bits_99_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_99_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_99_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_99_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_99_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_99_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_99_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_99_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_99_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_99_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_99_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_99_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_99_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_99_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_99_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_99_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_99_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_99_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_99_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_99_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_99_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_99_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_99_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_99_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_99_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_99_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_99_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_99_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_99_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_99_io_cout_group_29),
    .io_cout(Walloc33bits_99_io_cout),
    .io_s(Walloc33bits_99_io_s)
  );
  Walloc33bits Walloc33bits_100 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_100_io_src_in),
    .io_cin(Walloc33bits_100_io_cin),
    .io_cout_group_0(Walloc33bits_100_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_100_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_100_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_100_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_100_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_100_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_100_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_100_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_100_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_100_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_100_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_100_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_100_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_100_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_100_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_100_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_100_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_100_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_100_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_100_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_100_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_100_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_100_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_100_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_100_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_100_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_100_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_100_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_100_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_100_io_cout_group_29),
    .io_cout(Walloc33bits_100_io_cout),
    .io_s(Walloc33bits_100_io_s)
  );
  Walloc33bits Walloc33bits_101 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_101_io_src_in),
    .io_cin(Walloc33bits_101_io_cin),
    .io_cout_group_0(Walloc33bits_101_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_101_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_101_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_101_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_101_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_101_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_101_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_101_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_101_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_101_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_101_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_101_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_101_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_101_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_101_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_101_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_101_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_101_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_101_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_101_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_101_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_101_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_101_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_101_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_101_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_101_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_101_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_101_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_101_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_101_io_cout_group_29),
    .io_cout(Walloc33bits_101_io_cout),
    .io_s(Walloc33bits_101_io_s)
  );
  Walloc33bits Walloc33bits_102 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_102_io_src_in),
    .io_cin(Walloc33bits_102_io_cin),
    .io_cout_group_0(Walloc33bits_102_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_102_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_102_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_102_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_102_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_102_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_102_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_102_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_102_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_102_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_102_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_102_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_102_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_102_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_102_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_102_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_102_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_102_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_102_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_102_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_102_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_102_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_102_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_102_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_102_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_102_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_102_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_102_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_102_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_102_io_cout_group_29),
    .io_cout(Walloc33bits_102_io_cout),
    .io_s(Walloc33bits_102_io_s)
  );
  Walloc33bits Walloc33bits_103 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_103_io_src_in),
    .io_cin(Walloc33bits_103_io_cin),
    .io_cout_group_0(Walloc33bits_103_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_103_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_103_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_103_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_103_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_103_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_103_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_103_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_103_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_103_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_103_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_103_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_103_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_103_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_103_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_103_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_103_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_103_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_103_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_103_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_103_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_103_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_103_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_103_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_103_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_103_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_103_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_103_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_103_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_103_io_cout_group_29),
    .io_cout(Walloc33bits_103_io_cout),
    .io_s(Walloc33bits_103_io_s)
  );
  Walloc33bits Walloc33bits_104 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_104_io_src_in),
    .io_cin(Walloc33bits_104_io_cin),
    .io_cout_group_0(Walloc33bits_104_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_104_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_104_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_104_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_104_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_104_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_104_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_104_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_104_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_104_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_104_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_104_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_104_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_104_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_104_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_104_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_104_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_104_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_104_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_104_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_104_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_104_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_104_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_104_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_104_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_104_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_104_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_104_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_104_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_104_io_cout_group_29),
    .io_cout(Walloc33bits_104_io_cout),
    .io_s(Walloc33bits_104_io_s)
  );
  Walloc33bits Walloc33bits_105 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_105_io_src_in),
    .io_cin(Walloc33bits_105_io_cin),
    .io_cout_group_0(Walloc33bits_105_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_105_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_105_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_105_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_105_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_105_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_105_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_105_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_105_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_105_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_105_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_105_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_105_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_105_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_105_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_105_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_105_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_105_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_105_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_105_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_105_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_105_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_105_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_105_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_105_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_105_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_105_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_105_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_105_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_105_io_cout_group_29),
    .io_cout(Walloc33bits_105_io_cout),
    .io_s(Walloc33bits_105_io_s)
  );
  Walloc33bits Walloc33bits_106 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_106_io_src_in),
    .io_cin(Walloc33bits_106_io_cin),
    .io_cout_group_0(Walloc33bits_106_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_106_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_106_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_106_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_106_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_106_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_106_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_106_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_106_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_106_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_106_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_106_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_106_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_106_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_106_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_106_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_106_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_106_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_106_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_106_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_106_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_106_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_106_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_106_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_106_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_106_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_106_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_106_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_106_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_106_io_cout_group_29),
    .io_cout(Walloc33bits_106_io_cout),
    .io_s(Walloc33bits_106_io_s)
  );
  Walloc33bits Walloc33bits_107 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_107_io_src_in),
    .io_cin(Walloc33bits_107_io_cin),
    .io_cout_group_0(Walloc33bits_107_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_107_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_107_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_107_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_107_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_107_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_107_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_107_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_107_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_107_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_107_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_107_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_107_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_107_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_107_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_107_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_107_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_107_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_107_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_107_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_107_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_107_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_107_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_107_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_107_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_107_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_107_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_107_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_107_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_107_io_cout_group_29),
    .io_cout(Walloc33bits_107_io_cout),
    .io_s(Walloc33bits_107_io_s)
  );
  Walloc33bits Walloc33bits_108 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_108_io_src_in),
    .io_cin(Walloc33bits_108_io_cin),
    .io_cout_group_0(Walloc33bits_108_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_108_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_108_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_108_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_108_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_108_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_108_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_108_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_108_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_108_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_108_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_108_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_108_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_108_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_108_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_108_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_108_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_108_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_108_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_108_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_108_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_108_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_108_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_108_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_108_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_108_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_108_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_108_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_108_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_108_io_cout_group_29),
    .io_cout(Walloc33bits_108_io_cout),
    .io_s(Walloc33bits_108_io_s)
  );
  Walloc33bits Walloc33bits_109 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_109_io_src_in),
    .io_cin(Walloc33bits_109_io_cin),
    .io_cout_group_0(Walloc33bits_109_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_109_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_109_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_109_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_109_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_109_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_109_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_109_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_109_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_109_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_109_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_109_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_109_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_109_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_109_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_109_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_109_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_109_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_109_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_109_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_109_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_109_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_109_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_109_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_109_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_109_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_109_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_109_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_109_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_109_io_cout_group_29),
    .io_cout(Walloc33bits_109_io_cout),
    .io_s(Walloc33bits_109_io_s)
  );
  Walloc33bits Walloc33bits_110 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_110_io_src_in),
    .io_cin(Walloc33bits_110_io_cin),
    .io_cout_group_0(Walloc33bits_110_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_110_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_110_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_110_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_110_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_110_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_110_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_110_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_110_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_110_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_110_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_110_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_110_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_110_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_110_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_110_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_110_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_110_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_110_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_110_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_110_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_110_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_110_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_110_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_110_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_110_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_110_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_110_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_110_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_110_io_cout_group_29),
    .io_cout(Walloc33bits_110_io_cout),
    .io_s(Walloc33bits_110_io_s)
  );
  Walloc33bits Walloc33bits_111 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_111_io_src_in),
    .io_cin(Walloc33bits_111_io_cin),
    .io_cout_group_0(Walloc33bits_111_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_111_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_111_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_111_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_111_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_111_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_111_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_111_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_111_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_111_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_111_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_111_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_111_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_111_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_111_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_111_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_111_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_111_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_111_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_111_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_111_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_111_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_111_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_111_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_111_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_111_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_111_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_111_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_111_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_111_io_cout_group_29),
    .io_cout(Walloc33bits_111_io_cout),
    .io_s(Walloc33bits_111_io_s)
  );
  Walloc33bits Walloc33bits_112 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_112_io_src_in),
    .io_cin(Walloc33bits_112_io_cin),
    .io_cout_group_0(Walloc33bits_112_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_112_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_112_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_112_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_112_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_112_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_112_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_112_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_112_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_112_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_112_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_112_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_112_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_112_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_112_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_112_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_112_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_112_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_112_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_112_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_112_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_112_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_112_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_112_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_112_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_112_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_112_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_112_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_112_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_112_io_cout_group_29),
    .io_cout(Walloc33bits_112_io_cout),
    .io_s(Walloc33bits_112_io_s)
  );
  Walloc33bits Walloc33bits_113 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_113_io_src_in),
    .io_cin(Walloc33bits_113_io_cin),
    .io_cout_group_0(Walloc33bits_113_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_113_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_113_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_113_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_113_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_113_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_113_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_113_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_113_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_113_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_113_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_113_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_113_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_113_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_113_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_113_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_113_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_113_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_113_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_113_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_113_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_113_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_113_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_113_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_113_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_113_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_113_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_113_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_113_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_113_io_cout_group_29),
    .io_cout(Walloc33bits_113_io_cout),
    .io_s(Walloc33bits_113_io_s)
  );
  Walloc33bits Walloc33bits_114 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_114_io_src_in),
    .io_cin(Walloc33bits_114_io_cin),
    .io_cout_group_0(Walloc33bits_114_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_114_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_114_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_114_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_114_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_114_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_114_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_114_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_114_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_114_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_114_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_114_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_114_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_114_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_114_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_114_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_114_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_114_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_114_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_114_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_114_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_114_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_114_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_114_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_114_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_114_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_114_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_114_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_114_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_114_io_cout_group_29),
    .io_cout(Walloc33bits_114_io_cout),
    .io_s(Walloc33bits_114_io_s)
  );
  Walloc33bits Walloc33bits_115 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_115_io_src_in),
    .io_cin(Walloc33bits_115_io_cin),
    .io_cout_group_0(Walloc33bits_115_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_115_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_115_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_115_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_115_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_115_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_115_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_115_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_115_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_115_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_115_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_115_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_115_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_115_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_115_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_115_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_115_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_115_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_115_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_115_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_115_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_115_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_115_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_115_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_115_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_115_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_115_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_115_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_115_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_115_io_cout_group_29),
    .io_cout(Walloc33bits_115_io_cout),
    .io_s(Walloc33bits_115_io_s)
  );
  Walloc33bits Walloc33bits_116 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_116_io_src_in),
    .io_cin(Walloc33bits_116_io_cin),
    .io_cout_group_0(Walloc33bits_116_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_116_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_116_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_116_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_116_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_116_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_116_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_116_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_116_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_116_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_116_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_116_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_116_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_116_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_116_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_116_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_116_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_116_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_116_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_116_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_116_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_116_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_116_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_116_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_116_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_116_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_116_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_116_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_116_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_116_io_cout_group_29),
    .io_cout(Walloc33bits_116_io_cout),
    .io_s(Walloc33bits_116_io_s)
  );
  Walloc33bits Walloc33bits_117 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_117_io_src_in),
    .io_cin(Walloc33bits_117_io_cin),
    .io_cout_group_0(Walloc33bits_117_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_117_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_117_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_117_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_117_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_117_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_117_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_117_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_117_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_117_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_117_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_117_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_117_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_117_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_117_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_117_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_117_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_117_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_117_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_117_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_117_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_117_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_117_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_117_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_117_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_117_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_117_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_117_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_117_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_117_io_cout_group_29),
    .io_cout(Walloc33bits_117_io_cout),
    .io_s(Walloc33bits_117_io_s)
  );
  Walloc33bits Walloc33bits_118 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_118_io_src_in),
    .io_cin(Walloc33bits_118_io_cin),
    .io_cout_group_0(Walloc33bits_118_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_118_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_118_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_118_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_118_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_118_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_118_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_118_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_118_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_118_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_118_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_118_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_118_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_118_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_118_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_118_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_118_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_118_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_118_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_118_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_118_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_118_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_118_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_118_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_118_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_118_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_118_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_118_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_118_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_118_io_cout_group_29),
    .io_cout(Walloc33bits_118_io_cout),
    .io_s(Walloc33bits_118_io_s)
  );
  Walloc33bits Walloc33bits_119 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_119_io_src_in),
    .io_cin(Walloc33bits_119_io_cin),
    .io_cout_group_0(Walloc33bits_119_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_119_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_119_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_119_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_119_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_119_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_119_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_119_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_119_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_119_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_119_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_119_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_119_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_119_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_119_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_119_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_119_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_119_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_119_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_119_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_119_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_119_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_119_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_119_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_119_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_119_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_119_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_119_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_119_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_119_io_cout_group_29),
    .io_cout(Walloc33bits_119_io_cout),
    .io_s(Walloc33bits_119_io_s)
  );
  Walloc33bits Walloc33bits_120 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_120_io_src_in),
    .io_cin(Walloc33bits_120_io_cin),
    .io_cout_group_0(Walloc33bits_120_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_120_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_120_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_120_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_120_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_120_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_120_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_120_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_120_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_120_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_120_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_120_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_120_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_120_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_120_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_120_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_120_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_120_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_120_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_120_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_120_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_120_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_120_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_120_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_120_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_120_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_120_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_120_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_120_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_120_io_cout_group_29),
    .io_cout(Walloc33bits_120_io_cout),
    .io_s(Walloc33bits_120_io_s)
  );
  Walloc33bits Walloc33bits_121 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_121_io_src_in),
    .io_cin(Walloc33bits_121_io_cin),
    .io_cout_group_0(Walloc33bits_121_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_121_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_121_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_121_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_121_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_121_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_121_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_121_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_121_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_121_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_121_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_121_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_121_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_121_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_121_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_121_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_121_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_121_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_121_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_121_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_121_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_121_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_121_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_121_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_121_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_121_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_121_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_121_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_121_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_121_io_cout_group_29),
    .io_cout(Walloc33bits_121_io_cout),
    .io_s(Walloc33bits_121_io_s)
  );
  Walloc33bits Walloc33bits_122 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_122_io_src_in),
    .io_cin(Walloc33bits_122_io_cin),
    .io_cout_group_0(Walloc33bits_122_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_122_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_122_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_122_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_122_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_122_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_122_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_122_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_122_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_122_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_122_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_122_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_122_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_122_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_122_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_122_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_122_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_122_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_122_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_122_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_122_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_122_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_122_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_122_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_122_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_122_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_122_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_122_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_122_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_122_io_cout_group_29),
    .io_cout(Walloc33bits_122_io_cout),
    .io_s(Walloc33bits_122_io_s)
  );
  Walloc33bits Walloc33bits_123 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_123_io_src_in),
    .io_cin(Walloc33bits_123_io_cin),
    .io_cout_group_0(Walloc33bits_123_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_123_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_123_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_123_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_123_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_123_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_123_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_123_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_123_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_123_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_123_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_123_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_123_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_123_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_123_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_123_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_123_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_123_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_123_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_123_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_123_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_123_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_123_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_123_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_123_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_123_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_123_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_123_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_123_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_123_io_cout_group_29),
    .io_cout(Walloc33bits_123_io_cout),
    .io_s(Walloc33bits_123_io_s)
  );
  Walloc33bits Walloc33bits_124 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_124_io_src_in),
    .io_cin(Walloc33bits_124_io_cin),
    .io_cout_group_0(Walloc33bits_124_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_124_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_124_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_124_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_124_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_124_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_124_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_124_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_124_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_124_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_124_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_124_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_124_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_124_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_124_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_124_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_124_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_124_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_124_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_124_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_124_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_124_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_124_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_124_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_124_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_124_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_124_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_124_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_124_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_124_io_cout_group_29),
    .io_cout(Walloc33bits_124_io_cout),
    .io_s(Walloc33bits_124_io_s)
  );
  Walloc33bits Walloc33bits_125 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_125_io_src_in),
    .io_cin(Walloc33bits_125_io_cin),
    .io_cout_group_0(Walloc33bits_125_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_125_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_125_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_125_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_125_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_125_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_125_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_125_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_125_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_125_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_125_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_125_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_125_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_125_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_125_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_125_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_125_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_125_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_125_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_125_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_125_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_125_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_125_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_125_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_125_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_125_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_125_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_125_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_125_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_125_io_cout_group_29),
    .io_cout(Walloc33bits_125_io_cout),
    .io_s(Walloc33bits_125_io_s)
  );
  Walloc33bits Walloc33bits_126 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_126_io_src_in),
    .io_cin(Walloc33bits_126_io_cin),
    .io_cout_group_0(Walloc33bits_126_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_126_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_126_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_126_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_126_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_126_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_126_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_126_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_126_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_126_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_126_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_126_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_126_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_126_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_126_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_126_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_126_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_126_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_126_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_126_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_126_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_126_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_126_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_126_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_126_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_126_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_126_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_126_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_126_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_126_io_cout_group_29),
    .io_cout(Walloc33bits_126_io_cout),
    .io_s(Walloc33bits_126_io_s)
  );
  Walloc33bits Walloc33bits_127 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_127_io_src_in),
    .io_cin(Walloc33bits_127_io_cin),
    .io_cout_group_0(Walloc33bits_127_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_127_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_127_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_127_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_127_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_127_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_127_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_127_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_127_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_127_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_127_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_127_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_127_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_127_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_127_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_127_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_127_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_127_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_127_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_127_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_127_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_127_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_127_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_127_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_127_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_127_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_127_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_127_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_127_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_127_io_cout_group_29),
    .io_cout(Walloc33bits_127_io_cout),
    .io_s(Walloc33bits_127_io_s)
  );
  Walloc33bits Walloc33bits_128 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_128_io_src_in),
    .io_cin(Walloc33bits_128_io_cin),
    .io_cout_group_0(Walloc33bits_128_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_128_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_128_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_128_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_128_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_128_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_128_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_128_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_128_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_128_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_128_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_128_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_128_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_128_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_128_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_128_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_128_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_128_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_128_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_128_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_128_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_128_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_128_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_128_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_128_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_128_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_128_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_128_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_128_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_128_io_cout_group_29),
    .io_cout(Walloc33bits_128_io_cout),
    .io_s(Walloc33bits_128_io_s)
  );
  Walloc33bits Walloc33bits_129 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_129_io_src_in),
    .io_cin(Walloc33bits_129_io_cin),
    .io_cout_group_0(Walloc33bits_129_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_129_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_129_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_129_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_129_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_129_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_129_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_129_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_129_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_129_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_129_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_129_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_129_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_129_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_129_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_129_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_129_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_129_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_129_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_129_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_129_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_129_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_129_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_129_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_129_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_129_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_129_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_129_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_129_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_129_io_cout_group_29),
    .io_cout(Walloc33bits_129_io_cout),
    .io_s(Walloc33bits_129_io_s)
  );
  Walloc33bits Walloc33bits_130 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_130_io_src_in),
    .io_cin(Walloc33bits_130_io_cin),
    .io_cout_group_0(Walloc33bits_130_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_130_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_130_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_130_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_130_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_130_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_130_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_130_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_130_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_130_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_130_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_130_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_130_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_130_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_130_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_130_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_130_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_130_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_130_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_130_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_130_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_130_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_130_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_130_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_130_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_130_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_130_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_130_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_130_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_130_io_cout_group_29),
    .io_cout(Walloc33bits_130_io_cout),
    .io_s(Walloc33bits_130_io_s)
  );
  Walloc33bits Walloc33bits_131 ( // @[WallaceTest.scala 206:30]
    .io_src_in(Walloc33bits_131_io_src_in),
    .io_cin(Walloc33bits_131_io_cin),
    .io_cout_group_0(Walloc33bits_131_io_cout_group_0),
    .io_cout_group_1(Walloc33bits_131_io_cout_group_1),
    .io_cout_group_2(Walloc33bits_131_io_cout_group_2),
    .io_cout_group_3(Walloc33bits_131_io_cout_group_3),
    .io_cout_group_4(Walloc33bits_131_io_cout_group_4),
    .io_cout_group_5(Walloc33bits_131_io_cout_group_5),
    .io_cout_group_6(Walloc33bits_131_io_cout_group_6),
    .io_cout_group_7(Walloc33bits_131_io_cout_group_7),
    .io_cout_group_8(Walloc33bits_131_io_cout_group_8),
    .io_cout_group_9(Walloc33bits_131_io_cout_group_9),
    .io_cout_group_10(Walloc33bits_131_io_cout_group_10),
    .io_cout_group_11(Walloc33bits_131_io_cout_group_11),
    .io_cout_group_12(Walloc33bits_131_io_cout_group_12),
    .io_cout_group_13(Walloc33bits_131_io_cout_group_13),
    .io_cout_group_14(Walloc33bits_131_io_cout_group_14),
    .io_cout_group_15(Walloc33bits_131_io_cout_group_15),
    .io_cout_group_16(Walloc33bits_131_io_cout_group_16),
    .io_cout_group_17(Walloc33bits_131_io_cout_group_17),
    .io_cout_group_18(Walloc33bits_131_io_cout_group_18),
    .io_cout_group_19(Walloc33bits_131_io_cout_group_19),
    .io_cout_group_20(Walloc33bits_131_io_cout_group_20),
    .io_cout_group_21(Walloc33bits_131_io_cout_group_21),
    .io_cout_group_22(Walloc33bits_131_io_cout_group_22),
    .io_cout_group_23(Walloc33bits_131_io_cout_group_23),
    .io_cout_group_24(Walloc33bits_131_io_cout_group_24),
    .io_cout_group_25(Walloc33bits_131_io_cout_group_25),
    .io_cout_group_26(Walloc33bits_131_io_cout_group_26),
    .io_cout_group_27(Walloc33bits_131_io_cout_group_27),
    .io_cout_group_28(Walloc33bits_131_io_cout_group_28),
    .io_cout_group_29(Walloc33bits_131_io_cout_group_29),
    .io_cout(Walloc33bits_131_io_cout),
    .io_s(Walloc33bits_131_io_s)
  );
  assign io_result_hi = result[127:64]; // @[WallaceTest.scala 232:25]
  assign io_result_lo = result[63:0]; // @[WallaceTest.scala 233:25]
  assign gen_p_io_src = mulb[2:0]; // @[WallaceTest.scala 212:20]
  assign gen_p_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_1_io_src = mulb[4:2]; // @[WallaceTest.scala 212:20]
  assign gen_p_1_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_2_io_src = mulb[6:4]; // @[WallaceTest.scala 212:20]
  assign gen_p_2_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_3_io_src = mulb[8:6]; // @[WallaceTest.scala 212:20]
  assign gen_p_3_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_4_io_src = mulb[10:8]; // @[WallaceTest.scala 212:20]
  assign gen_p_4_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_5_io_src = mulb[12:10]; // @[WallaceTest.scala 212:20]
  assign gen_p_5_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_6_io_src = mulb[14:12]; // @[WallaceTest.scala 212:20]
  assign gen_p_6_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_7_io_src = mulb[16:14]; // @[WallaceTest.scala 212:20]
  assign gen_p_7_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_8_io_src = mulb[18:16]; // @[WallaceTest.scala 212:20]
  assign gen_p_8_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_9_io_src = mulb[20:18]; // @[WallaceTest.scala 212:20]
  assign gen_p_9_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_10_io_src = mulb[22:20]; // @[WallaceTest.scala 212:20]
  assign gen_p_10_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_11_io_src = mulb[24:22]; // @[WallaceTest.scala 212:20]
  assign gen_p_11_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_12_io_src = mulb[26:24]; // @[WallaceTest.scala 212:20]
  assign gen_p_12_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_13_io_src = mulb[28:26]; // @[WallaceTest.scala 212:20]
  assign gen_p_13_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_14_io_src = mulb[30:28]; // @[WallaceTest.scala 212:20]
  assign gen_p_14_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_15_io_src = mulb[32:30]; // @[WallaceTest.scala 212:20]
  assign gen_p_15_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_16_io_src = mulb[34:32]; // @[WallaceTest.scala 212:20]
  assign gen_p_16_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_17_io_src = mulb[36:34]; // @[WallaceTest.scala 212:20]
  assign gen_p_17_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_18_io_src = mulb[38:36]; // @[WallaceTest.scala 212:20]
  assign gen_p_18_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_19_io_src = mulb[40:38]; // @[WallaceTest.scala 212:20]
  assign gen_p_19_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_20_io_src = mulb[42:40]; // @[WallaceTest.scala 212:20]
  assign gen_p_20_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_21_io_src = mulb[44:42]; // @[WallaceTest.scala 212:20]
  assign gen_p_21_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_22_io_src = mulb[46:44]; // @[WallaceTest.scala 212:20]
  assign gen_p_22_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_23_io_src = mulb[48:46]; // @[WallaceTest.scala 212:20]
  assign gen_p_23_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_24_io_src = mulb[50:48]; // @[WallaceTest.scala 212:20]
  assign gen_p_24_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_25_io_src = mulb[52:50]; // @[WallaceTest.scala 212:20]
  assign gen_p_25_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_26_io_src = mulb[54:52]; // @[WallaceTest.scala 212:20]
  assign gen_p_26_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_27_io_src = mulb[56:54]; // @[WallaceTest.scala 212:20]
  assign gen_p_27_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_28_io_src = mulb[58:56]; // @[WallaceTest.scala 212:20]
  assign gen_p_28_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_29_io_src = mulb[60:58]; // @[WallaceTest.scala 212:20]
  assign gen_p_29_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_30_io_src = mulb[62:60]; // @[WallaceTest.scala 212:20]
  assign gen_p_30_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_31_io_src = mulb[64:62]; // @[WallaceTest.scala 212:20]
  assign gen_p_31_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign gen_p_32_io_src = mulb[66:64]; // @[WallaceTest.scala 212:20]
  assign gen_p_32_io_x = io_multiplicand; // @[WallaceTest.scala 213:12]
  assign switch_clock = clock;
  assign switch_reset = reset;
  assign switch_io_in_0 = gen_p_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_1 = gen_p_1_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_2 = gen_p_2_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_3 = gen_p_3_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_4 = gen_p_4_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_5 = gen_p_5_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_6 = gen_p_6_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_7 = gen_p_7_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_8 = gen_p_8_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_9 = gen_p_9_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_10 = gen_p_10_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_11 = gen_p_11_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_12 = gen_p_12_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_13 = gen_p_13_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_14 = gen_p_14_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_15 = gen_p_15_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_16 = gen_p_16_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_17 = gen_p_17_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_18 = gen_p_18_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_19 = gen_p_19_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_20 = gen_p_20_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_21 = gen_p_21_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_22 = gen_p_22_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_23 = gen_p_23_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_24 = gen_p_24_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_25 = gen_p_25_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_26 = gen_p_26_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_27 = gen_p_27_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_28 = gen_p_28_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_29 = gen_p_29_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_30 = gen_p_30_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_31 = gen_p_31_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_in_32 = gen_p_32_io_p; // @[WallaceTest.scala 214:13]
  assign switch_io_cin_0 = gen_p_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_1 = gen_p_1_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_2 = gen_p_2_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_3 = gen_p_3_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_4 = gen_p_4_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_5 = gen_p_5_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_6 = gen_p_6_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_7 = gen_p_7_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_8 = gen_p_8_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_9 = gen_p_9_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_10 = gen_p_10_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_11 = gen_p_11_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_12 = gen_p_12_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_13 = gen_p_13_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_14 = gen_p_14_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_15 = gen_p_15_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_16 = gen_p_16_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_17 = gen_p_17_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_18 = gen_p_18_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_19 = gen_p_19_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_20 = gen_p_20_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_21 = gen_p_21_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_22 = gen_p_22_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_23 = gen_p_23_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_24 = gen_p_24_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_25 = gen_p_25_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_26 = gen_p_26_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_27 = gen_p_27_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_28 = gen_p_28_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_29 = gen_p_29_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_30 = gen_p_30_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_31 = gen_p_31_io_c; // @[WallaceTest.scala 215:14]
  assign switch_io_cin_32 = gen_p_32_io_c; // @[WallaceTest.scala 215:14]
  assign Walloc33bits_io_src_in = switch_io_out_0; // @[WallaceTest.scala 218:16]
  assign Walloc33bits_io_cin = switch_io_cout[31:2]; // @[WallaceTest.scala 219:23]
  assign Walloc33bits_1_io_src_in = switch_io_out_1; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_1_io_cin = {hi,lo}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_2_io_src_in = switch_io_out_2; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_2_io_cin = {hi_1,lo_1}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_3_io_src_in = switch_io_out_3; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_3_io_cin = {hi_2,lo_2}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_4_io_src_in = switch_io_out_4; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_4_io_cin = {hi_3,lo_3}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_5_io_src_in = switch_io_out_5; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_5_io_cin = {hi_4,lo_4}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_6_io_src_in = switch_io_out_6; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_6_io_cin = {hi_5,lo_5}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_7_io_src_in = switch_io_out_7; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_7_io_cin = {hi_6,lo_6}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_8_io_src_in = switch_io_out_8; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_8_io_cin = {hi_7,lo_7}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_9_io_src_in = switch_io_out_9; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_9_io_cin = {hi_8,lo_8}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_10_io_src_in = switch_io_out_10; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_10_io_cin = {hi_9,lo_9}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_11_io_src_in = switch_io_out_11; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_11_io_cin = {hi_10,lo_10}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_12_io_src_in = switch_io_out_12; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_12_io_cin = {hi_11,lo_11}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_13_io_src_in = switch_io_out_13; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_13_io_cin = {hi_12,lo_12}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_14_io_src_in = switch_io_out_14; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_14_io_cin = {hi_13,lo_13}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_15_io_src_in = switch_io_out_15; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_15_io_cin = {hi_14,lo_14}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_16_io_src_in = switch_io_out_16; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_16_io_cin = {hi_15,lo_15}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_17_io_src_in = switch_io_out_17; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_17_io_cin = {hi_16,lo_16}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_18_io_src_in = switch_io_out_18; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_18_io_cin = {hi_17,lo_17}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_19_io_src_in = switch_io_out_19; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_19_io_cin = {hi_18,lo_18}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_20_io_src_in = switch_io_out_20; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_20_io_cin = {hi_19,lo_19}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_21_io_src_in = switch_io_out_21; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_21_io_cin = {hi_20,lo_20}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_22_io_src_in = switch_io_out_22; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_22_io_cin = {hi_21,lo_21}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_23_io_src_in = switch_io_out_23; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_23_io_cin = {hi_22,lo_22}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_24_io_src_in = switch_io_out_24; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_24_io_cin = {hi_23,lo_23}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_25_io_src_in = switch_io_out_25; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_25_io_cin = {hi_24,lo_24}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_26_io_src_in = switch_io_out_26; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_26_io_cin = {hi_25,lo_25}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_27_io_src_in = switch_io_out_27; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_27_io_cin = {hi_26,lo_26}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_28_io_src_in = switch_io_out_28; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_28_io_cin = {hi_27,lo_27}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_29_io_src_in = switch_io_out_29; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_29_io_cin = {hi_28,lo_28}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_30_io_src_in = switch_io_out_30; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_30_io_cin = {hi_29,lo_29}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_31_io_src_in = switch_io_out_31; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_31_io_cin = {hi_30,lo_30}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_32_io_src_in = switch_io_out_32; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_32_io_cin = {hi_31,lo_31}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_33_io_src_in = switch_io_out_33; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_33_io_cin = {hi_32,lo_32}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_34_io_src_in = switch_io_out_34; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_34_io_cin = {hi_33,lo_33}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_35_io_src_in = switch_io_out_35; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_35_io_cin = {hi_34,lo_34}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_36_io_src_in = switch_io_out_36; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_36_io_cin = {hi_35,lo_35}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_37_io_src_in = switch_io_out_37; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_37_io_cin = {hi_36,lo_36}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_38_io_src_in = switch_io_out_38; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_38_io_cin = {hi_37,lo_37}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_39_io_src_in = switch_io_out_39; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_39_io_cin = {hi_38,lo_38}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_40_io_src_in = switch_io_out_40; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_40_io_cin = {hi_39,lo_39}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_41_io_src_in = switch_io_out_41; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_41_io_cin = {hi_40,lo_40}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_42_io_src_in = switch_io_out_42; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_42_io_cin = {hi_41,lo_41}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_43_io_src_in = switch_io_out_43; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_43_io_cin = {hi_42,lo_42}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_44_io_src_in = switch_io_out_44; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_44_io_cin = {hi_43,lo_43}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_45_io_src_in = switch_io_out_45; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_45_io_cin = {hi_44,lo_44}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_46_io_src_in = switch_io_out_46; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_46_io_cin = {hi_45,lo_45}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_47_io_src_in = switch_io_out_47; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_47_io_cin = {hi_46,lo_46}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_48_io_src_in = switch_io_out_48; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_48_io_cin = {hi_47,lo_47}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_49_io_src_in = switch_io_out_49; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_49_io_cin = {hi_48,lo_48}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_50_io_src_in = switch_io_out_50; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_50_io_cin = {hi_49,lo_49}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_51_io_src_in = switch_io_out_51; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_51_io_cin = {hi_50,lo_50}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_52_io_src_in = switch_io_out_52; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_52_io_cin = {hi_51,lo_51}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_53_io_src_in = switch_io_out_53; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_53_io_cin = {hi_52,lo_52}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_54_io_src_in = switch_io_out_54; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_54_io_cin = {hi_53,lo_53}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_55_io_src_in = switch_io_out_55; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_55_io_cin = {hi_54,lo_54}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_56_io_src_in = switch_io_out_56; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_56_io_cin = {hi_55,lo_55}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_57_io_src_in = switch_io_out_57; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_57_io_cin = {hi_56,lo_56}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_58_io_src_in = switch_io_out_58; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_58_io_cin = {hi_57,lo_57}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_59_io_src_in = switch_io_out_59; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_59_io_cin = {hi_58,lo_58}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_60_io_src_in = switch_io_out_60; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_60_io_cin = {hi_59,lo_59}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_61_io_src_in = switch_io_out_61; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_61_io_cin = {hi_60,lo_60}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_62_io_src_in = switch_io_out_62; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_62_io_cin = {hi_61,lo_61}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_63_io_src_in = switch_io_out_63; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_63_io_cin = {hi_62,lo_62}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_64_io_src_in = switch_io_out_64; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_64_io_cin = {hi_63,lo_63}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_65_io_src_in = switch_io_out_65; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_65_io_cin = {hi_64,lo_64}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_66_io_src_in = switch_io_out_66; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_66_io_cin = {hi_65,lo_65}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_67_io_src_in = switch_io_out_67; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_67_io_cin = {hi_66,lo_66}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_68_io_src_in = switch_io_out_68; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_68_io_cin = {hi_67,lo_67}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_69_io_src_in = switch_io_out_69; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_69_io_cin = {hi_68,lo_68}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_70_io_src_in = switch_io_out_70; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_70_io_cin = {hi_69,lo_69}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_71_io_src_in = switch_io_out_71; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_71_io_cin = {hi_70,lo_70}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_72_io_src_in = switch_io_out_72; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_72_io_cin = {hi_71,lo_71}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_73_io_src_in = switch_io_out_73; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_73_io_cin = {hi_72,lo_72}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_74_io_src_in = switch_io_out_74; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_74_io_cin = {hi_73,lo_73}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_75_io_src_in = switch_io_out_75; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_75_io_cin = {hi_74,lo_74}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_76_io_src_in = switch_io_out_76; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_76_io_cin = {hi_75,lo_75}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_77_io_src_in = switch_io_out_77; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_77_io_cin = {hi_76,lo_76}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_78_io_src_in = switch_io_out_78; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_78_io_cin = {hi_77,lo_77}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_79_io_src_in = switch_io_out_79; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_79_io_cin = {hi_78,lo_78}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_80_io_src_in = switch_io_out_80; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_80_io_cin = {hi_79,lo_79}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_81_io_src_in = switch_io_out_81; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_81_io_cin = {hi_80,lo_80}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_82_io_src_in = switch_io_out_82; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_82_io_cin = {hi_81,lo_81}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_83_io_src_in = switch_io_out_83; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_83_io_cin = {hi_82,lo_82}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_84_io_src_in = switch_io_out_84; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_84_io_cin = {hi_83,lo_83}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_85_io_src_in = switch_io_out_85; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_85_io_cin = {hi_84,lo_84}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_86_io_src_in = switch_io_out_86; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_86_io_cin = {hi_85,lo_85}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_87_io_src_in = switch_io_out_87; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_87_io_cin = {hi_86,lo_86}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_88_io_src_in = switch_io_out_88; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_88_io_cin = {hi_87,lo_87}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_89_io_src_in = switch_io_out_89; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_89_io_cin = {hi_88,lo_88}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_90_io_src_in = switch_io_out_90; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_90_io_cin = {hi_89,lo_89}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_91_io_src_in = switch_io_out_91; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_91_io_cin = {hi_90,lo_90}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_92_io_src_in = switch_io_out_92; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_92_io_cin = {hi_91,lo_91}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_93_io_src_in = switch_io_out_93; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_93_io_cin = {hi_92,lo_92}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_94_io_src_in = switch_io_out_94; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_94_io_cin = {hi_93,lo_93}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_95_io_src_in = switch_io_out_95; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_95_io_cin = {hi_94,lo_94}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_96_io_src_in = switch_io_out_96; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_96_io_cin = {hi_95,lo_95}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_97_io_src_in = switch_io_out_97; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_97_io_cin = {hi_96,lo_96}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_98_io_src_in = switch_io_out_98; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_98_io_cin = {hi_97,lo_97}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_99_io_src_in = switch_io_out_99; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_99_io_cin = {hi_98,lo_98}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_100_io_src_in = switch_io_out_100; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_100_io_cin = {hi_99,lo_99}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_101_io_src_in = switch_io_out_101; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_101_io_cin = {hi_100,lo_100}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_102_io_src_in = switch_io_out_102; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_102_io_cin = {hi_101,lo_101}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_103_io_src_in = switch_io_out_103; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_103_io_cin = {hi_102,lo_102}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_104_io_src_in = switch_io_out_104; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_104_io_cin = {hi_103,lo_103}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_105_io_src_in = switch_io_out_105; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_105_io_cin = {hi_104,lo_104}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_106_io_src_in = switch_io_out_106; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_106_io_cin = {hi_105,lo_105}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_107_io_src_in = switch_io_out_107; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_107_io_cin = {hi_106,lo_106}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_108_io_src_in = switch_io_out_108; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_108_io_cin = {hi_107,lo_107}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_109_io_src_in = switch_io_out_109; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_109_io_cin = {hi_108,lo_108}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_110_io_src_in = switch_io_out_110; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_110_io_cin = {hi_109,lo_109}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_111_io_src_in = switch_io_out_111; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_111_io_cin = {hi_110,lo_110}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_112_io_src_in = switch_io_out_112; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_112_io_cin = {hi_111,lo_111}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_113_io_src_in = switch_io_out_113; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_113_io_cin = {hi_112,lo_112}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_114_io_src_in = switch_io_out_114; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_114_io_cin = {hi_113,lo_113}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_115_io_src_in = switch_io_out_115; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_115_io_cin = {hi_114,lo_114}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_116_io_src_in = switch_io_out_116; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_116_io_cin = {hi_115,lo_115}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_117_io_src_in = switch_io_out_117; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_117_io_cin = {hi_116,lo_116}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_118_io_src_in = switch_io_out_118; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_118_io_cin = {hi_117,lo_117}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_119_io_src_in = switch_io_out_119; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_119_io_cin = {hi_118,lo_118}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_120_io_src_in = switch_io_out_120; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_120_io_cin = {hi_119,lo_119}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_121_io_src_in = switch_io_out_121; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_121_io_cin = {hi_120,lo_120}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_122_io_src_in = switch_io_out_122; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_122_io_cin = {hi_121,lo_121}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_123_io_src_in = switch_io_out_123; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_123_io_cin = {hi_122,lo_122}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_124_io_src_in = switch_io_out_124; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_124_io_cin = {hi_123,lo_123}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_125_io_src_in = switch_io_out_125; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_125_io_cin = {hi_124,lo_124}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_126_io_src_in = switch_io_out_126; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_126_io_cin = {hi_125,lo_125}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_127_io_src_in = switch_io_out_127; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_127_io_cin = {hi_126,lo_126}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_128_io_src_in = switch_io_out_128; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_128_io_cin = {hi_127,lo_127}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_129_io_src_in = switch_io_out_129; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_129_io_cin = {hi_128,lo_128}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_130_io_src_in = switch_io_out_130; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_130_io_cin = {hi_129,lo_129}; // @[WallaceTest.scala 224:37]
  assign Walloc33bits_131_io_src_in = switch_io_out_131; // @[WallaceTest.scala 223:18]
  assign Walloc33bits_131_io_cin = {hi_130,lo_130}; // @[WallaceTest.scala 224:37]
endmodule
module unit(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input         io_flush,
  input         io_mulw,
  input  [1:0]  io_mul_signed,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_mul_ready,
  output        io_out_valid,
  output [63:0] io_result_hi,
  output [63:0] io_result_lo
);
  wire  walloc_64_mul_clock; // @[WallaceTest.scala 265:20]
  wire  walloc_64_mul_reset; // @[WallaceTest.scala 265:20]
  wire [131:0] walloc_64_mul_io_multiplicand; // @[WallaceTest.scala 265:20]
  wire [65:0] walloc_64_mul_io_multiplier; // @[WallaceTest.scala 265:20]
  wire [63:0] walloc_64_mul_io_result_hi; // @[WallaceTest.scala 265:20]
  wire [63:0] walloc_64_mul_io_result_lo; // @[WallaceTest.scala 265:20]
  wire  _a_T_2 = io_mul_valid & io_mul_signed[1]; // @[WallaceTest.scala 254:24]
  wire  _a_T_3 = io_mul_valid & io_mul_signed[1] & io_mulw; // @[WallaceTest.scala 254:41]
  wire [99:0] _a_T_7 = io_multiplicand[31] ? 100'hfffffffffffffffffffffffff : 100'h0; // @[Bitwise.scala 77:12]
  wire [163:0] _a_T_8 = {_a_T_7,io_multiplicand}; // @[Cat.scala 33:92]
  wire  _a_T_12 = _a_T_2 & ~io_mulw; // @[WallaceTest.scala 255:41]
  wire [67:0] _a_T_16 = io_multiplicand[63] ? 68'hfffffffffffffffff : 68'h0; // @[Bitwise.scala 77:12]
  wire [131:0] _a_T_17 = {_a_T_16,io_multiplicand}; // @[Cat.scala 33:92]
  wire [63:0] _a_T_19 = io_mul_valid ? io_multiplicand : 64'h0; // @[WallaceTest.scala 256:10]
  wire [131:0] _a_T_20 = _a_T_2 & ~io_mulw ? _a_T_17 : {{68'd0}, _a_T_19}; // @[WallaceTest.scala 255:10]
  wire [163:0] _a_T_21 = io_mul_valid & io_mul_signed[1] & io_mulw ? _a_T_8 : {{32'd0}, _a_T_20}; // @[WallaceTest.scala 254:10]
  wire [163:0] _a_T_22 = io_flush ? 164'h0 : _a_T_21; // @[WallaceTest.scala 253:10]
  wire [99:0] _b_T_7 = io_multiplier[31] ? 100'hfffffffffffffffffffffffff : 100'h0; // @[Bitwise.scala 77:12]
  wire [163:0] _b_T_8 = {_b_T_7,io_multiplier}; // @[Cat.scala 33:92]
  wire [67:0] _b_T_16 = io_multiplier[63] ? 68'hfffffffffffffffff : 68'h0; // @[Bitwise.scala 77:12]
  wire [131:0] _b_T_17 = {_b_T_16,io_multiplier}; // @[Cat.scala 33:92]
  wire [63:0] _b_T_19 = io_mul_valid ? io_multiplier : 64'h0; // @[WallaceTest.scala 262:10]
  wire [131:0] _b_T_20 = _a_T_12 ? _b_T_17 : {{68'd0}, _b_T_19}; // @[WallaceTest.scala 261:10]
  wire [163:0] _b_T_21 = _a_T_3 ? _b_T_8 : {{32'd0}, _b_T_20}; // @[WallaceTest.scala 260:10]
  wire [163:0] _b_T_22 = io_flush ? 164'h0 : _b_T_21; // @[WallaceTest.scala 259:10]
  walloc_64_mul walloc_64_mul ( // @[WallaceTest.scala 265:20]
    .clock(walloc_64_mul_clock),
    .reset(walloc_64_mul_reset),
    .io_multiplicand(walloc_64_mul_io_multiplicand),
    .io_multiplier(walloc_64_mul_io_multiplier),
    .io_result_hi(walloc_64_mul_io_result_hi),
    .io_result_lo(walloc_64_mul_io_result_lo)
  );
  assign io_mul_ready = 1'h1; // @[WallaceTest.scala 273:15]
  assign io_out_valid = io_mul_valid; // @[WallaceTest.scala 272:15]
  assign io_result_hi = walloc_64_mul_io_result_hi; // @[WallaceTest.scala 269:15]
  assign io_result_lo = walloc_64_mul_io_result_lo; // @[WallaceTest.scala 270:15]
  assign walloc_64_mul_clock = clock;
  assign walloc_64_mul_reset = reset;
  assign walloc_64_mul_io_multiplicand = _a_T_22[131:0]; // @[WallaceTest.scala 250:15 253:5]
  assign walloc_64_mul_io_multiplier = _b_T_22[65:0]; // @[WallaceTest.scala 251:15 259:5]
endmodule
